magic
tech scmos
timestamp 1625156677
<< metal1 >>
rect 856 3703 858 3707
rect 862 3703 865 3707
rect 869 3703 872 3707
rect 1872 3703 1874 3707
rect 1878 3703 1881 3707
rect 1885 3703 1888 3707
rect 2904 3703 2906 3707
rect 2910 3703 2913 3707
rect 2917 3703 2920 3707
rect 3928 3703 3930 3707
rect 3934 3703 3937 3707
rect 3941 3703 3944 3707
rect 4952 3703 4954 3707
rect 4958 3703 4961 3707
rect 4965 3703 4968 3707
rect 492 3688 494 3692
rect 698 3688 719 3691
rect 1108 3688 1110 3692
rect 1780 3688 1782 3692
rect 2946 3688 2953 3691
rect 3294 3688 3302 3691
rect 302 3678 313 3681
rect 398 3671 401 3681
rect 370 3668 385 3671
rect 398 3668 406 3671
rect 510 3668 529 3671
rect 570 3668 577 3671
rect 686 3668 702 3671
rect 766 3671 769 3681
rect 1542 3678 1553 3681
rect 1626 3678 1630 3682
rect 3110 3678 3118 3681
rect 3318 3678 3326 3681
rect 4090 3678 4097 3681
rect 4186 3678 4193 3681
rect 4710 3678 4718 3681
rect 5042 3678 5043 3682
rect 766 3668 774 3671
rect 782 3668 790 3671
rect 1350 3668 1377 3671
rect 170 3658 177 3661
rect 270 3658 281 3661
rect 670 3661 673 3668
rect 1478 3662 1481 3671
rect 1510 3668 1521 3671
rect 1610 3668 1617 3671
rect 670 3658 681 3661
rect 902 3658 921 3661
rect 926 3658 942 3661
rect 982 3658 990 3661
rect 1150 3658 1158 3661
rect 1450 3658 1465 3661
rect 1582 3658 1590 3661
rect 1742 3661 1745 3671
rect 2438 3668 2446 3671
rect 2686 3668 2694 3671
rect 3518 3668 3530 3671
rect 3742 3671 3746 3674
rect 3738 3668 3746 3671
rect 3934 3668 3950 3671
rect 4398 3668 4409 3671
rect 4450 3668 4473 3671
rect 4558 3668 4566 3671
rect 1742 3658 1750 3661
rect 1862 3661 1865 3668
rect 1862 3658 1873 3661
rect 1942 3658 1950 3661
rect 1986 3658 1993 3661
rect 2098 3658 2105 3661
rect 2582 3658 2590 3661
rect 2642 3658 2649 3661
rect 2766 3658 2778 3661
rect 3270 3658 3281 3661
rect 3406 3658 3434 3661
rect 3726 3658 3746 3661
rect 3934 3658 3966 3661
rect 4326 3661 4329 3668
rect 4398 3662 4402 3664
rect 4318 3658 4329 3661
rect 4458 3658 4473 3661
rect 4558 3658 4574 3661
rect 5054 3658 5062 3661
rect 5158 3658 5169 3661
rect 270 3656 274 3658
rect 1726 3652 1729 3658
rect 758 3648 766 3651
rect 894 3648 905 3651
rect 1254 3648 1265 3651
rect 1302 3648 1313 3651
rect 1350 3648 1358 3651
rect 1401 3648 1406 3652
rect 1530 3648 1534 3652
rect 1542 3648 1553 3651
rect 1590 3648 1601 3651
rect 1721 3648 1729 3652
rect 2174 3648 2177 3658
rect 2774 3657 2778 3658
rect 3270 3657 3274 3658
rect 3430 3657 3434 3658
rect 3742 3657 3746 3658
rect 5158 3657 5162 3658
rect 2234 3648 2241 3651
rect 2350 3648 2366 3651
rect 2874 3648 2881 3651
rect 338 3638 366 3641
rect 1270 3641 1273 3648
rect 1550 3642 1553 3648
rect 1262 3638 1273 3641
rect 1822 3638 1838 3641
rect 2122 3638 2150 3641
rect 2318 3641 2321 3648
rect 2310 3638 2321 3641
rect 2486 3638 2494 3641
rect 3762 3638 3765 3642
rect 4010 3638 4013 3642
rect 5139 3638 5142 3642
rect 445 3618 446 3622
rect 557 3618 558 3622
rect 858 3618 873 3621
rect 1028 3618 1030 3622
rect 1186 3618 1190 3622
rect 1242 3618 1243 3622
rect 2290 3618 2291 3622
rect 2677 3618 2678 3622
rect 2724 3618 2726 3622
rect 4389 3618 4390 3622
rect 344 3603 346 3607
rect 350 3603 353 3607
rect 357 3603 360 3607
rect 1368 3603 1370 3607
rect 1374 3603 1377 3607
rect 1381 3603 1384 3607
rect 2392 3603 2394 3607
rect 2398 3603 2401 3607
rect 2405 3603 2408 3607
rect 3416 3603 3418 3607
rect 3422 3603 3425 3607
rect 3429 3603 3432 3607
rect 4440 3603 4442 3607
rect 4446 3603 4449 3607
rect 4453 3603 4456 3607
rect 285 3588 286 3592
rect 626 3588 627 3592
rect 1220 3588 1222 3592
rect 4829 3588 4830 3592
rect 214 3568 241 3571
rect 258 3568 265 3571
rect 678 3568 686 3571
rect 1322 3568 1345 3571
rect 1502 3568 1513 3571
rect 1517 3568 1518 3572
rect 1742 3568 1758 3571
rect 2622 3568 2630 3571
rect 2646 3568 2657 3571
rect 3226 3568 3229 3572
rect 670 3566 674 3568
rect 1502 3566 1506 3568
rect 1742 3566 1746 3568
rect 54 3558 65 3561
rect 98 3558 105 3561
rect 182 3558 193 3561
rect 214 3561 218 3564
rect 2654 3562 2657 3568
rect 214 3558 222 3561
rect 262 3558 273 3561
rect 590 3558 601 3561
rect 22 3548 38 3551
rect 118 3551 121 3558
rect 110 3548 121 3551
rect 198 3551 201 3558
rect 190 3548 201 3551
rect 350 3548 377 3551
rect 26 3538 33 3541
rect 54 3538 57 3548
rect 374 3542 377 3548
rect 418 3548 425 3551
rect 670 3551 673 3561
rect 702 3558 713 3561
rect 1462 3558 1470 3561
rect 1690 3558 1697 3561
rect 1890 3558 1897 3561
rect 2246 3558 2254 3561
rect 3006 3558 3017 3561
rect 654 3548 673 3551
rect 714 3548 721 3551
rect 814 3548 822 3551
rect 854 3548 878 3551
rect 902 3548 910 3551
rect 1142 3548 1150 3551
rect 1166 3551 1169 3558
rect 1166 3548 1177 3551
rect 1250 3548 1257 3551
rect 1262 3548 1278 3551
rect 1542 3548 1553 3551
rect 62 3538 81 3541
rect 398 3541 401 3548
rect 382 3538 401 3541
rect 470 3541 473 3548
rect 1550 3542 1553 3548
rect 1574 3542 1577 3551
rect 1614 3542 1617 3551
rect 1774 3548 1782 3551
rect 1946 3548 1969 3551
rect 2062 3548 2073 3551
rect 2358 3548 2366 3551
rect 2494 3551 2497 3558
rect 3748 3557 3750 3561
rect 3898 3557 3900 3561
rect 4222 3558 4230 3561
rect 4614 3558 4625 3561
rect 4702 3558 4710 3561
rect 5118 3558 5126 3561
rect 5278 3558 5286 3561
rect 2478 3548 2497 3551
rect 2558 3548 2574 3551
rect 2582 3548 2590 3551
rect 2686 3551 2690 3554
rect 2686 3548 2694 3551
rect 3082 3548 3089 3551
rect 3162 3548 3169 3551
rect 462 3538 473 3541
rect 690 3538 697 3541
rect 794 3538 801 3541
rect 806 3538 822 3541
rect 862 3538 905 3541
rect 974 3538 985 3541
rect 1094 3538 1102 3541
rect 1242 3538 1249 3541
rect 1662 3541 1665 3548
rect 2070 3542 2073 3548
rect 3306 3548 3313 3551
rect 3342 3548 3350 3551
rect 3382 3548 3398 3551
rect 3602 3548 3609 3551
rect 3722 3548 3737 3551
rect 3762 3548 3785 3551
rect 3910 3548 3950 3551
rect 4046 3551 4050 3553
rect 4010 3548 4017 3551
rect 4046 3548 4065 3551
rect 4134 3548 4145 3551
rect 4366 3551 4370 3554
rect 4614 3552 4617 3558
rect 4350 3548 4370 3551
rect 4398 3548 4409 3551
rect 4470 3548 4481 3551
rect 4550 3548 4558 3551
rect 4594 3548 4601 3551
rect 4694 3551 4697 3558
rect 4674 3548 4681 3551
rect 4686 3548 4697 3551
rect 4778 3548 4785 3551
rect 4806 3548 4817 3551
rect 4886 3548 4913 3551
rect 4942 3548 4950 3551
rect 5054 3548 5062 3551
rect 5222 3551 5226 3553
rect 4398 3542 4401 3548
rect 1662 3538 1673 3541
rect 1758 3538 1772 3541
rect 2030 3538 2041 3541
rect 2490 3538 2505 3541
rect 2670 3538 2681 3541
rect 2716 3538 2718 3542
rect 2834 3538 2841 3541
rect 2846 3538 2854 3541
rect 2914 3538 2937 3541
rect 2978 3538 2985 3541
rect 3022 3538 3030 3541
rect 3062 3538 3070 3541
rect 3154 3538 3169 3541
rect 3382 3538 3414 3541
rect 3770 3538 3785 3541
rect 3826 3538 3833 3541
rect 4058 3538 4065 3541
rect 4214 3538 4225 3541
rect 4426 3538 4433 3541
rect 4438 3538 4446 3541
rect 4550 3538 4553 3548
rect 4562 3538 4569 3541
rect 4598 3538 4601 3548
rect 4806 3542 4809 3548
rect 4886 3546 4890 3548
rect 5222 3548 5233 3551
rect 4606 3538 4614 3541
rect 4934 3538 4942 3541
rect 5054 3538 5089 3541
rect 694 3528 697 3538
rect 1742 3532 1745 3538
rect 782 3528 793 3531
rect 1106 3528 1110 3532
rect 1630 3528 1641 3531
rect 1738 3528 1745 3532
rect 1758 3532 1761 3538
rect 1830 3528 1838 3531
rect 2382 3528 2390 3531
rect 2630 3528 2633 3538
rect 2678 3532 2681 3538
rect 2794 3528 2809 3531
rect 3022 3528 3025 3538
rect 3621 3528 3622 3532
rect 3662 3528 3670 3531
rect 4894 3528 4897 3538
rect 5074 3528 5081 3531
rect 508 3518 510 3522
rect 1318 3518 1326 3521
rect 1382 3518 1390 3521
rect 1786 3518 1807 3521
rect 2138 3518 2139 3522
rect 2162 3518 2169 3521
rect 2765 3518 2766 3522
rect 2892 3518 2894 3522
rect 3042 3518 3043 3522
rect 4922 3518 4923 3522
rect 4996 3518 4998 3522
rect 5290 3518 5297 3521
rect 856 3503 858 3507
rect 862 3503 865 3507
rect 869 3503 872 3507
rect 1872 3503 1874 3507
rect 1878 3503 1881 3507
rect 1885 3503 1888 3507
rect 2904 3503 2906 3507
rect 2910 3503 2913 3507
rect 2917 3503 2920 3507
rect 3928 3503 3930 3507
rect 3934 3503 3937 3507
rect 3941 3503 3944 3507
rect 4952 3503 4954 3507
rect 4958 3503 4961 3507
rect 4965 3503 4968 3507
rect 36 3488 38 3492
rect 498 3488 505 3491
rect 722 3488 724 3492
rect 854 3488 862 3491
rect 1058 3488 1059 3492
rect 1218 3488 1220 3492
rect 1284 3488 1286 3492
rect 1636 3488 1638 3492
rect 2060 3488 2062 3492
rect 2162 3488 2164 3492
rect 2260 3488 2262 3492
rect 2820 3488 2822 3492
rect 626 3478 633 3482
rect 1402 3478 1406 3482
rect 1482 3478 1489 3482
rect 1858 3478 1862 3482
rect 3086 3478 3097 3481
rect 4174 3481 4177 3488
rect 4166 3478 4177 3481
rect 4474 3478 4478 3482
rect 4582 3478 4601 3481
rect 630 3472 633 3478
rect 1486 3472 1489 3478
rect 86 3468 94 3471
rect 154 3468 161 3471
rect 382 3468 393 3471
rect 450 3468 457 3471
rect 470 3468 478 3471
rect 542 3468 553 3471
rect 642 3468 649 3471
rect 782 3468 790 3471
rect 866 3468 881 3471
rect 1090 3468 1097 3471
rect 1306 3468 1313 3471
rect 1462 3468 1473 3471
rect 1578 3468 1585 3471
rect 1590 3468 1601 3471
rect 1654 3468 1662 3471
rect 1690 3468 1705 3471
rect 1774 3468 1785 3471
rect 550 3462 553 3468
rect 1462 3462 1465 3468
rect 1598 3462 1601 3468
rect 26 3458 33 3461
rect 322 3458 369 3461
rect 558 3458 569 3461
rect 606 3458 614 3461
rect 774 3458 790 3461
rect 798 3458 817 3461
rect 858 3458 889 3461
rect 894 3458 913 3461
rect 982 3458 1006 3461
rect 1854 3461 1857 3468
rect 1934 3468 1953 3471
rect 1970 3468 1977 3471
rect 2094 3468 2102 3471
rect 2190 3468 2201 3471
rect 2374 3468 2390 3471
rect 1838 3458 1857 3461
rect 1950 3458 1953 3468
rect 2454 3461 2457 3471
rect 2486 3468 2494 3471
rect 2970 3468 2977 3471
rect 2994 3468 3001 3471
rect 3278 3468 3290 3471
rect 4046 3468 4054 3471
rect 2454 3458 2462 3461
rect 2610 3458 2617 3461
rect 2862 3458 2878 3461
rect 2886 3458 2894 3461
rect 2950 3458 2958 3461
rect 3318 3458 3326 3461
rect 3822 3458 3830 3461
rect 4122 3458 4129 3461
rect 4194 3458 4201 3461
rect 4254 3461 4257 3471
rect 4262 3468 4273 3471
rect 4378 3468 4385 3471
rect 4242 3458 4257 3461
rect 4270 3462 4273 3468
rect 4758 3462 4761 3471
rect 4374 3458 4382 3461
rect 4622 3458 4641 3461
rect 4802 3458 4817 3461
rect 4838 3461 4841 3471
rect 4926 3468 4934 3471
rect 4946 3468 4953 3471
rect 5038 3468 5073 3471
rect 4826 3458 4841 3461
rect 4846 3458 4854 3461
rect 5038 3458 5062 3461
rect 5206 3458 5217 3461
rect 566 3452 569 3458
rect 814 3452 817 3458
rect 190 3448 201 3451
rect 270 3448 278 3451
rect 382 3448 390 3451
rect 1506 3448 1510 3452
rect 1814 3451 1817 3458
rect 1814 3448 1825 3451
rect 1854 3448 1857 3458
rect 2494 3451 2497 3458
rect 5206 3457 5210 3458
rect 2494 3448 2505 3451
rect 2598 3448 2609 3451
rect 4254 3448 4265 3451
rect 5102 3448 5110 3451
rect 174 3438 182 3441
rect 526 3438 534 3441
rect 1062 3441 1066 3444
rect 4254 3442 4257 3448
rect 1062 3438 1073 3441
rect 1554 3438 1558 3442
rect 1806 3438 1814 3441
rect 4438 3438 4454 3441
rect 4558 3438 4566 3441
rect 5187 3438 5190 3442
rect 1366 3428 1374 3431
rect 3046 3428 3049 3438
rect 1733 3418 1734 3422
rect 1957 3418 1958 3422
rect 2004 3418 2006 3422
rect 2349 3418 2350 3422
rect 2436 3418 2438 3422
rect 2764 3418 2766 3422
rect 2861 3418 2862 3422
rect 2949 3418 2950 3422
rect 4980 3418 4982 3422
rect 344 3403 346 3407
rect 350 3403 353 3407
rect 357 3403 360 3407
rect 1368 3403 1370 3407
rect 1374 3403 1377 3407
rect 1381 3403 1384 3407
rect 2392 3403 2394 3407
rect 2398 3403 2401 3407
rect 2405 3403 2408 3407
rect 3416 3403 3418 3407
rect 3422 3403 3425 3407
rect 3429 3403 3432 3407
rect 4440 3403 4442 3407
rect 4446 3403 4449 3407
rect 4453 3403 4456 3407
rect 852 3388 854 3392
rect 3402 3388 3404 3392
rect 5110 3372 5113 3381
rect 158 3368 166 3371
rect 629 3368 630 3372
rect 790 3368 801 3371
rect 998 3368 1009 3371
rect 1086 3368 1097 3371
rect 2150 3368 2158 3371
rect 2812 3368 2814 3372
rect 2962 3368 2977 3371
rect 3486 3368 3497 3371
rect 3548 3368 3550 3372
rect 3594 3368 3597 3372
rect 3970 3368 3977 3371
rect 4842 3368 4843 3372
rect 78 3361 81 3368
rect 798 3362 801 3368
rect 1006 3362 1009 3368
rect 1094 3362 1097 3368
rect 78 3358 89 3361
rect 606 3358 617 3361
rect 945 3358 953 3362
rect 990 3358 1001 3361
rect 1026 3358 1030 3362
rect 1174 3358 1185 3361
rect 1206 3358 1217 3361
rect 1502 3358 1510 3361
rect 1774 3361 1777 3368
rect 1766 3358 1777 3361
rect 1806 3358 1817 3361
rect 1854 3358 1865 3361
rect 10 3348 17 3351
rect 22 3348 30 3351
rect 34 3348 41 3351
rect 118 3351 122 3354
rect 114 3348 122 3351
rect 186 3348 193 3351
rect 26 3338 33 3341
rect 78 3338 89 3341
rect 334 3341 337 3351
rect 398 3348 406 3351
rect 334 3338 369 3341
rect 478 3341 481 3358
rect 950 3352 953 3358
rect 1862 3352 1865 3358
rect 590 3348 609 3351
rect 690 3348 697 3351
rect 1398 3348 1422 3351
rect 1494 3348 1502 3351
rect 1758 3348 1769 3351
rect 1778 3348 1793 3351
rect 2030 3351 2033 3361
rect 2118 3358 2126 3361
rect 2318 3361 2321 3368
rect 3486 3366 3490 3368
rect 2974 3362 2978 3364
rect 2302 3358 2321 3361
rect 2382 3358 2409 3361
rect 3126 3358 3134 3361
rect 2014 3348 2033 3351
rect 2070 3348 2078 3351
rect 2254 3348 2265 3351
rect 2702 3348 2713 3351
rect 3158 3348 3177 3351
rect 3250 3348 3257 3351
rect 3674 3348 3681 3351
rect 4342 3351 4346 3353
rect 4222 3348 4233 3351
rect 470 3338 481 3341
rect 498 3340 505 3341
rect 494 3338 505 3340
rect 590 3338 593 3348
rect 754 3338 761 3341
rect 1122 3338 1129 3341
rect 1294 3338 1302 3341
rect 1422 3338 1430 3341
rect 1438 3338 1454 3341
rect 1542 3341 1545 3348
rect 1518 3338 1529 3341
rect 1534 3338 1545 3341
rect 1594 3338 1609 3341
rect 2254 3338 2257 3348
rect 2702 3342 2705 3348
rect 4342 3348 4353 3351
rect 4422 3351 4425 3361
rect 4898 3358 4905 3361
rect 4394 3348 4409 3351
rect 4422 3348 4457 3351
rect 4646 3348 4654 3351
rect 4910 3351 4913 3358
rect 4910 3348 4921 3351
rect 5030 3348 5049 3351
rect 4350 3342 4353 3348
rect 2498 3338 2505 3341
rect 2546 3338 2553 3341
rect 2670 3338 2678 3341
rect 2950 3338 2961 3341
rect 2994 3338 3001 3341
rect 3078 3338 3094 3341
rect 3110 3338 3129 3341
rect 3454 3338 3473 3341
rect 3478 3338 3486 3341
rect 3510 3338 3521 3341
rect 3858 3338 3873 3341
rect 4370 3338 4377 3341
rect 4606 3338 4622 3341
rect 4926 3338 4961 3341
rect 4974 3338 5001 3341
rect 5086 3338 5094 3341
rect 5302 3338 5310 3341
rect 814 3332 817 3338
rect 990 3332 993 3338
rect 374 3328 385 3331
rect 482 3328 486 3332
rect 810 3328 817 3332
rect 986 3328 993 3332
rect 1294 3328 1297 3338
rect 1430 3328 1433 3338
rect 3510 3332 3513 3338
rect 2186 3328 2190 3332
rect 2370 3328 2377 3331
rect 2534 3328 2545 3331
rect 3018 3328 3025 3331
rect 3238 3328 3246 3331
rect 4366 3328 4369 3338
rect 4422 3328 4430 3331
rect 4958 3328 4961 3338
rect 69 3318 70 3322
rect 140 3318 142 3322
rect 226 3318 247 3321
rect 1332 3318 1334 3322
rect 1684 3318 1686 3322
rect 1980 3318 1982 3322
rect 2037 3318 2038 3322
rect 2236 3318 2238 3322
rect 2394 3318 2409 3321
rect 2458 3318 2460 3322
rect 2932 3318 2934 3322
rect 3286 3318 3294 3321
rect 5266 3318 5267 3322
rect 856 3303 858 3307
rect 862 3303 865 3307
rect 869 3303 872 3307
rect 1872 3303 1874 3307
rect 1878 3303 1881 3307
rect 1885 3303 1888 3307
rect 2904 3303 2906 3307
rect 2910 3303 2913 3307
rect 2917 3303 2920 3307
rect 3928 3303 3930 3307
rect 3934 3303 3937 3307
rect 3941 3303 3944 3307
rect 4952 3303 4954 3307
rect 4958 3303 4961 3307
rect 4965 3303 4968 3307
rect 342 3288 358 3291
rect 644 3288 646 3292
rect 797 3288 798 3292
rect 940 3288 942 3292
rect 1132 3288 1134 3292
rect 1348 3288 1350 3292
rect 2170 3288 2171 3292
rect 2982 3288 2998 3291
rect 3406 3288 3422 3291
rect 4364 3288 4366 3292
rect 4930 3288 4931 3292
rect 5053 3288 5054 3292
rect 850 3278 862 3281
rect 2170 3278 2185 3281
rect 22 3258 38 3261
rect 138 3258 145 3261
rect 150 3258 166 3261
rect 214 3261 217 3271
rect 354 3268 369 3271
rect 574 3271 577 3278
rect 574 3268 585 3271
rect 606 3268 614 3271
rect 710 3268 721 3271
rect 1078 3271 1081 3278
rect 1070 3268 1081 3271
rect 1086 3268 1105 3271
rect 1310 3268 1321 3271
rect 1510 3268 1521 3271
rect 1558 3268 1569 3271
rect 1586 3268 1593 3271
rect 1654 3268 1662 3271
rect 2014 3268 2025 3271
rect 2150 3268 2161 3271
rect 2190 3268 2201 3271
rect 2206 3268 2222 3271
rect 2242 3268 2249 3271
rect 2434 3268 2441 3271
rect 2470 3268 2489 3271
rect 2558 3271 2561 3281
rect 2910 3278 2926 3281
rect 3242 3278 3254 3281
rect 3270 3278 3281 3281
rect 2518 3268 2545 3271
rect 2558 3268 2566 3271
rect 2574 3268 2582 3271
rect 2726 3271 2729 3278
rect 2714 3268 2721 3271
rect 2726 3268 2737 3271
rect 2742 3268 2761 3271
rect 198 3258 217 3261
rect 466 3258 481 3261
rect 526 3258 558 3261
rect 686 3258 705 3261
rect 758 3258 790 3261
rect 902 3258 905 3268
rect 1190 3258 1222 3261
rect 1446 3261 1449 3268
rect 1566 3262 1569 3268
rect 1422 3258 1449 3261
rect 1662 3258 1673 3261
rect 1678 3258 1697 3261
rect 1822 3258 1838 3261
rect 2070 3258 2089 3261
rect 2278 3258 2286 3261
rect 2430 3258 2446 3261
rect 2662 3258 2678 3261
rect 2902 3258 2937 3261
rect 3030 3261 3033 3271
rect 3092 3268 3094 3272
rect 3126 3268 3137 3271
rect 3030 3258 3065 3261
rect 3230 3261 3233 3271
rect 3418 3268 3433 3271
rect 3742 3268 3777 3271
rect 3990 3271 3993 3281
rect 4562 3278 4569 3281
rect 4942 3272 4945 3281
rect 4950 3278 4958 3281
rect 5022 3272 5025 3281
rect 5030 3278 5038 3281
rect 3974 3268 3993 3271
rect 4006 3268 4025 3271
rect 4134 3268 4146 3271
rect 3222 3258 3233 3261
rect 3250 3258 3257 3261
rect 3498 3258 3505 3261
rect 3954 3258 3961 3261
rect 4006 3258 4009 3268
rect 4390 3262 4393 3271
rect 4682 3268 4689 3271
rect 4694 3268 4721 3271
rect 4878 3268 4886 3271
rect 5002 3268 5009 3271
rect 4466 3258 4473 3261
rect 4478 3258 4497 3261
rect 4518 3258 4529 3261
rect 4814 3258 4825 3261
rect 4998 3258 5017 3261
rect 5038 3258 5046 3261
rect 5134 3261 5137 3281
rect 5142 3268 5150 3271
rect 5122 3258 5137 3261
rect 102 3251 105 3258
rect 94 3248 105 3251
rect 674 3248 681 3251
rect 686 3248 689 3258
rect 1162 3248 1169 3251
rect 1510 3251 1513 3258
rect 1502 3248 1513 3251
rect 1582 3251 1585 3258
rect 1574 3248 1585 3251
rect 1662 3252 1665 3258
rect 1694 3252 1697 3258
rect 1710 3248 1726 3251
rect 1964 3248 1966 3252
rect 2002 3248 2006 3252
rect 2014 3248 2022 3251
rect 2086 3248 2089 3258
rect 2134 3248 2142 3251
rect 2262 3248 2281 3251
rect 2390 3248 2406 3251
rect 2462 3248 2473 3251
rect 2790 3251 2793 3258
rect 2774 3248 2793 3251
rect 2934 3251 2937 3258
rect 3222 3256 3226 3258
rect 2930 3248 2937 3251
rect 3406 3248 3422 3251
rect 3474 3248 3478 3252
rect 4998 3248 5001 3258
rect 694 3242 698 3244
rect 244 3238 246 3242
rect 342 3238 358 3241
rect 1494 3241 1498 3244
rect 2086 3242 2090 3244
rect 1486 3238 1498 3241
rect 1620 3238 1622 3242
rect 1868 3238 1870 3242
rect 4420 3238 4422 3242
rect 18 3218 19 3222
rect 170 3218 171 3222
rect 2301 3218 2302 3222
rect 2690 3218 2691 3222
rect 2813 3218 2814 3222
rect 3340 3218 3342 3222
rect 5277 3218 5278 3222
rect 344 3203 346 3207
rect 350 3203 353 3207
rect 357 3203 360 3207
rect 1368 3203 1370 3207
rect 1374 3203 1377 3207
rect 1381 3203 1384 3207
rect 2392 3203 2394 3207
rect 2398 3203 2401 3207
rect 2405 3203 2408 3207
rect 3416 3203 3418 3207
rect 3422 3203 3425 3207
rect 3429 3203 3432 3207
rect 4440 3203 4442 3207
rect 4446 3203 4449 3207
rect 4453 3203 4456 3207
rect 290 3188 291 3192
rect 738 3188 740 3192
rect 866 3188 873 3191
rect 2442 3188 2444 3192
rect 3173 3188 3174 3192
rect 4042 3188 4044 3192
rect 4468 3188 4470 3192
rect 38 3172 41 3181
rect 950 3168 958 3171
rect 1206 3168 1214 3171
rect 1286 3168 1294 3171
rect 3574 3168 3585 3171
rect 4835 3168 4838 3172
rect 314 3158 321 3161
rect 454 3161 457 3168
rect 3574 3162 3577 3168
rect 438 3158 457 3161
rect 482 3158 489 3161
rect 1454 3158 1465 3161
rect 382 3151 386 3154
rect 1462 3152 1466 3154
rect 382 3148 393 3151
rect 662 3148 697 3151
rect 1134 3148 1145 3151
rect 1218 3148 1225 3151
rect 1394 3148 1401 3151
rect 1534 3151 1537 3161
rect 1746 3158 1753 3161
rect 1937 3158 1945 3162
rect 1942 3152 1945 3158
rect 1526 3148 1537 3151
rect 1554 3148 1593 3151
rect 1702 3148 1713 3151
rect 194 3138 201 3141
rect 218 3138 225 3141
rect 494 3138 502 3141
rect 526 3141 529 3148
rect 1526 3142 1529 3148
rect 1710 3142 1713 3148
rect 2302 3151 2305 3161
rect 2322 3158 2329 3161
rect 2286 3148 2305 3151
rect 2342 3148 2358 3151
rect 2526 3148 2534 3151
rect 2582 3148 2622 3151
rect 2646 3151 2650 3154
rect 2702 3152 2705 3161
rect 2734 3158 2742 3161
rect 3129 3158 3137 3162
rect 3134 3152 3137 3158
rect 2630 3148 2650 3151
rect 2686 3148 2702 3151
rect 3206 3151 3209 3161
rect 3270 3158 3281 3161
rect 3206 3148 3225 3151
rect 3282 3148 3289 3151
rect 3342 3151 3345 3161
rect 3414 3158 3422 3161
rect 3462 3158 3470 3161
rect 3478 3158 3489 3161
rect 3486 3152 3490 3154
rect 3334 3148 3345 3151
rect 3454 3148 3462 3151
rect 3542 3151 3545 3161
rect 3562 3158 3569 3161
rect 3526 3148 3545 3151
rect 3658 3148 3665 3151
rect 518 3138 529 3141
rect 702 3138 721 3141
rect 1378 3138 1393 3141
rect 1410 3138 1417 3141
rect 1514 3138 1521 3141
rect 1558 3138 1569 3141
rect 1626 3138 1633 3141
rect 1654 3138 1665 3141
rect 1766 3141 1769 3148
rect 1766 3138 1777 3141
rect 1806 3141 1809 3148
rect 3334 3146 3338 3148
rect 3946 3148 3953 3151
rect 4626 3148 4633 3151
rect 4894 3148 4918 3151
rect 5118 3148 5126 3151
rect 5138 3148 5161 3151
rect 1786 3138 1793 3141
rect 1798 3138 1809 3141
rect 2070 3138 2081 3141
rect 2098 3138 2105 3141
rect 2166 3138 2185 3141
rect 2270 3138 2281 3141
rect 2322 3138 2329 3141
rect 2402 3138 2425 3141
rect 2470 3138 2489 3141
rect 2610 3138 2617 3141
rect 2718 3138 2737 3141
rect 2830 3138 2849 3141
rect 3014 3138 3025 3141
rect 3222 3138 3238 3141
rect 3254 3138 3273 3141
rect 3362 3138 3377 3141
rect 3622 3138 3641 3141
rect 3650 3138 3657 3141
rect 4242 3138 4249 3141
rect 334 3128 342 3131
rect 1276 3128 1278 3132
rect 1310 3128 1321 3131
rect 1566 3131 1569 3138
rect 2078 3132 2081 3138
rect 1566 3128 1577 3131
rect 1582 3128 1590 3131
rect 2358 3131 2361 3138
rect 2358 3128 2369 3131
rect 3574 3128 3593 3131
rect 3654 3128 3657 3138
rect 4694 3132 4697 3142
rect 4894 3138 4921 3141
rect 5118 3138 5153 3141
rect 4918 3132 4921 3138
rect 4946 3128 4953 3131
rect 172 3118 174 3122
rect 612 3118 614 3122
rect 828 3118 830 3122
rect 1036 3118 1038 3122
rect 1092 3118 1094 3122
rect 1254 3118 1262 3121
rect 1834 3118 1836 3122
rect 1996 3118 1998 3122
rect 2042 3118 2044 3122
rect 2122 3118 2124 3122
rect 2212 3118 2214 3122
rect 2866 3118 2868 3122
rect 2948 3118 2950 3122
rect 4514 3118 4516 3122
rect 5169 3118 5182 3121
rect 5294 3118 5302 3121
rect 856 3103 858 3107
rect 862 3103 865 3107
rect 869 3103 872 3107
rect 1872 3103 1874 3107
rect 1878 3103 1881 3107
rect 1885 3103 1888 3107
rect 2904 3103 2906 3107
rect 2910 3103 2913 3107
rect 2917 3103 2920 3107
rect 3928 3103 3930 3107
rect 3934 3103 3937 3107
rect 3941 3103 3944 3107
rect 4952 3103 4954 3107
rect 4958 3103 4961 3107
rect 4965 3103 4968 3107
rect 332 3088 334 3092
rect 541 3088 542 3092
rect 578 3088 580 3092
rect 882 3088 883 3092
rect 1082 3088 1084 3092
rect 1206 3088 1214 3091
rect 1526 3088 1534 3091
rect 1650 3088 1651 3092
rect 2445 3088 2446 3092
rect 2878 3088 2894 3091
rect 3820 3088 3822 3092
rect 3876 3088 3878 3092
rect 4220 3088 4222 3092
rect 4572 3088 4574 3092
rect 4788 3088 4790 3092
rect 4908 3088 4910 3092
rect 130 3078 145 3081
rect 108 3068 121 3071
rect 502 3068 534 3071
rect 662 3068 670 3071
rect 766 3071 769 3081
rect 2126 3072 2129 3081
rect 2154 3078 2169 3081
rect 2238 3078 2257 3081
rect 3452 3078 3454 3082
rect 766 3068 774 3071
rect 838 3068 873 3071
rect 990 3062 993 3071
rect 1166 3068 1174 3071
rect 1222 3068 1233 3071
rect 1306 3068 1313 3071
rect 1318 3068 1345 3071
rect 1482 3068 1489 3071
rect 26 3058 33 3061
rect 166 3058 174 3061
rect 390 3058 398 3061
rect 426 3058 433 3061
rect 638 3058 662 3061
rect 958 3058 966 3061
rect 1038 3061 1041 3068
rect 1602 3068 1609 3071
rect 1630 3068 1641 3071
rect 2086 3068 2094 3071
rect 2134 3068 2145 3071
rect 2174 3068 2182 3071
rect 2190 3068 2209 3071
rect 2390 3068 2417 3071
rect 2458 3068 2465 3071
rect 2566 3068 2574 3071
rect 2622 3068 2633 3071
rect 2670 3068 2689 3071
rect 2822 3068 2841 3071
rect 3054 3068 3073 3071
rect 3238 3068 3249 3071
rect 3370 3068 3377 3071
rect 3654 3071 3657 3081
rect 4374 3078 4393 3081
rect 3638 3068 3657 3071
rect 3702 3068 3710 3071
rect 3730 3068 3737 3071
rect 1030 3058 1041 3061
rect 1278 3058 1286 3061
rect 1294 3058 1313 3061
rect 1330 3058 1337 3061
rect 1574 3058 1614 3061
rect 2078 3058 2102 3061
rect 2422 3058 2441 3061
rect 2542 3058 2574 3061
rect 2646 3058 2665 3061
rect 2986 3058 2993 3061
rect 3030 3058 3049 3061
rect 3098 3058 3105 3061
rect 3506 3058 3513 3061
rect 3534 3058 3537 3068
rect 4518 3071 4521 3081
rect 4502 3068 4521 3071
rect 4650 3068 4651 3072
rect 4750 3068 4761 3071
rect 4806 3068 4825 3071
rect 4862 3068 4881 3071
rect 4926 3068 4942 3071
rect 4982 3068 4990 3071
rect 3754 3058 3761 3061
rect 3922 3058 3929 3061
rect 4134 3058 4150 3061
rect 4166 3061 4169 3068
rect 4166 3058 4177 3061
rect 4358 3058 4366 3061
rect 4382 3058 4390 3061
rect 4702 3058 4721 3061
rect 4734 3058 4753 3061
rect 4850 3058 4865 3061
rect 4982 3058 5006 3061
rect 5210 3058 5217 3061
rect 1310 3052 1313 3058
rect 890 3048 897 3051
rect 1022 3048 1033 3051
rect 1242 3048 1246 3052
rect 1286 3048 1297 3051
rect 2106 3048 2110 3052
rect 2118 3048 2137 3051
rect 2438 3048 2441 3058
rect 2646 3048 2649 3058
rect 2686 3048 2694 3051
rect 3030 3048 3033 3058
rect 3185 3048 3190 3052
rect 3342 3048 3353 3051
rect 3350 3042 3353 3048
rect 3470 3048 3481 3051
rect 3490 3048 3494 3052
rect 4042 3048 4049 3051
rect 4734 3048 4737 3058
rect 4830 3051 4833 3058
rect 4830 3048 4841 3051
rect 98 3038 105 3041
rect 757 3038 758 3042
rect 1206 3038 1214 3041
rect 2258 3038 2265 3041
rect 2804 3038 2806 3042
rect 3366 3041 3369 3048
rect 3358 3038 3369 3041
rect 3462 3041 3465 3048
rect 3550 3046 3554 3048
rect 3462 3038 3473 3041
rect 3550 3038 3577 3041
rect 4310 3038 4334 3041
rect 1866 3018 1867 3022
rect 2077 3018 2078 3022
rect 2242 3018 2243 3022
rect 2290 3018 2292 3022
rect 2932 3018 2934 3022
rect 3306 3018 3307 3022
rect 3330 3018 3331 3022
rect 344 3003 346 3007
rect 350 3003 353 3007
rect 357 3003 360 3007
rect 1368 3003 1370 3007
rect 1374 3003 1377 3007
rect 1381 3003 1384 3007
rect 2392 3003 2394 3007
rect 2398 3003 2401 3007
rect 2405 3003 2408 3007
rect 3416 3003 3418 3007
rect 3422 3003 3425 3007
rect 3429 3003 3432 3007
rect 4440 3003 4442 3007
rect 4446 3003 4449 3007
rect 4453 3003 4456 3007
rect 410 2988 411 2992
rect 514 2988 516 2992
rect 578 2988 579 2992
rect 1122 2988 1123 2992
rect 2709 2988 2710 2992
rect 2837 2988 2838 2992
rect 2972 2988 2974 2992
rect 3205 2988 3206 2992
rect 3837 2988 3838 2992
rect 3874 2988 3876 2992
rect 4186 2988 4190 2992
rect 4276 2988 4278 2992
rect 4380 2988 4382 2992
rect 3526 2972 3529 2981
rect 38 2968 54 2971
rect 86 2968 113 2971
rect 770 2968 771 2972
rect 1170 2968 1177 2971
rect 2090 2968 2091 2972
rect 2246 2968 2265 2971
rect 2564 2968 2566 2972
rect 3234 2968 3241 2971
rect 3334 2968 3345 2971
rect 4506 2968 4513 2971
rect 54 2958 65 2961
rect 86 2961 90 2964
rect 86 2958 94 2961
rect 170 2958 177 2961
rect 186 2958 190 2962
rect 318 2958 329 2961
rect 70 2951 73 2958
rect 62 2948 73 2951
rect 122 2948 137 2951
rect 282 2948 297 2951
rect 330 2948 337 2951
rect 446 2951 449 2961
rect 1202 2958 1209 2961
rect 1566 2958 1574 2961
rect 1790 2961 1793 2968
rect 1782 2958 1793 2961
rect 1866 2958 1889 2961
rect 2126 2958 2134 2961
rect 394 2948 409 2951
rect 446 2948 465 2951
rect 722 2948 729 2951
rect 1150 2948 1161 2951
rect 1190 2948 1206 2951
rect 1158 2942 1161 2948
rect 1514 2948 1529 2951
rect 1730 2948 1737 2951
rect 1830 2948 1838 2951
rect 2082 2948 2089 2951
rect 2166 2951 2170 2954
rect 2166 2948 2177 2951
rect 2262 2948 2265 2968
rect 2286 2961 2289 2968
rect 2278 2958 2289 2961
rect 2518 2958 2529 2961
rect 2686 2961 2689 2968
rect 3342 2962 3345 2968
rect 2670 2958 2689 2961
rect 2814 2958 2825 2961
rect 2862 2958 2873 2961
rect 3914 2958 3937 2961
rect 4430 2958 4438 2961
rect 5158 2958 5166 2961
rect 2526 2952 2529 2958
rect 2334 2948 2345 2951
rect 302 2938 321 2941
rect 350 2938 377 2941
rect 470 2938 481 2941
rect 686 2938 694 2941
rect 374 2932 377 2938
rect 934 2932 937 2942
rect 1174 2938 1185 2941
rect 1670 2938 1682 2941
rect 1782 2938 1793 2941
rect 1950 2941 1953 2948
rect 1974 2941 1977 2948
rect 1942 2938 1953 2941
rect 1966 2938 1977 2941
rect 2042 2938 2049 2941
rect 2074 2938 2081 2941
rect 2190 2938 2209 2941
rect 2230 2938 2238 2941
rect 2342 2938 2345 2948
rect 2838 2948 2854 2951
rect 3030 2948 3065 2951
rect 2530 2938 2537 2941
rect 2630 2941 2633 2948
rect 3062 2942 3065 2948
rect 2630 2938 2641 2941
rect 2778 2938 2785 2941
rect 2990 2938 3006 2941
rect 3086 2938 3097 2941
rect 3198 2941 3201 2951
rect 3398 2948 3422 2951
rect 3610 2948 3617 2951
rect 3642 2948 3649 2951
rect 3814 2948 3830 2951
rect 4078 2948 4086 2951
rect 4158 2948 4166 2951
rect 4738 2948 4745 2951
rect 3182 2938 3201 2941
rect 3356 2938 3358 2942
rect 3546 2938 3553 2941
rect 3614 2938 3617 2948
rect 4878 2948 4886 2951
rect 4954 2948 4990 2951
rect 5022 2948 5038 2951
rect 5094 2948 5126 2951
rect 4878 2946 4882 2948
rect 3658 2938 3665 2941
rect 3986 2938 3993 2941
rect 4162 2938 4169 2941
rect 4398 2938 4406 2941
rect 4458 2938 4465 2941
rect 4718 2938 4737 2941
rect 5094 2938 5129 2941
rect 1766 2931 1770 2933
rect 2670 2932 2673 2938
rect 3302 2932 3305 2938
rect 1766 2928 1774 2931
rect 2050 2928 2054 2932
rect 2150 2928 2161 2931
rect 2630 2928 2641 2931
rect 2666 2928 2673 2932
rect 3166 2928 3177 2931
rect 3298 2928 3305 2932
rect 3470 2931 3473 2938
rect 3470 2928 3481 2931
rect 3494 2928 3497 2938
rect 3630 2932 3633 2938
rect 3626 2928 3633 2932
rect 2158 2922 2161 2928
rect 4054 2928 4065 2931
rect 4070 2928 4078 2931
rect 4554 2928 4561 2931
rect 4734 2928 4737 2938
rect 4958 2928 4974 2931
rect 5010 2928 5011 2932
rect 1802 2918 1803 2922
rect 2362 2918 2364 2922
rect 3244 2918 3246 2922
rect 3437 2918 3438 2922
rect 3565 2918 3566 2922
rect 3708 2918 3710 2922
rect 4585 2918 4590 2922
rect 4902 2918 4910 2921
rect 856 2903 858 2907
rect 862 2903 865 2907
rect 869 2903 872 2907
rect 1872 2903 1874 2907
rect 1878 2903 1881 2907
rect 1885 2903 1888 2907
rect 2904 2903 2906 2907
rect 2910 2903 2913 2907
rect 2917 2903 2920 2907
rect 3928 2903 3930 2907
rect 3934 2903 3937 2907
rect 3941 2903 3944 2907
rect 4952 2903 4954 2907
rect 4958 2903 4961 2907
rect 4965 2903 4968 2907
rect 26 2888 28 2892
rect 314 2888 316 2892
rect 706 2888 708 2892
rect 762 2888 764 2892
rect 1509 2888 1510 2892
rect 3404 2888 3406 2892
rect 3572 2888 3574 2892
rect 3740 2888 3742 2892
rect 3981 2888 3982 2892
rect 4422 2888 4438 2891
rect 158 2878 169 2881
rect 1574 2878 1585 2881
rect 1782 2878 1790 2881
rect 1870 2878 1902 2881
rect 158 2872 161 2878
rect 134 2868 142 2871
rect 670 2868 689 2871
rect 802 2868 809 2871
rect 814 2868 822 2871
rect 1254 2868 1257 2878
rect 1494 2868 1502 2871
rect 1518 2868 1526 2871
rect 1546 2868 1553 2871
rect 1586 2868 1593 2871
rect 414 2858 430 2861
rect 626 2858 633 2861
rect 1542 2858 1558 2861
rect 1686 2858 1694 2861
rect 1758 2861 1761 2871
rect 1910 2868 1918 2871
rect 2078 2871 2081 2881
rect 2942 2878 2958 2881
rect 3138 2878 3145 2881
rect 2062 2868 2081 2871
rect 2278 2868 2286 2871
rect 2378 2868 2401 2871
rect 2438 2868 2449 2871
rect 2812 2868 2814 2872
rect 2886 2868 2910 2871
rect 3118 2871 3121 2878
rect 3110 2868 3121 2871
rect 3146 2868 3153 2871
rect 3158 2868 3180 2871
rect 3246 2868 3257 2871
rect 3318 2871 3321 2881
rect 3902 2878 3913 2881
rect 4010 2878 4017 2882
rect 4166 2878 4177 2881
rect 4014 2872 4017 2878
rect 3306 2868 3321 2871
rect 1730 2858 1761 2861
rect 1794 2858 1801 2861
rect 1938 2858 1945 2861
rect 2126 2861 2129 2868
rect 3254 2862 3257 2868
rect 2118 2858 2129 2861
rect 2270 2858 2294 2861
rect 2386 2858 2409 2861
rect 2590 2858 2630 2861
rect 2978 2858 2985 2861
rect 2990 2858 2998 2861
rect 3014 2858 3046 2861
rect 3326 2861 3329 2871
rect 3486 2868 3494 2871
rect 3298 2858 3329 2861
rect 3450 2858 3457 2861
rect 3590 2861 3593 2871
rect 3590 2858 3609 2861
rect 3666 2858 3673 2861
rect 3758 2861 3761 2871
rect 3790 2868 3798 2871
rect 3814 2862 3817 2871
rect 3838 2868 3857 2871
rect 3894 2868 3902 2871
rect 4150 2871 4153 2878
rect 4142 2868 4153 2871
rect 4158 2868 4166 2871
rect 4214 2871 4217 2881
rect 4794 2878 4801 2881
rect 4202 2868 4217 2871
rect 4294 2868 4305 2871
rect 3758 2858 3769 2861
rect 3958 2858 3966 2861
rect 4070 2858 4086 2861
rect 4194 2858 4233 2861
rect 4638 2858 4641 2868
rect 4822 2858 4841 2861
rect 4846 2858 4854 2861
rect 4870 2858 4897 2861
rect 5122 2858 5137 2861
rect 5226 2858 5233 2861
rect 1998 2848 2006 2851
rect 2422 2848 2430 2851
rect 2698 2848 2705 2851
rect 2782 2848 2790 2851
rect 3274 2848 3281 2851
rect 3638 2851 3641 2858
rect 3630 2848 3641 2851
rect 3806 2848 3817 2851
rect 4046 2848 4057 2851
rect 4094 2848 4105 2851
rect 4910 2848 4937 2851
rect 106 2838 108 2842
rect 1562 2838 1563 2842
rect 1574 2838 1582 2841
rect 2062 2838 2070 2841
rect 2634 2838 2635 2842
rect 2670 2838 2678 2841
rect 2794 2838 2801 2841
rect 4666 2838 4682 2841
rect 1610 2818 1611 2822
rect 4693 2818 4694 2822
rect 4725 2818 4726 2822
rect 4786 2818 4787 2822
rect 4898 2818 4899 2822
rect 344 2803 346 2807
rect 350 2803 353 2807
rect 357 2803 360 2807
rect 1368 2803 1370 2807
rect 1374 2803 1377 2807
rect 1381 2803 1384 2807
rect 2392 2803 2394 2807
rect 2398 2803 2401 2807
rect 2405 2803 2408 2807
rect 3416 2803 3418 2807
rect 3422 2803 3425 2807
rect 3429 2803 3432 2807
rect 4440 2803 4442 2807
rect 4446 2803 4449 2807
rect 4453 2803 4456 2807
rect 378 2788 379 2792
rect 821 2788 822 2792
rect 922 2788 924 2792
rect 1234 2788 1235 2792
rect 2053 2788 2054 2792
rect 3021 2788 3022 2792
rect 3469 2788 3470 2792
rect 94 2768 102 2771
rect 534 2768 542 2771
rect 766 2768 782 2771
rect 1627 2768 1630 2772
rect 1954 2768 1961 2771
rect 1982 2768 1990 2771
rect 2326 2768 2334 2771
rect 2870 2771 2873 2781
rect 2870 2768 2894 2771
rect 2922 2768 2953 2771
rect 3802 2768 3803 2772
rect 3970 2768 3977 2771
rect 4339 2768 4342 2772
rect 126 2748 134 2751
rect 186 2748 217 2751
rect 318 2751 321 2761
rect 798 2761 801 2768
rect 782 2758 801 2761
rect 1194 2758 1201 2761
rect 1706 2758 1713 2761
rect 1806 2758 1814 2761
rect 1982 2758 1993 2761
rect 2410 2758 2417 2761
rect 2794 2758 2801 2761
rect 2842 2758 2849 2761
rect 3278 2758 3286 2761
rect 3634 2758 3641 2761
rect 3850 2758 3857 2761
rect 310 2748 321 2751
rect 354 2748 377 2751
rect 582 2748 590 2751
rect 134 2738 142 2741
rect 182 2738 185 2748
rect 310 2742 313 2748
rect 746 2748 753 2751
rect 962 2748 969 2751
rect 1046 2748 1078 2751
rect 1122 2748 1145 2751
rect 1202 2748 1209 2751
rect 518 2738 526 2741
rect 1070 2738 1086 2741
rect 1158 2741 1161 2748
rect 1938 2748 1945 2751
rect 2030 2748 2049 2751
rect 2758 2748 2793 2751
rect 2966 2748 2974 2751
rect 3602 2748 3609 2751
rect 3614 2748 3630 2751
rect 3662 2748 3670 2751
rect 3830 2748 3838 2751
rect 3918 2748 3942 2751
rect 4094 2751 4097 2761
rect 4134 2758 4142 2761
rect 4438 2758 4446 2761
rect 5270 2758 5278 2761
rect 4094 2748 4113 2751
rect 2790 2742 2793 2748
rect 1150 2738 1161 2741
rect 1522 2738 1537 2741
rect 1678 2738 1689 2741
rect 1694 2738 1702 2741
rect 1842 2738 1849 2741
rect 2214 2738 2226 2741
rect 2830 2738 2833 2748
rect 4094 2742 4097 2748
rect 4422 2751 4426 2754
rect 4422 2748 4430 2751
rect 4470 2748 4494 2751
rect 4762 2748 4769 2751
rect 4838 2748 4857 2751
rect 4934 2748 4966 2751
rect 5106 2748 5113 2751
rect 3034 2738 3049 2741
rect 3180 2738 3182 2742
rect 3942 2738 3958 2741
rect 3986 2738 3993 2741
rect 4118 2738 4137 2741
rect 218 2728 233 2731
rect 1126 2728 1134 2731
rect 1862 2728 1873 2731
rect 2310 2731 2314 2733
rect 4230 2732 4233 2742
rect 4734 2738 4742 2741
rect 4806 2738 4814 2741
rect 2310 2728 2321 2731
rect 3214 2728 3225 2731
rect 854 2718 862 2721
rect 1717 2718 1718 2722
rect 2100 2718 2102 2722
rect 2658 2718 2660 2722
rect 3100 2718 3102 2722
rect 3372 2718 3374 2722
rect 3516 2718 3518 2722
rect 3572 2718 3574 2722
rect 3962 2718 3969 2721
rect 4458 2718 4465 2721
rect 4578 2718 4585 2721
rect 4614 2718 4622 2721
rect 4668 2718 4670 2722
rect 4725 2718 4726 2722
rect 856 2703 858 2707
rect 862 2703 865 2707
rect 869 2703 872 2707
rect 1872 2703 1874 2707
rect 1878 2703 1881 2707
rect 1885 2703 1888 2707
rect 2904 2703 2906 2707
rect 2910 2703 2913 2707
rect 2917 2703 2920 2707
rect 3928 2703 3930 2707
rect 3934 2703 3937 2707
rect 3941 2703 3944 2707
rect 4952 2703 4954 2707
rect 4958 2703 4961 2707
rect 4965 2703 4968 2707
rect 61 2688 62 2692
rect 562 2688 563 2692
rect 690 2688 692 2692
rect 770 2688 772 2692
rect 837 2688 838 2692
rect 858 2688 873 2691
rect 2050 2688 2052 2692
rect 2341 2688 2342 2692
rect 2402 2688 2409 2691
rect 2418 2688 2419 2692
rect 2602 2688 2604 2692
rect 2930 2688 2937 2691
rect 3138 2688 3139 2692
rect 3586 2688 3588 2692
rect 3934 2688 3950 2691
rect 4938 2688 4940 2692
rect 270 2678 281 2681
rect 414 2678 422 2682
rect 738 2678 742 2682
rect 1190 2678 1201 2681
rect 2110 2678 2121 2681
rect 2126 2678 2134 2681
rect 2282 2678 2286 2682
rect 2910 2678 2937 2681
rect 414 2672 417 2678
rect 38 2668 54 2671
rect 354 2668 369 2671
rect 618 2668 625 2671
rect 722 2668 729 2671
rect 746 2668 753 2671
rect 1054 2668 1062 2671
rect 1350 2668 1358 2671
rect 1958 2668 1966 2671
rect 2110 2671 2113 2678
rect 4086 2672 4089 2681
rect 4286 2678 4294 2682
rect 2010 2668 2017 2671
rect 2102 2668 2113 2671
rect 2198 2668 2209 2671
rect 2286 2668 2297 2671
rect 2350 2668 2361 2671
rect 2382 2668 2398 2671
rect 2630 2668 2649 2671
rect 2878 2668 2886 2671
rect 3146 2668 3161 2671
rect 3214 2668 3222 2671
rect 3270 2668 3281 2671
rect 3294 2668 3305 2671
rect 3326 2668 3334 2671
rect 3886 2668 3894 2671
rect 4262 2671 4265 2678
rect 4286 2672 4289 2678
rect 4262 2668 4273 2671
rect 4618 2668 4633 2671
rect 4826 2668 4833 2671
rect 4966 2668 4993 2671
rect 5146 2668 5153 2671
rect 94 2658 102 2661
rect 466 2658 473 2661
rect 558 2658 577 2661
rect 618 2658 633 2661
rect 1058 2658 1065 2661
rect 1166 2658 1177 2661
rect 1214 2658 1222 2661
rect 1430 2658 1438 2661
rect 1622 2658 1630 2661
rect 2286 2662 2289 2668
rect 2098 2658 2137 2661
rect 2310 2661 2313 2668
rect 2310 2658 2321 2661
rect 2550 2658 2558 2661
rect 2706 2658 2721 2661
rect 2810 2658 2817 2661
rect 2870 2658 2889 2661
rect 3294 2662 3297 2668
rect 3170 2658 3185 2661
rect 3322 2658 3337 2661
rect 3502 2658 3510 2661
rect 3882 2658 3897 2661
rect 4150 2661 4153 2668
rect 4106 2658 4113 2661
rect 4118 2658 4153 2661
rect 4302 2658 4313 2661
rect 4506 2658 4513 2661
rect 4818 2658 4841 2661
rect 4846 2658 4865 2661
rect 5138 2658 5161 2661
rect 5262 2658 5270 2661
rect 102 2648 113 2651
rect 482 2648 489 2651
rect 574 2648 577 2658
rect 982 2656 986 2658
rect 982 2648 993 2651
rect 1002 2648 1009 2651
rect 1150 2648 1169 2651
rect 1366 2648 1374 2651
rect 2074 2648 2081 2651
rect 3278 2651 3281 2658
rect 3270 2648 3281 2651
rect 3814 2648 3822 2651
rect 3838 2651 3841 2658
rect 4302 2652 4305 2658
rect 3830 2648 3841 2651
rect 4094 2648 4105 2651
rect 4194 2648 4201 2651
rect 4862 2648 4865 2658
rect 4882 2648 4889 2651
rect 5174 2648 5182 2651
rect 142 2641 145 2648
rect 4862 2642 4866 2644
rect 134 2638 145 2641
rect 1514 2638 1517 2642
rect 1610 2638 1613 2642
rect 1982 2638 1990 2641
rect 3638 2638 3646 2641
rect 4338 2638 4345 2641
rect 4572 2638 4574 2642
rect 4684 2638 4686 2642
rect 5070 2638 5094 2641
rect 5162 2638 5163 2642
rect 1302 2628 1305 2638
rect 5070 2628 5073 2638
rect 5133 2628 5134 2632
rect 3066 2618 3070 2622
rect 4762 2618 4764 2622
rect 4813 2618 4814 2622
rect 5285 2618 5286 2622
rect 344 2603 346 2607
rect 350 2603 353 2607
rect 357 2603 360 2607
rect 1368 2603 1370 2607
rect 1374 2603 1377 2607
rect 1381 2603 1384 2607
rect 2392 2603 2394 2607
rect 2398 2603 2401 2607
rect 2405 2603 2408 2607
rect 3416 2603 3418 2607
rect 3422 2603 3425 2607
rect 3429 2603 3432 2607
rect 4440 2603 4442 2607
rect 4446 2603 4449 2607
rect 4453 2603 4456 2607
rect 92 2588 94 2592
rect 346 2588 350 2592
rect 450 2588 451 2592
rect 578 2588 579 2592
rect 693 2588 694 2592
rect 717 2588 718 2592
rect 850 2588 851 2592
rect 893 2588 894 2592
rect 1334 2588 1342 2591
rect 1354 2588 1361 2591
rect 1706 2588 1707 2592
rect 3053 2588 3054 2592
rect 4266 2588 4268 2592
rect 4332 2588 4334 2592
rect 3982 2572 3985 2581
rect 4478 2572 4481 2581
rect 2614 2568 2622 2571
rect 3122 2568 3129 2571
rect 4171 2568 4174 2572
rect 4382 2568 4393 2571
rect 4498 2568 4505 2571
rect 5140 2568 5142 2572
rect 742 2561 745 2568
rect 4390 2562 4393 2568
rect 742 2558 753 2561
rect 866 2558 881 2561
rect 2390 2558 2406 2561
rect 3074 2558 3081 2561
rect 3374 2558 3385 2561
rect 3394 2558 3398 2562
rect 3934 2558 3977 2561
rect 4486 2558 4505 2561
rect 4578 2558 4582 2562
rect 4854 2558 4865 2561
rect 4862 2552 4865 2558
rect 22 2548 38 2551
rect 154 2548 161 2551
rect 170 2548 185 2551
rect 230 2548 262 2551
rect 366 2548 390 2551
rect 646 2548 657 2551
rect 694 2548 702 2551
rect 706 2548 713 2551
rect 898 2548 932 2551
rect 942 2548 977 2551
rect 46 2538 62 2541
rect 110 2538 118 2541
rect 258 2538 265 2541
rect 366 2538 369 2548
rect 654 2542 657 2548
rect 974 2542 977 2548
rect 1598 2548 1614 2551
rect 2170 2548 2177 2551
rect 2562 2548 2577 2551
rect 2846 2548 2854 2551
rect 3054 2548 3062 2551
rect 3102 2548 3110 2551
rect 3398 2548 3441 2551
rect 3766 2548 3774 2551
rect 3846 2548 3865 2551
rect 3870 2548 3894 2551
rect 4238 2548 4249 2551
rect 4550 2548 4558 2551
rect 4586 2548 4609 2551
rect 4974 2548 5001 2551
rect 5222 2548 5257 2551
rect 4246 2542 4249 2548
rect 702 2538 710 2541
rect 786 2538 793 2541
rect 1838 2538 1866 2541
rect 2046 2538 2058 2541
rect 2382 2538 2398 2541
rect 3438 2538 3473 2541
rect 4058 2538 4073 2541
rect 4294 2538 4302 2541
rect 4354 2538 4361 2541
rect 4398 2538 4406 2541
rect 4594 2538 4601 2541
rect 4622 2538 4625 2548
rect 4738 2538 4745 2541
rect 4790 2538 4793 2548
rect 4886 2541 4889 2548
rect 4878 2538 4889 2541
rect 5014 2538 5017 2548
rect 5254 2542 5257 2548
rect 5270 2538 5281 2541
rect 274 2528 289 2531
rect 610 2528 625 2531
rect 958 2528 966 2531
rect 1030 2528 1041 2531
rect 2814 2528 2825 2531
rect 3358 2531 3362 2533
rect 3358 2528 3369 2531
rect 3946 2528 3961 2531
rect 4358 2528 4361 2538
rect 5270 2532 5273 2538
rect 1156 2518 1158 2522
rect 3934 2518 3950 2521
rect 4014 2518 4022 2521
rect 4772 2518 4774 2522
rect 4869 2518 4870 2522
rect 4978 2518 4979 2522
rect 5042 2518 5044 2522
rect 5218 2518 5220 2522
rect 856 2503 858 2507
rect 862 2503 865 2507
rect 869 2503 872 2507
rect 1872 2503 1874 2507
rect 1878 2503 1881 2507
rect 1885 2503 1888 2507
rect 2904 2503 2906 2507
rect 2910 2503 2913 2507
rect 2917 2503 2920 2507
rect 3928 2503 3930 2507
rect 3934 2503 3937 2507
rect 3941 2503 3944 2507
rect 4952 2503 4954 2507
rect 4958 2503 4961 2507
rect 4965 2503 4968 2507
rect 146 2488 148 2492
rect 458 2488 460 2492
rect 604 2488 606 2492
rect 650 2488 652 2492
rect 690 2488 692 2492
rect 794 2488 801 2491
rect 858 2488 859 2492
rect 1558 2488 1566 2491
rect 2870 2488 2886 2491
rect 4085 2488 4086 2492
rect 4882 2488 4883 2492
rect 102 2478 113 2481
rect 186 2478 201 2481
rect 2510 2478 2521 2481
rect 3822 2478 3830 2482
rect 3934 2478 3942 2481
rect 4482 2478 4489 2482
rect 70 2471 74 2472
rect 78 2471 81 2478
rect 70 2468 81 2471
rect 110 2472 113 2478
rect 2518 2472 2521 2478
rect 222 2468 233 2471
rect 246 2468 260 2471
rect 298 2468 313 2471
rect 398 2468 409 2471
rect 222 2462 225 2468
rect 246 2462 249 2468
rect 370 2458 385 2461
rect 438 2461 441 2471
rect 678 2462 681 2471
rect 830 2468 849 2471
rect 1114 2468 1121 2471
rect 1158 2468 1174 2471
rect 1190 2468 1201 2471
rect 1238 2468 1246 2471
rect 1262 2468 1289 2471
rect 1326 2468 1334 2471
rect 1342 2468 1358 2471
rect 1438 2468 1446 2471
rect 430 2458 441 2461
rect 530 2458 553 2461
rect 866 2458 897 2461
rect 930 2458 945 2461
rect 1086 2458 1126 2461
rect 1218 2458 1225 2461
rect 1322 2458 1337 2461
rect 1582 2461 1585 2471
rect 1942 2468 1953 2471
rect 2162 2468 2170 2471
rect 2266 2468 2273 2471
rect 1574 2458 1585 2461
rect 2534 2461 2537 2471
rect 2646 2468 2658 2471
rect 3022 2468 3025 2478
rect 3822 2472 3825 2478
rect 4486 2472 4489 2478
rect 3646 2468 3681 2471
rect 3786 2468 3793 2471
rect 3838 2468 3852 2471
rect 3938 2468 3969 2471
rect 4402 2468 4409 2471
rect 4414 2468 4430 2471
rect 4610 2468 4617 2471
rect 4622 2468 4630 2471
rect 4846 2468 4857 2471
rect 4862 2468 4870 2471
rect 1574 2456 1578 2458
rect 246 2448 257 2451
rect 862 2448 886 2451
rect 906 2448 913 2451
rect 1198 2448 1209 2451
rect 1206 2442 1209 2448
rect 262 2438 289 2441
rect 1298 2438 1306 2441
rect 2518 2441 2521 2461
rect 2526 2458 2537 2461
rect 3338 2458 3345 2461
rect 3534 2461 3537 2468
rect 3534 2458 3545 2461
rect 3646 2458 3654 2461
rect 3774 2458 3798 2461
rect 3806 2458 3825 2461
rect 4242 2458 4249 2461
rect 4502 2458 4513 2461
rect 4594 2458 4601 2461
rect 4654 2458 4670 2461
rect 4686 2458 4705 2461
rect 4710 2458 4729 2461
rect 4766 2461 4769 2468
rect 4766 2458 4777 2461
rect 4826 2458 4833 2461
rect 5026 2458 5033 2461
rect 5150 2458 5158 2461
rect 2526 2456 2530 2458
rect 3310 2452 3313 2458
rect 3358 2456 3362 2458
rect 3305 2448 3313 2452
rect 3718 2451 3721 2458
rect 3710 2448 3721 2451
rect 3822 2448 3825 2458
rect 4118 2452 4121 2458
rect 4510 2452 4513 2458
rect 4118 2448 4127 2452
rect 4446 2448 4454 2451
rect 4814 2448 4825 2451
rect 2518 2438 2526 2441
rect 2578 2438 2581 2442
rect 3878 2441 3881 2448
rect 3854 2438 3881 2441
rect 4006 2441 4009 2448
rect 3890 2438 3897 2441
rect 4006 2438 4017 2441
rect 4205 2438 4206 2442
rect 4518 2438 4526 2441
rect 4902 2438 4910 2441
rect 354 2418 361 2421
rect 386 2418 387 2422
rect 1130 2418 1131 2422
rect 3621 2418 3622 2422
rect 4173 2418 4174 2422
rect 4573 2418 4574 2422
rect 5205 2418 5206 2422
rect 344 2403 346 2407
rect 350 2403 353 2407
rect 357 2403 360 2407
rect 1368 2403 1370 2407
rect 1374 2403 1377 2407
rect 1381 2403 1384 2407
rect 2392 2403 2394 2407
rect 2398 2403 2401 2407
rect 2405 2403 2408 2407
rect 3416 2403 3418 2407
rect 3422 2403 3425 2407
rect 3429 2403 3432 2407
rect 4440 2403 4442 2407
rect 4446 2403 4449 2407
rect 4453 2403 4456 2407
rect 85 2388 86 2392
rect 274 2388 275 2392
rect 554 2388 556 2392
rect 842 2388 849 2391
rect 1556 2388 1558 2392
rect 1612 2388 1614 2392
rect 2164 2388 2166 2392
rect 3452 2388 3454 2392
rect 5181 2388 5182 2392
rect 5213 2378 5214 2382
rect 6 2368 17 2371
rect 418 2368 425 2371
rect 594 2368 601 2371
rect 634 2368 662 2371
rect 1022 2368 1030 2371
rect 1802 2368 1809 2371
rect 1970 2368 1977 2371
rect 2010 2368 2025 2371
rect 2862 2368 2889 2371
rect 2894 2368 2902 2371
rect 3250 2368 3266 2371
rect 3990 2368 3998 2371
rect 4243 2368 4246 2372
rect 4942 2368 4950 2371
rect 14 2362 17 2368
rect 46 2358 54 2361
rect 118 2361 121 2368
rect 2886 2362 2890 2364
rect 62 2358 73 2361
rect 118 2358 137 2361
rect 202 2358 209 2361
rect 238 2358 249 2361
rect 406 2358 425 2361
rect 710 2358 721 2361
rect 822 2358 830 2361
rect 990 2358 998 2361
rect 1130 2358 1137 2361
rect 1166 2358 1177 2361
rect 1668 2358 1670 2362
rect 2966 2361 2969 2368
rect 2958 2358 2969 2361
rect 3274 2358 3278 2362
rect 3330 2358 3334 2362
rect 3350 2358 3358 2361
rect 3522 2358 3529 2361
rect 230 2348 238 2351
rect 518 2351 521 2358
rect 614 2351 617 2358
rect 518 2348 529 2351
rect 606 2348 617 2351
rect 814 2348 822 2351
rect 942 2348 950 2351
rect 1062 2351 1065 2358
rect 1034 2348 1041 2351
rect 1046 2348 1065 2351
rect 1170 2348 1177 2351
rect 1894 2348 1902 2351
rect 1910 2348 1918 2351
rect 142 2338 150 2341
rect 342 2338 358 2341
rect 454 2338 465 2341
rect 885 2338 886 2342
rect 1066 2338 1073 2341
rect 1134 2338 1145 2341
rect 1518 2338 1529 2341
rect 1890 2338 1897 2341
rect 2030 2341 2033 2348
rect 2306 2348 2313 2351
rect 2942 2342 2945 2351
rect 3006 2348 3030 2351
rect 3058 2348 3081 2351
rect 3166 2348 3174 2351
rect 3626 2348 3657 2351
rect 3670 2348 3689 2351
rect 3734 2351 3737 2361
rect 3938 2358 3953 2361
rect 4274 2358 4281 2361
rect 4398 2358 4409 2361
rect 4774 2358 4801 2361
rect 5014 2361 5017 2368
rect 5014 2358 5025 2361
rect 5142 2358 5169 2361
rect 3718 2348 3737 2351
rect 3802 2348 3809 2351
rect 3826 2348 3833 2351
rect 4078 2351 4081 2358
rect 4398 2352 4401 2358
rect 4078 2348 4089 2351
rect 4330 2348 4361 2351
rect 4594 2348 4625 2351
rect 4854 2348 4865 2351
rect 4914 2348 4921 2351
rect 2030 2338 2042 2341
rect 2482 2338 2497 2341
rect 3018 2338 3025 2341
rect 3170 2338 3177 2341
rect 142 2328 145 2338
rect 350 2328 374 2331
rect 1030 2328 1038 2331
rect 1182 2328 1185 2338
rect 1518 2332 1521 2338
rect 2830 2328 2841 2331
rect 2942 2328 2950 2331
rect 3054 2331 3057 2338
rect 3046 2328 3057 2331
rect 3174 2328 3177 2338
rect 3510 2338 3521 2341
rect 3670 2338 3673 2348
rect 3686 2338 3705 2341
rect 3786 2338 3793 2341
rect 3798 2338 3801 2348
rect 3846 2338 3865 2341
rect 3902 2338 3910 2341
rect 3926 2338 3942 2341
rect 4358 2338 4361 2348
rect 4430 2338 4446 2341
rect 4450 2338 4457 2341
rect 4646 2338 4654 2341
rect 4702 2338 4724 2341
rect 4798 2338 4801 2348
rect 4854 2338 4857 2348
rect 4886 2338 4894 2341
rect 4902 2338 4910 2341
rect 4922 2338 4929 2341
rect 4990 2338 4998 2341
rect 5074 2338 5076 2342
rect 5094 2338 5106 2341
rect 5302 2338 5310 2341
rect 3182 2328 3190 2331
rect 3246 2331 3249 2338
rect 3518 2332 3521 2338
rect 3238 2328 3249 2331
rect 3822 2328 3830 2331
rect 4262 2331 4266 2333
rect 4270 2331 4273 2338
rect 5094 2332 5097 2338
rect 4262 2328 4273 2331
rect 4294 2328 4302 2331
rect 402 2318 403 2322
rect 2882 2318 2889 2321
rect 3089 2318 3102 2321
rect 3206 2321 3209 2328
rect 3206 2318 3217 2321
rect 3306 2318 3307 2322
rect 3554 2318 3556 2322
rect 3610 2318 3612 2322
rect 4377 2318 4398 2321
rect 4450 2318 4457 2321
rect 4532 2318 4534 2322
rect 4954 2318 4969 2321
rect 5005 2318 5006 2322
rect 856 2303 858 2307
rect 862 2303 865 2307
rect 869 2303 872 2307
rect 1872 2303 1874 2307
rect 1878 2303 1881 2307
rect 1885 2303 1888 2307
rect 2904 2303 2906 2307
rect 2910 2303 2913 2307
rect 2917 2303 2920 2307
rect 3928 2303 3930 2307
rect 3934 2303 3937 2307
rect 3941 2303 3944 2307
rect 4952 2303 4954 2307
rect 4958 2303 4961 2307
rect 4965 2303 4968 2307
rect 26 2288 28 2292
rect 140 2288 142 2292
rect 268 2288 270 2292
rect 394 2288 395 2292
rect 506 2288 508 2292
rect 628 2288 630 2292
rect 898 2288 905 2291
rect 1316 2288 1318 2292
rect 1394 2288 1401 2291
rect 1477 2288 1478 2292
rect 1522 2288 1523 2292
rect 1621 2288 1622 2292
rect 1970 2288 1971 2292
rect 2149 2288 2150 2292
rect 2174 2288 2182 2291
rect 2620 2288 2622 2292
rect 3554 2288 3556 2292
rect 4186 2288 4188 2292
rect 4818 2288 4820 2292
rect 1166 2272 1169 2278
rect 326 2268 334 2271
rect 478 2262 481 2271
rect 590 2268 601 2271
rect 694 2268 705 2271
rect 878 2268 886 2271
rect 1166 2268 1170 2272
rect 1350 2268 1358 2271
rect 1502 2271 1505 2281
rect 3990 2278 3998 2282
rect 4342 2278 4353 2281
rect 4630 2278 4638 2281
rect 4754 2278 4761 2282
rect 1486 2268 1497 2271
rect 1502 2268 1510 2271
rect 1594 2268 1601 2271
rect 1890 2268 1913 2271
rect 1946 2268 1961 2271
rect 2270 2268 2281 2271
rect 2374 2268 2385 2271
rect 2734 2271 2738 2274
rect 3990 2272 3993 2278
rect 4342 2272 4345 2278
rect 4758 2272 4761 2278
rect 2734 2268 2745 2271
rect 2942 2268 2961 2271
rect 2998 2268 3014 2271
rect 3062 2268 3073 2271
rect 3334 2268 3345 2271
rect 3386 2268 3398 2271
rect 3802 2268 3809 2271
rect 598 2262 601 2268
rect 174 2258 193 2261
rect 450 2258 457 2261
rect 562 2258 577 2261
rect 670 2258 689 2261
rect 950 2258 990 2261
rect 1262 2258 1278 2261
rect 1562 2258 1569 2261
rect 1838 2258 1857 2261
rect 2966 2261 2969 2268
rect 3334 2262 3337 2268
rect 2966 2258 2977 2261
rect 3098 2258 3105 2261
rect 3654 2258 3678 2261
rect 3766 2258 3769 2268
rect 3822 2261 3825 2271
rect 4070 2268 4078 2271
rect 4442 2268 4449 2271
rect 4474 2268 4481 2271
rect 4502 2268 4510 2271
rect 4670 2268 4678 2271
rect 5058 2268 5073 2271
rect 5134 2268 5142 2271
rect 5166 2268 5185 2271
rect 5234 2268 5241 2271
rect 3806 2258 3825 2261
rect 3854 2261 3857 2268
rect 3854 2258 3865 2261
rect 4050 2258 4057 2261
rect 4062 2258 4086 2261
rect 4114 2258 4121 2261
rect 4310 2261 4313 2268
rect 4310 2258 4321 2261
rect 4402 2258 4409 2261
rect 4462 2258 4486 2261
rect 4514 2258 4521 2261
rect 4578 2258 4585 2261
rect 4638 2261 4641 2268
rect 4662 2261 4665 2268
rect 4638 2258 4649 2261
rect 4654 2258 4665 2261
rect 4670 2258 4681 2261
rect 4702 2258 4713 2261
rect 4938 2258 4953 2261
rect 5046 2261 5049 2268
rect 5038 2258 5049 2261
rect 5110 2258 5134 2261
rect 5226 2258 5233 2261
rect 190 2252 193 2258
rect 670 2248 673 2258
rect 890 2248 905 2251
rect 1358 2248 1369 2251
rect 2118 2248 2129 2251
rect 3302 2248 3313 2251
rect 3954 2248 3961 2251
rect 4390 2248 4401 2251
rect 5230 2248 5233 2258
rect 5270 2251 5273 2271
rect 5270 2248 5278 2251
rect 1366 2241 1369 2248
rect 1366 2238 1398 2241
rect 1434 2238 1436 2242
rect 2026 2238 2028 2242
rect 3990 2241 3994 2244
rect 3978 2238 3994 2241
rect 4758 2241 4762 2244
rect 4758 2238 4785 2241
rect 4022 2228 4025 2238
rect 1546 2218 1547 2222
rect 1878 2218 1886 2221
rect 3044 2218 3046 2222
rect 3146 2218 3147 2222
rect 3186 2218 3188 2222
rect 3252 2218 3254 2222
rect 3682 2218 3683 2222
rect 4186 2218 4188 2222
rect 4252 2218 4254 2222
rect 4922 2218 4923 2222
rect 4994 2218 4995 2222
rect 344 2203 346 2207
rect 350 2203 353 2207
rect 357 2203 360 2207
rect 1368 2203 1370 2207
rect 1374 2203 1377 2207
rect 1381 2203 1384 2207
rect 2392 2203 2394 2207
rect 2398 2203 2401 2207
rect 2405 2203 2408 2207
rect 3416 2203 3418 2207
rect 3422 2203 3425 2207
rect 3429 2203 3432 2207
rect 4440 2203 4442 2207
rect 4446 2203 4449 2207
rect 4453 2203 4456 2207
rect 324 2188 326 2192
rect 570 2188 571 2192
rect 1717 2188 1718 2192
rect 2173 2188 2174 2192
rect 2394 2188 2409 2191
rect 2506 2188 2508 2192
rect 2946 2188 2948 2192
rect 3002 2188 3004 2192
rect 3652 2188 3654 2192
rect 3698 2188 3700 2192
rect 4370 2188 4372 2192
rect 5301 2188 5302 2192
rect 46 2168 54 2171
rect 166 2168 174 2171
rect 686 2168 697 2171
rect 1546 2168 1547 2172
rect 1638 2168 1646 2171
rect 3572 2168 3574 2172
rect 4310 2168 4321 2171
rect 4614 2171 4617 2181
rect 4594 2168 4617 2171
rect 4949 2168 4950 2172
rect 686 2162 689 2168
rect 74 2158 81 2161
rect 442 2158 449 2161
rect 410 2148 433 2151
rect 538 2148 569 2151
rect 618 2148 625 2151
rect 702 2151 705 2161
rect 746 2158 750 2162
rect 1286 2158 1294 2161
rect 2102 2158 2113 2161
rect 2434 2158 2438 2162
rect 2614 2158 2623 2162
rect 2764 2158 2766 2162
rect 4022 2158 4030 2161
rect 4214 2161 4217 2168
rect 4310 2162 4313 2168
rect 4206 2158 4217 2161
rect 4598 2158 4601 2168
rect 4702 2158 4713 2161
rect 4898 2158 4905 2161
rect 5006 2158 5014 2161
rect 5030 2161 5033 2168
rect 5030 2158 5041 2161
rect 5106 2158 5110 2162
rect 2614 2152 2617 2158
rect 4206 2156 4210 2158
rect 702 2148 721 2151
rect 730 2148 745 2151
rect 934 2148 942 2151
rect 62 2138 70 2141
rect 382 2141 385 2148
rect 702 2142 705 2148
rect 1686 2148 1702 2151
rect 1806 2148 1814 2151
rect 1902 2148 1921 2151
rect 2146 2148 2153 2151
rect 2186 2148 2193 2151
rect 2418 2148 2433 2151
rect 2450 2148 2457 2151
rect 3042 2148 3049 2151
rect 3210 2148 3217 2151
rect 3254 2148 3262 2151
rect 3290 2148 3297 2151
rect 3382 2151 3386 2154
rect 4606 2152 4610 2154
rect 3382 2148 3393 2151
rect 3510 2148 3545 2151
rect 3814 2148 3833 2151
rect 3926 2148 3969 2151
rect 4054 2148 4073 2151
rect 4294 2148 4305 2151
rect 4450 2148 4457 2151
rect 4518 2148 4553 2151
rect 4714 2148 4721 2151
rect 4726 2148 4758 2151
rect 4802 2148 4817 2151
rect 4950 2148 4958 2151
rect 5090 2148 5102 2151
rect 5134 2148 5145 2151
rect 2566 2146 2570 2148
rect 382 2138 393 2141
rect 730 2138 737 2141
rect 830 2138 878 2141
rect 1606 2138 1625 2141
rect 1654 2138 1666 2141
rect 1726 2138 1745 2141
rect 1862 2138 1878 2141
rect 2182 2138 2201 2141
rect 2230 2138 2241 2141
rect 2274 2138 2281 2141
rect 2382 2138 2398 2141
rect 2414 2138 2422 2141
rect 2698 2138 2705 2141
rect 3318 2138 3326 2141
rect 3390 2138 3393 2148
rect 3410 2138 3433 2141
rect 3542 2138 3545 2148
rect 3906 2138 3913 2141
rect 4054 2138 4057 2148
rect 4294 2142 4297 2148
rect 4406 2141 4409 2148
rect 4398 2138 4409 2141
rect 4518 2138 4521 2148
rect 4550 2142 4553 2148
rect 4646 2138 4654 2141
rect 4854 2138 4862 2141
rect 4878 2138 4886 2141
rect 4914 2138 4921 2141
rect 5158 2138 5177 2141
rect 5246 2138 5249 2148
rect 5258 2138 5265 2141
rect 1654 2132 1657 2138
rect 382 2128 393 2131
rect 786 2128 793 2131
rect 866 2128 886 2131
rect 2414 2128 2417 2138
rect 3182 2128 3190 2131
rect 4030 2131 4033 2138
rect 4030 2128 4046 2131
rect 4206 2131 4210 2133
rect 5014 2132 5017 2138
rect 4206 2128 4217 2131
rect 4554 2128 4558 2132
rect 4886 2128 4894 2131
rect 4902 2128 4913 2131
rect 5014 2128 5022 2132
rect 5158 2128 5161 2138
rect 85 2118 86 2122
rect 222 2118 230 2121
rect 250 2118 255 2122
rect 498 2118 519 2121
rect 2690 2118 2691 2122
rect 2902 2118 2918 2121
rect 3366 2118 3374 2121
rect 3406 2118 3422 2121
rect 3450 2118 3452 2122
rect 3874 2118 3876 2122
rect 4490 2118 4492 2122
rect 856 2103 858 2107
rect 862 2103 865 2107
rect 869 2103 872 2107
rect 1872 2103 1874 2107
rect 1878 2103 1881 2107
rect 1885 2103 1888 2107
rect 2904 2103 2906 2107
rect 2910 2103 2913 2107
rect 2917 2103 2920 2107
rect 3928 2103 3930 2107
rect 3934 2103 3937 2107
rect 3941 2103 3944 2107
rect 4952 2103 4954 2107
rect 4958 2103 4961 2107
rect 4965 2103 4968 2107
rect 237 2088 238 2092
rect 405 2088 406 2092
rect 429 2088 430 2092
rect 620 2088 622 2092
rect 770 2088 772 2092
rect 1420 2088 1422 2092
rect 2109 2088 2110 2092
rect 2189 2088 2190 2092
rect 2662 2088 2670 2091
rect 2842 2088 2843 2092
rect 2898 2088 2900 2092
rect 3650 2088 3652 2092
rect 3716 2088 3718 2092
rect 3902 2088 3910 2091
rect 4018 2088 4020 2092
rect 4524 2088 4526 2092
rect 4626 2088 4628 2092
rect 4682 2088 4684 2092
rect 4748 2088 4750 2092
rect 4794 2088 4796 2092
rect 4850 2088 4852 2092
rect 4930 2088 4932 2092
rect 5090 2088 5091 2092
rect 1018 2078 1022 2082
rect 1570 2078 1577 2081
rect 1710 2078 1721 2081
rect 62 2062 65 2071
rect 190 2071 193 2078
rect 1310 2072 1313 2078
rect 2318 2072 2321 2081
rect 2534 2078 2545 2081
rect 2590 2078 2601 2081
rect 3204 2078 3206 2082
rect 3354 2078 3361 2082
rect 3358 2072 3361 2078
rect 3750 2076 3754 2078
rect 190 2068 201 2071
rect 534 2068 542 2071
rect 958 2068 977 2071
rect 1310 2068 1314 2072
rect 34 2058 49 2061
rect 326 2058 337 2061
rect 390 2058 398 2061
rect 514 2058 521 2061
rect 530 2058 553 2061
rect 686 2058 694 2061
rect 898 2058 905 2061
rect 974 2058 993 2061
rect 1034 2058 1049 2061
rect 1526 2061 1529 2071
rect 1858 2068 1865 2071
rect 1870 2068 1886 2071
rect 1526 2058 1537 2061
rect 1786 2058 1794 2061
rect 2046 2061 2049 2071
rect 2358 2068 2366 2071
rect 2542 2068 2553 2071
rect 1862 2058 1897 2061
rect 2014 2058 2049 2061
rect 2542 2062 2545 2068
rect 2742 2062 2745 2071
rect 3158 2062 3161 2071
rect 3236 2068 3238 2072
rect 3442 2068 3457 2071
rect 3522 2068 3529 2071
rect 4046 2068 4054 2071
rect 4198 2068 4206 2071
rect 4250 2068 4265 2071
rect 4270 2068 4278 2071
rect 4374 2068 4386 2071
rect 4878 2068 4897 2071
rect 4906 2068 4913 2071
rect 2350 2058 2374 2061
rect 2794 2058 2817 2061
rect 3086 2058 3110 2061
rect 3494 2058 3502 2061
rect 3594 2058 3596 2062
rect 4062 2058 4081 2061
rect 4902 2058 4910 2061
rect 5038 2058 5057 2061
rect 5078 2061 5081 2071
rect 5074 2058 5081 2061
rect 5094 2068 5105 2071
rect 5094 2062 5097 2068
rect 5114 2058 5140 2061
rect 62 2048 73 2051
rect 318 2051 321 2058
rect 318 2048 329 2051
rect 574 2048 582 2051
rect 990 2048 993 2058
rect 1790 2056 1794 2058
rect 998 2048 1017 2051
rect 1770 2048 1777 2051
rect 2062 2048 2073 2051
rect 2394 2048 2417 2051
rect 2718 2048 2745 2051
rect 3158 2048 3185 2051
rect 3342 2051 3345 2058
rect 3306 2048 3313 2051
rect 3334 2048 3345 2051
rect 3494 2048 3505 2051
rect 4134 2048 4142 2051
rect 4222 2051 4225 2058
rect 4222 2048 4233 2051
rect 5070 2048 5078 2051
rect 398 2042 402 2044
rect 170 2038 177 2041
rect 390 2038 398 2041
rect 998 2038 1006 2041
rect 1746 2038 1753 2041
rect 3114 2038 3115 2042
rect 3178 2038 3198 2041
rect 3226 2038 3233 2041
rect 3557 2038 3558 2042
rect 4114 2038 4121 2041
rect 4170 2038 4172 2042
rect 4570 2038 4572 2042
rect 5194 2038 5196 2042
rect 2146 2028 2150 2032
rect 2670 2028 2673 2038
rect 3413 2028 3414 2032
rect 5058 2028 5059 2032
rect 18 2018 19 2022
rect 210 2018 211 2022
rect 2349 2018 2350 2022
rect 2378 2018 2379 2022
rect 344 2003 346 2007
rect 350 2003 353 2007
rect 357 2003 360 2007
rect 1368 2003 1370 2007
rect 1374 2003 1377 2007
rect 1381 2003 1384 2007
rect 2392 2003 2394 2007
rect 2398 2003 2401 2007
rect 2405 2003 2408 2007
rect 3416 2003 3418 2007
rect 3422 2003 3425 2007
rect 3429 2003 3432 2007
rect 4440 2003 4442 2007
rect 4446 2003 4449 2007
rect 4453 2003 4456 2007
rect 170 1988 174 1992
rect 402 1988 403 1992
rect 1282 1988 1283 1992
rect 1357 1988 1358 1992
rect 1476 1988 1478 1992
rect 2797 1988 2798 1992
rect 4164 1988 4166 1992
rect 4210 1988 4212 1992
rect 5004 1988 5006 1992
rect 1420 1978 1422 1982
rect 1838 1972 1841 1981
rect 2610 1978 2614 1982
rect 226 1968 233 1971
rect 266 1968 273 1971
rect 1054 1968 1062 1971
rect 4004 1968 4006 1972
rect 4315 1968 4318 1972
rect 414 1958 425 1961
rect 534 1961 537 1968
rect 534 1958 561 1961
rect 858 1958 870 1961
rect 90 1948 97 1951
rect 106 1948 121 1951
rect 334 1948 342 1951
rect 394 1948 401 1951
rect 478 1951 482 1954
rect 478 1948 489 1951
rect 510 1948 518 1951
rect 590 1948 598 1951
rect 134 1938 145 1941
rect 194 1938 201 1941
rect 330 1938 361 1941
rect 638 1941 641 1948
rect 842 1948 881 1951
rect 894 1948 910 1951
rect 930 1948 937 1951
rect 1062 1951 1065 1958
rect 1674 1957 1676 1961
rect 3290 1958 3297 1961
rect 3406 1961 3409 1968
rect 3406 1958 3417 1961
rect 4350 1958 4361 1961
rect 1062 1948 1073 1951
rect 1114 1948 1121 1951
rect 602 1938 609 1941
rect 630 1938 641 1941
rect 894 1938 897 1948
rect 946 1938 953 1941
rect 1086 1941 1089 1948
rect 1526 1948 1537 1951
rect 1550 1948 1558 1951
rect 1602 1948 1620 1951
rect 1694 1948 1726 1951
rect 1754 1948 1761 1951
rect 1950 1948 1958 1951
rect 2342 1948 2350 1951
rect 2358 1948 2377 1951
rect 2558 1948 2569 1951
rect 2642 1948 2649 1951
rect 1534 1942 1537 1948
rect 1062 1938 1073 1941
rect 1086 1938 1097 1941
rect 1330 1938 1337 1941
rect 1646 1938 1654 1941
rect 1694 1938 1697 1948
rect 1742 1938 1750 1941
rect 2194 1938 2209 1941
rect 2358 1941 2361 1948
rect 2566 1942 2569 1948
rect 2830 1948 2841 1951
rect 2830 1942 2833 1948
rect 3270 1948 3281 1951
rect 2354 1938 2361 1941
rect 2466 1938 2473 1941
rect 2482 1938 2489 1941
rect 2654 1938 2666 1941
rect 2902 1938 2929 1941
rect 3174 1938 3198 1941
rect 3246 1938 3254 1941
rect 3358 1938 3361 1948
rect 3462 1941 3465 1951
rect 3470 1948 3502 1951
rect 3718 1948 3742 1951
rect 3794 1948 3809 1951
rect 3966 1948 3974 1951
rect 4102 1948 4110 1951
rect 3446 1938 3465 1941
rect 3838 1938 3850 1941
rect 4046 1941 4049 1948
rect 4038 1938 4049 1941
rect 4102 1938 4105 1948
rect 4374 1948 4409 1951
rect 4494 1951 4497 1961
rect 4490 1948 4497 1951
rect 4836 1958 4838 1962
rect 4510 1951 4513 1958
rect 4510 1948 4521 1951
rect 4406 1942 4409 1948
rect 4130 1938 4137 1941
rect 4450 1938 4481 1941
rect 4542 1938 4550 1941
rect 4746 1938 4753 1941
rect 5226 1938 5233 1941
rect 214 1932 217 1938
rect 210 1928 217 1932
rect 510 1931 513 1938
rect 510 1928 526 1931
rect 838 1928 854 1931
rect 950 1928 953 1938
rect 2062 1931 2065 1938
rect 2662 1936 2666 1938
rect 2054 1928 2065 1931
rect 2818 1928 2825 1931
rect 3246 1928 3249 1938
rect 3402 1928 3409 1931
rect 3414 1928 3441 1931
rect 3942 1928 3961 1931
rect 4334 1931 4338 1933
rect 4334 1928 4342 1931
rect 242 1918 244 1922
rect 810 1918 815 1922
rect 1866 1918 1867 1922
rect 1978 1918 1980 1922
rect 2090 1918 2091 1922
rect 2506 1918 2508 1922
rect 2578 1918 2579 1922
rect 2962 1918 2964 1922
rect 3516 1918 3518 1922
rect 3572 1918 3574 1922
rect 3942 1921 3945 1928
rect 3934 1918 3945 1921
rect 4570 1918 4572 1922
rect 4658 1918 4660 1922
rect 4714 1918 4716 1922
rect 4770 1918 4772 1922
rect 5266 1918 5268 1922
rect 856 1903 858 1907
rect 862 1903 865 1907
rect 869 1903 872 1907
rect 1872 1903 1874 1907
rect 1878 1903 1881 1907
rect 1885 1903 1888 1907
rect 2904 1903 2906 1907
rect 2910 1903 2913 1907
rect 2917 1903 2920 1907
rect 3928 1903 3930 1907
rect 3934 1903 3937 1907
rect 3941 1903 3944 1907
rect 4952 1903 4954 1907
rect 4958 1903 4961 1907
rect 4965 1903 4968 1907
rect 26 1888 28 1892
rect 194 1888 195 1892
rect 410 1888 412 1892
rect 458 1888 459 1892
rect 500 1888 502 1892
rect 538 1888 539 1892
rect 882 1888 889 1891
rect 1170 1888 1172 1892
rect 1556 1888 1558 1892
rect 1834 1888 1835 1892
rect 2237 1888 2238 1892
rect 2434 1888 2435 1892
rect 3484 1888 3486 1892
rect 4074 1888 4076 1892
rect 4140 1888 4142 1892
rect 4802 1888 4804 1892
rect 4858 1888 4860 1892
rect 4924 1888 4926 1892
rect 4996 1888 4998 1892
rect 5052 1888 5054 1892
rect 138 1878 153 1881
rect 270 1878 278 1882
rect 322 1878 329 1882
rect 554 1878 561 1881
rect 758 1878 769 1881
rect 862 1878 878 1881
rect 110 1871 113 1878
rect 270 1872 273 1878
rect 326 1872 329 1878
rect 100 1868 113 1871
rect 294 1868 313 1871
rect 718 1868 737 1871
rect 174 1858 182 1861
rect 286 1858 297 1861
rect 326 1858 345 1861
rect 902 1861 905 1871
rect 1086 1868 1094 1871
rect 1598 1871 1601 1878
rect 1590 1868 1601 1871
rect 1750 1868 1758 1871
rect 1814 1868 1822 1871
rect 1918 1871 1921 1881
rect 2914 1878 2926 1881
rect 3242 1878 3254 1881
rect 4178 1878 4185 1882
rect 3238 1874 3242 1878
rect 1830 1868 1849 1871
rect 1894 1868 1921 1871
rect 830 1858 849 1861
rect 902 1858 914 1861
rect 942 1861 945 1868
rect 942 1858 953 1861
rect 1006 1858 1014 1861
rect 1082 1858 1121 1861
rect 2062 1861 2065 1871
rect 2318 1868 2326 1871
rect 2418 1868 2425 1871
rect 2442 1868 2457 1871
rect 2602 1868 2609 1871
rect 2778 1868 2793 1871
rect 2822 1868 2838 1871
rect 2922 1868 2937 1871
rect 2062 1858 2094 1861
rect 2254 1861 2258 1864
rect 2990 1862 2993 1871
rect 3138 1868 3145 1871
rect 3150 1868 3161 1871
rect 3326 1871 3330 1872
rect 3334 1871 3337 1878
rect 4182 1872 4185 1878
rect 3326 1868 3337 1871
rect 3438 1868 3457 1871
rect 3158 1862 3161 1868
rect 4394 1868 4409 1871
rect 4438 1868 4462 1871
rect 4654 1868 4670 1871
rect 2250 1858 2258 1861
rect 2346 1858 2353 1861
rect 2634 1858 2649 1861
rect 2902 1858 2942 1861
rect 3050 1858 3057 1861
rect 3126 1858 3142 1861
rect 3354 1858 3361 1861
rect 3542 1858 3550 1861
rect 4302 1861 4305 1868
rect 4258 1858 4265 1861
rect 4294 1858 4305 1861
rect 4618 1858 4625 1861
rect 4830 1861 4833 1871
rect 4954 1868 4969 1871
rect 5182 1868 5201 1871
rect 4666 1858 4681 1861
rect 4830 1858 4838 1861
rect 286 1852 289 1858
rect 326 1852 329 1858
rect 910 1856 914 1858
rect 822 1848 833 1851
rect 1058 1848 1065 1851
rect 2398 1848 2422 1851
rect 3198 1851 3201 1858
rect 4190 1856 4194 1858
rect 5278 1856 5282 1858
rect 3190 1848 3201 1851
rect 3374 1848 3385 1851
rect 3394 1848 3398 1852
rect 4542 1848 4553 1851
rect 5278 1848 5289 1851
rect 2486 1838 2513 1841
rect 2554 1838 2577 1841
rect 3718 1841 3721 1848
rect 3710 1838 3721 1841
rect 4466 1838 4486 1841
rect 214 1828 217 1838
rect 690 1818 692 1822
rect 1077 1818 1078 1822
rect 1866 1818 1868 1822
rect 1970 1818 1972 1822
rect 2053 1818 2054 1822
rect 2122 1818 2123 1822
rect 2741 1818 2742 1822
rect 4084 1818 4086 1822
rect 4314 1818 4315 1822
rect 4746 1818 4748 1822
rect 5098 1818 5100 1822
rect 344 1803 346 1807
rect 350 1803 353 1807
rect 357 1803 360 1807
rect 1368 1803 1370 1807
rect 1374 1803 1377 1807
rect 1381 1803 1384 1807
rect 2392 1803 2394 1807
rect 2398 1803 2401 1807
rect 2405 1803 2408 1807
rect 3416 1803 3418 1807
rect 3422 1803 3425 1807
rect 3429 1803 3432 1807
rect 4440 1803 4442 1807
rect 4446 1803 4449 1807
rect 4453 1803 4456 1807
rect 117 1788 118 1792
rect 162 1788 163 1792
rect 202 1788 204 1792
rect 522 1788 524 1792
rect 1580 1788 1582 1792
rect 1810 1788 1812 1792
rect 1898 1788 1900 1792
rect 2618 1788 2619 1792
rect 3554 1788 3555 1792
rect 894 1772 897 1781
rect 4742 1772 4745 1781
rect 4878 1772 4881 1781
rect 54 1768 78 1771
rect 134 1768 142 1771
rect 390 1768 398 1771
rect 2322 1768 2323 1772
rect 4326 1768 4350 1771
rect 4858 1768 4865 1771
rect 46 1758 57 1761
rect 286 1761 289 1768
rect 270 1758 289 1761
rect 146 1748 161 1751
rect 422 1748 438 1751
rect 774 1751 777 1761
rect 978 1758 982 1762
rect 1042 1758 1046 1762
rect 1054 1758 1065 1761
rect 762 1748 777 1751
rect 790 1748 822 1751
rect 958 1748 966 1751
rect 1034 1748 1041 1751
rect 1062 1748 1081 1751
rect 1126 1751 1129 1761
rect 1774 1758 1782 1761
rect 2126 1758 2137 1761
rect 1110 1748 1129 1751
rect 230 1738 238 1741
rect 246 1738 262 1741
rect 346 1738 361 1741
rect 478 1738 489 1741
rect 802 1738 817 1741
rect 938 1738 945 1741
rect 962 1738 969 1741
rect 1078 1738 1081 1748
rect 1678 1751 1681 1758
rect 1654 1748 1681 1751
rect 1854 1748 1870 1751
rect 2334 1751 2337 1761
rect 2366 1758 2374 1761
rect 2646 1761 2649 1768
rect 2646 1758 2657 1761
rect 4282 1758 4289 1761
rect 4426 1758 4430 1762
rect 4594 1758 4598 1762
rect 4626 1758 4630 1762
rect 4810 1758 4814 1762
rect 4862 1758 4873 1761
rect 5286 1758 5302 1761
rect 3190 1753 3194 1758
rect 2334 1748 2350 1751
rect 2382 1748 2409 1751
rect 2422 1748 2433 1751
rect 2734 1748 2750 1751
rect 2902 1748 2918 1751
rect 1098 1738 1113 1741
rect 1406 1738 1422 1741
rect 1678 1738 1681 1748
rect 2422 1742 2425 1748
rect 1750 1738 1761 1741
rect 2022 1738 2033 1741
rect 2582 1741 2585 1748
rect 2582 1738 2593 1741
rect 2670 1738 2689 1741
rect 2702 1738 2710 1741
rect 2850 1738 2862 1741
rect 2946 1738 2961 1741
rect 3358 1738 3370 1741
rect 3466 1738 3489 1741
rect 3518 1741 3521 1748
rect 3958 1751 3962 1753
rect 3822 1748 3849 1751
rect 3854 1748 3865 1751
rect 3862 1742 3865 1748
rect 3958 1748 3982 1751
rect 4174 1748 4193 1751
rect 4398 1748 4414 1751
rect 4574 1748 4593 1751
rect 4598 1748 4614 1751
rect 4618 1748 4625 1751
rect 4782 1748 4806 1751
rect 4834 1748 4841 1751
rect 4978 1748 4985 1751
rect 5158 1748 5188 1751
rect 5254 1748 5270 1751
rect 3510 1738 3521 1741
rect 3978 1738 3985 1741
rect 4174 1738 4177 1748
rect 4310 1738 4324 1741
rect 4478 1738 4505 1741
rect 4534 1738 4550 1741
rect 4610 1738 4617 1741
rect 4670 1738 4678 1741
rect 4766 1738 4769 1748
rect 4790 1738 4798 1741
rect 4998 1738 5006 1741
rect 5158 1738 5161 1748
rect 5214 1738 5225 1741
rect 5266 1738 5273 1741
rect 706 1728 713 1731
rect 814 1728 817 1738
rect 926 1728 937 1731
rect 1070 1728 1073 1738
rect 3734 1728 3745 1731
rect 4234 1728 4246 1731
rect 4514 1728 4521 1731
rect 334 1718 342 1721
rect 2076 1718 2078 1722
rect 2226 1718 2228 1722
rect 2270 1718 2278 1721
rect 2794 1718 2796 1722
rect 2922 1718 2929 1721
rect 3082 1718 3084 1722
rect 3138 1718 3140 1722
rect 3602 1718 3603 1722
rect 4090 1718 4092 1722
rect 4146 1718 4148 1722
rect 856 1703 858 1707
rect 862 1703 865 1707
rect 869 1703 872 1707
rect 1872 1703 1874 1707
rect 1878 1703 1881 1707
rect 1885 1703 1888 1707
rect 2904 1703 2906 1707
rect 2910 1703 2913 1707
rect 2917 1703 2920 1707
rect 3928 1703 3930 1707
rect 3934 1703 3937 1707
rect 3941 1703 3944 1707
rect 4952 1703 4954 1707
rect 4958 1703 4961 1707
rect 4965 1703 4968 1707
rect 84 1688 86 1692
rect 140 1688 142 1692
rect 196 1688 198 1692
rect 596 1688 598 1692
rect 1020 1688 1022 1692
rect 1618 1688 1620 1692
rect 1762 1688 1764 1692
rect 1842 1688 1844 1692
rect 2050 1688 2052 1692
rect 2106 1688 2108 1692
rect 2389 1688 2390 1692
rect 2698 1688 2705 1691
rect 2844 1688 2846 1692
rect 3693 1688 3694 1692
rect 4466 1688 4468 1692
rect 4882 1688 4883 1692
rect 4982 1688 4990 1691
rect 5042 1688 5044 1692
rect 5276 1688 5278 1692
rect 2298 1678 2310 1681
rect 2410 1678 2425 1681
rect 2542 1678 2550 1681
rect 3318 1678 3329 1681
rect 3318 1672 3321 1678
rect 354 1668 361 1671
rect 674 1668 689 1671
rect 706 1668 713 1671
rect 774 1668 782 1671
rect 906 1668 913 1671
rect 1142 1662 1145 1671
rect 1330 1668 1337 1671
rect 1382 1668 1398 1671
rect 1674 1668 1681 1671
rect 378 1658 385 1661
rect 418 1658 457 1661
rect 778 1658 785 1661
rect 1050 1658 1057 1661
rect 1170 1658 1177 1661
rect 1710 1661 1713 1671
rect 1870 1668 1894 1671
rect 1918 1668 1929 1671
rect 2218 1668 2225 1671
rect 2318 1668 2337 1671
rect 2410 1668 2433 1671
rect 2454 1668 2465 1671
rect 2494 1668 2510 1671
rect 2518 1668 2526 1671
rect 2862 1668 2878 1671
rect 3390 1668 3430 1671
rect 3454 1671 3457 1681
rect 3594 1678 3601 1681
rect 4374 1678 4382 1681
rect 3438 1668 3457 1671
rect 3550 1668 3558 1671
rect 1918 1662 1921 1668
rect 2454 1662 2457 1668
rect 1702 1658 1713 1661
rect 1726 1658 1734 1661
rect 2150 1658 2174 1661
rect 2182 1658 2201 1661
rect 2238 1658 2246 1661
rect 2566 1658 2585 1661
rect 2660 1658 2690 1661
rect 3014 1658 3022 1661
rect 3126 1658 3134 1661
rect 3398 1658 3422 1661
rect 3458 1658 3465 1661
rect 3574 1658 3582 1661
rect 3670 1658 3689 1661
rect 4278 1661 4281 1671
rect 4294 1668 4313 1671
rect 4346 1668 4353 1671
rect 4410 1668 4417 1671
rect 4594 1668 4601 1671
rect 4638 1668 4652 1671
rect 4702 1668 4710 1671
rect 4278 1658 4297 1661
rect 4326 1658 4342 1661
rect 4518 1661 4521 1668
rect 4406 1658 4417 1661
rect 4510 1658 4521 1661
rect 4638 1658 4649 1661
rect 4682 1658 4689 1661
rect 4694 1658 4718 1661
rect 4758 1661 4761 1668
rect 4994 1668 5009 1671
rect 5014 1668 5025 1671
rect 5202 1668 5214 1671
rect 5242 1668 5249 1671
rect 4758 1658 4769 1661
rect 5118 1658 5129 1661
rect 5238 1658 5246 1661
rect 634 1648 638 1652
rect 858 1648 873 1651
rect 958 1648 966 1651
rect 1126 1648 1145 1651
rect 1182 1648 1193 1651
rect 1318 1648 1326 1651
rect 1890 1648 1897 1651
rect 1950 1648 1961 1651
rect 2246 1648 2257 1651
rect 2342 1651 2345 1658
rect 2342 1648 2353 1651
rect 2470 1651 2473 1658
rect 2686 1656 2690 1658
rect 2470 1648 2481 1651
rect 3370 1648 3377 1651
rect 3622 1648 3630 1651
rect 3686 1648 3689 1658
rect 4638 1652 4641 1658
rect 4734 1648 4745 1651
rect 1182 1642 1185 1648
rect 294 1638 302 1641
rect 1670 1638 1678 1641
rect 2650 1638 2652 1642
rect 4502 1641 4505 1648
rect 4518 1641 4522 1644
rect 4502 1638 4513 1641
rect 4518 1638 4545 1641
rect 506 1628 508 1632
rect 1102 1628 1105 1638
rect 413 1618 414 1622
rect 1205 1618 1206 1622
rect 1722 1618 1723 1622
rect 2205 1618 2206 1622
rect 3154 1618 3156 1622
rect 3597 1618 3598 1622
rect 4130 1618 4132 1622
rect 4196 1618 4198 1622
rect 4573 1618 4574 1622
rect 4722 1618 4723 1622
rect 5093 1618 5094 1622
rect 344 1603 346 1607
rect 350 1603 353 1607
rect 357 1603 360 1607
rect 1368 1603 1370 1607
rect 1374 1603 1377 1607
rect 1381 1603 1384 1607
rect 2392 1603 2394 1607
rect 2398 1603 2401 1607
rect 2405 1603 2408 1607
rect 3416 1603 3418 1607
rect 3422 1603 3425 1607
rect 3429 1603 3432 1607
rect 4440 1603 4442 1607
rect 4446 1603 4449 1607
rect 4453 1603 4456 1607
rect 325 1588 326 1592
rect 450 1588 454 1592
rect 572 1588 574 1592
rect 1490 1588 1491 1592
rect 1701 1588 1702 1592
rect 1813 1588 1814 1592
rect 1877 1588 1878 1592
rect 2125 1588 2126 1592
rect 2794 1588 2796 1592
rect 4658 1588 4660 1592
rect 4934 1588 4942 1591
rect 130 1568 131 1572
rect 974 1568 982 1571
rect 1054 1568 1062 1571
rect 1538 1568 1541 1572
rect 2546 1568 2549 1572
rect 2738 1568 2740 1572
rect 3002 1568 3004 1572
rect 3462 1568 3473 1571
rect 4978 1568 4980 1572
rect 5178 1568 5180 1572
rect 54 1558 62 1561
rect 142 1558 153 1561
rect 370 1558 374 1562
rect 22 1548 38 1551
rect 46 1548 54 1551
rect 278 1548 302 1551
rect 346 1548 369 1551
rect 386 1548 401 1551
rect 622 1551 625 1561
rect 658 1558 662 1562
rect 750 1558 761 1561
rect 838 1558 846 1561
rect 1078 1558 1089 1561
rect 1646 1558 1655 1562
rect 1854 1558 1865 1561
rect 2070 1558 2081 1561
rect 2418 1558 2422 1562
rect 2430 1558 2441 1561
rect 3342 1561 3345 1568
rect 3462 1566 3466 1568
rect 3334 1558 3345 1561
rect 606 1548 625 1551
rect 742 1548 750 1551
rect 806 1551 810 1554
rect 798 1548 810 1551
rect 866 1548 873 1551
rect 990 1551 994 1554
rect 1646 1552 1649 1558
rect 986 1548 994 1551
rect 1102 1548 1118 1551
rect 10 1538 17 1541
rect 26 1538 33 1541
rect 70 1538 97 1541
rect 182 1541 185 1548
rect 150 1538 169 1541
rect 174 1538 185 1541
rect 334 1538 342 1541
rect 726 1538 729 1548
rect 1022 1541 1025 1548
rect 1022 1538 1033 1541
rect 1062 1538 1070 1541
rect 1086 1538 1089 1548
rect 1502 1548 1510 1551
rect 1614 1548 1622 1551
rect 1710 1548 1721 1551
rect 1942 1548 1950 1551
rect 1958 1548 1966 1551
rect 2094 1548 2102 1551
rect 2126 1548 2153 1551
rect 2366 1551 2370 1554
rect 2366 1548 2374 1551
rect 2382 1548 2417 1551
rect 2450 1548 2473 1551
rect 2902 1548 2918 1551
rect 3038 1551 3042 1553
rect 3034 1548 3042 1551
rect 3070 1548 3078 1551
rect 3090 1548 3097 1551
rect 1710 1538 1713 1548
rect 1898 1538 1921 1541
rect 1990 1538 1993 1548
rect 2038 1538 2041 1548
rect 3374 1548 3385 1551
rect 3422 1551 3426 1554
rect 3422 1548 3449 1551
rect 2074 1538 2081 1541
rect 2202 1538 2209 1541
rect 2334 1538 2348 1541
rect 3354 1538 3361 1541
rect 3446 1538 3449 1548
rect 3714 1548 3721 1551
rect 3914 1548 3921 1551
rect 4542 1548 4553 1551
rect 4558 1548 4577 1551
rect 4586 1548 4609 1551
rect 4718 1551 4722 1554
rect 4718 1548 4729 1551
rect 4814 1548 4825 1551
rect 5066 1548 5081 1551
rect 5086 1548 5094 1551
rect 5118 1548 5137 1551
rect 5142 1548 5158 1551
rect 3694 1538 3713 1541
rect 3982 1538 3998 1541
rect 4486 1541 4489 1548
rect 4542 1542 4545 1548
rect 4486 1538 4497 1541
rect 4614 1538 4622 1541
rect 4630 1538 4641 1541
rect 4726 1538 4729 1548
rect 4814 1542 4817 1548
rect 5038 1541 5041 1548
rect 5038 1538 5049 1541
rect 5054 1538 5062 1541
rect 770 1528 777 1531
rect 1070 1528 1073 1538
rect 1122 1528 1129 1531
rect 1754 1528 1761 1531
rect 1950 1528 1961 1531
rect 2194 1528 2201 1531
rect 2526 1531 2530 1533
rect 2518 1528 2530 1531
rect 3286 1528 3297 1531
rect 3710 1528 3713 1538
rect 4926 1528 4929 1538
rect 226 1518 233 1521
rect 250 1518 271 1521
rect 506 1518 508 1522
rect 2850 1518 2852 1522
rect 2956 1518 2958 1522
rect 3406 1518 3414 1521
rect 4114 1518 4116 1522
rect 4266 1518 4268 1522
rect 4322 1518 4324 1522
rect 4378 1518 4380 1522
rect 4738 1518 4739 1522
rect 4858 1518 4860 1522
rect 5266 1518 5268 1522
rect 856 1503 858 1507
rect 862 1503 865 1507
rect 869 1503 872 1507
rect 1872 1503 1874 1507
rect 1878 1503 1881 1507
rect 1885 1503 1888 1507
rect 2904 1503 2906 1507
rect 2910 1503 2913 1507
rect 2917 1503 2920 1507
rect 3928 1503 3930 1507
rect 3934 1503 3937 1507
rect 3941 1503 3944 1507
rect 4952 1503 4954 1507
rect 4958 1503 4961 1507
rect 4965 1503 4968 1507
rect 284 1488 286 1492
rect 532 1488 534 1492
rect 588 1488 590 1492
rect 717 1488 718 1492
rect 1444 1488 1446 1492
rect 1834 1488 1835 1492
rect 1989 1488 1990 1492
rect 2298 1488 2299 1492
rect 2340 1488 2342 1492
rect 2612 1488 2614 1492
rect 3725 1488 3726 1492
rect 4829 1488 4830 1492
rect 4934 1488 4942 1491
rect 5013 1488 5014 1492
rect 14 1478 25 1481
rect 66 1478 73 1482
rect 158 1478 166 1481
rect 350 1478 366 1481
rect 1222 1478 1230 1482
rect 2774 1478 2786 1481
rect 70 1472 73 1478
rect 46 1468 57 1471
rect 166 1471 169 1478
rect 46 1462 49 1468
rect 150 1461 153 1471
rect 166 1468 177 1471
rect 198 1468 209 1471
rect 326 1468 345 1471
rect 486 1468 505 1471
rect 734 1468 745 1471
rect 778 1468 785 1471
rect 1158 1468 1161 1478
rect 1222 1472 1225 1478
rect 1302 1471 1305 1478
rect 1262 1468 1273 1471
rect 1302 1468 1313 1471
rect 1402 1468 1417 1471
rect 1586 1468 1587 1472
rect 1622 1471 1626 1474
rect 1622 1468 1633 1471
rect 1678 1468 1697 1471
rect 1842 1468 1849 1471
rect 1910 1471 1913 1478
rect 2782 1477 2786 1478
rect 3190 1478 3198 1481
rect 3426 1478 3449 1481
rect 3578 1478 3593 1481
rect 3598 1478 3606 1481
rect 3638 1478 3646 1481
rect 3954 1478 3961 1481
rect 1902 1468 1913 1471
rect 206 1462 209 1468
rect 150 1458 182 1461
rect 326 1458 329 1468
rect 734 1462 737 1468
rect 398 1458 422 1461
rect 494 1458 502 1461
rect 678 1458 694 1461
rect 750 1458 758 1461
rect 1242 1458 1257 1461
rect 1302 1458 1310 1461
rect 1326 1458 1334 1461
rect 1734 1458 1742 1461
rect 1782 1458 1801 1461
rect 1942 1461 1945 1471
rect 2034 1468 2041 1471
rect 2118 1468 2126 1471
rect 2306 1468 2313 1471
rect 2358 1468 2366 1471
rect 2414 1468 2449 1471
rect 2490 1468 2497 1471
rect 2734 1468 2753 1471
rect 2758 1468 2769 1471
rect 2926 1468 2929 1478
rect 3510 1468 3545 1471
rect 3606 1468 3617 1471
rect 3670 1468 3681 1471
rect 3702 1468 3710 1471
rect 4218 1468 4219 1472
rect 4382 1468 4401 1471
rect 4434 1468 4449 1471
rect 1942 1458 1953 1461
rect 2042 1458 2049 1461
rect 2126 1458 2145 1461
rect 2758 1462 2761 1468
rect 2498 1458 2505 1461
rect 3174 1458 3182 1461
rect 3206 1461 3209 1468
rect 3606 1462 3609 1468
rect 3678 1462 3681 1468
rect 3198 1458 3209 1461
rect 4478 1462 4481 1471
rect 4542 1468 4553 1471
rect 4742 1468 4761 1471
rect 4862 1468 4881 1471
rect 4954 1468 4964 1471
rect 5066 1468 5073 1471
rect 4542 1462 4545 1468
rect 4078 1458 4086 1461
rect 4334 1458 4353 1461
rect 4518 1458 4529 1461
rect 4894 1458 4897 1468
rect 4918 1458 4926 1461
rect 5054 1458 5065 1461
rect 5134 1458 5158 1461
rect 5186 1458 5193 1461
rect 222 1456 226 1458
rect 74 1448 81 1451
rect 130 1449 132 1453
rect 214 1448 225 1451
rect 694 1448 713 1451
rect 1362 1448 1364 1452
rect 1650 1448 1652 1452
rect 4422 1448 4430 1451
rect 4866 1448 4873 1451
rect 4982 1448 4993 1451
rect 694 1442 697 1448
rect 3450 1438 3457 1441
rect 4644 1438 4646 1442
rect 93 1418 94 1422
rect 1482 1418 1483 1422
rect 2386 1418 2390 1422
rect 2546 1418 2550 1422
rect 4724 1418 4726 1422
rect 344 1403 346 1407
rect 350 1403 353 1407
rect 357 1403 360 1407
rect 1368 1403 1370 1407
rect 1374 1403 1377 1407
rect 1381 1403 1384 1407
rect 2392 1403 2394 1407
rect 2398 1403 2401 1407
rect 2405 1403 2408 1407
rect 3416 1403 3418 1407
rect 3422 1403 3425 1407
rect 3429 1403 3432 1407
rect 4440 1403 4442 1407
rect 4446 1403 4449 1407
rect 4453 1403 4456 1407
rect 162 1388 164 1392
rect 1762 1388 1764 1392
rect 1986 1388 1990 1392
rect 2178 1388 2179 1392
rect 2301 1388 2302 1392
rect 2794 1388 2795 1392
rect 5114 1388 5115 1392
rect 1834 1378 1836 1382
rect 2074 1378 2076 1382
rect 2682 1378 2684 1382
rect 14 1368 30 1371
rect 42 1368 49 1371
rect 850 1368 881 1371
rect 954 1368 961 1371
rect 1109 1368 1110 1372
rect 4650 1368 4652 1372
rect 4706 1368 4708 1372
rect 4762 1368 4764 1372
rect 5006 1368 5033 1371
rect 5242 1368 5257 1371
rect 30 1358 38 1361
rect 406 1358 414 1361
rect 510 1358 529 1361
rect 822 1361 825 1368
rect 822 1358 833 1361
rect 854 1358 870 1361
rect 1078 1358 1097 1361
rect 2322 1358 2329 1361
rect 2358 1358 2369 1361
rect 2806 1358 2817 1361
rect 2842 1358 2846 1362
rect 2906 1358 2926 1361
rect 2942 1361 2945 1368
rect 2942 1358 2953 1361
rect 4510 1361 4513 1368
rect 5006 1362 5010 1364
rect 4510 1358 4521 1361
rect 5018 1358 5025 1361
rect 5066 1358 5073 1361
rect 5126 1358 5137 1361
rect 5230 1361 5233 1368
rect 5222 1358 5233 1361
rect 206 1348 217 1351
rect 530 1348 537 1351
rect 662 1348 670 1351
rect 1070 1351 1073 1358
rect 1070 1348 1081 1351
rect 1110 1348 1126 1351
rect 214 1342 217 1348
rect 126 1338 145 1341
rect 190 1338 209 1341
rect 350 1341 353 1348
rect 326 1338 353 1341
rect 462 1341 465 1348
rect 462 1338 473 1341
rect 502 1338 513 1341
rect 586 1338 593 1341
rect 798 1338 817 1341
rect 918 1341 921 1348
rect 910 1338 921 1341
rect 970 1338 972 1342
rect 1054 1341 1057 1348
rect 2126 1348 2134 1351
rect 2202 1348 2209 1351
rect 2302 1348 2318 1351
rect 2418 1348 2449 1351
rect 2742 1348 2761 1351
rect 2878 1348 2897 1351
rect 3194 1348 3201 1351
rect 1054 1338 1065 1341
rect 1862 1338 1870 1341
rect 2134 1338 2142 1341
rect 2150 1338 2169 1341
rect 2710 1338 2718 1341
rect 2974 1338 2982 1341
rect 3102 1341 3105 1348
rect 3350 1348 3358 1351
rect 3434 1348 3441 1351
rect 3846 1351 3850 1353
rect 3838 1348 3850 1351
rect 3890 1348 3905 1351
rect 4086 1348 4102 1351
rect 4566 1348 4585 1351
rect 4622 1348 4630 1351
rect 5090 1348 5113 1351
rect 3066 1338 3073 1341
rect 3086 1338 3105 1341
rect 3614 1338 3633 1341
rect 3934 1338 3962 1341
rect 4174 1338 4185 1341
rect 4206 1338 4214 1341
rect 4326 1338 4334 1341
rect 4566 1338 4569 1348
rect 4622 1338 4633 1341
rect 5094 1338 5102 1341
rect 5162 1338 5169 1341
rect 126 1328 134 1331
rect 246 1328 262 1331
rect 314 1328 318 1332
rect 590 1328 593 1338
rect 898 1328 902 1332
rect 2922 1328 2934 1331
rect 2974 1328 2977 1338
rect 2986 1328 2990 1332
rect 3414 1328 3433 1331
rect 3806 1328 3817 1331
rect 4326 1328 4329 1338
rect 5182 1332 5185 1338
rect 4542 1328 4558 1331
rect 5178 1328 5185 1332
rect 493 1318 494 1322
rect 714 1318 716 1322
rect 770 1318 772 1322
rect 2570 1318 2572 1322
rect 2626 1318 2628 1322
rect 3058 1318 3059 1322
rect 3414 1321 3417 1328
rect 3406 1318 3417 1321
rect 4946 1318 4948 1322
rect 5250 1318 5257 1321
rect 856 1303 858 1307
rect 862 1303 865 1307
rect 869 1303 872 1307
rect 1872 1303 1874 1307
rect 1878 1303 1881 1307
rect 1885 1303 1888 1307
rect 2904 1303 2906 1307
rect 2910 1303 2913 1307
rect 2917 1303 2920 1307
rect 3928 1303 3930 1307
rect 3934 1303 3937 1307
rect 3941 1303 3944 1307
rect 4952 1303 4954 1307
rect 4958 1303 4961 1307
rect 4965 1303 4968 1307
rect 69 1288 70 1292
rect 394 1288 395 1292
rect 562 1288 564 1292
rect 642 1288 644 1292
rect 1426 1288 1428 1292
rect 2634 1288 2636 1292
rect 4692 1288 4694 1292
rect 4874 1288 4876 1292
rect 4986 1288 5001 1291
rect 5146 1288 5147 1292
rect 5226 1288 5233 1291
rect 298 1278 305 1281
rect 498 1278 502 1282
rect 966 1278 977 1281
rect 1358 1278 1374 1281
rect 2694 1278 2710 1281
rect 4126 1278 4138 1281
rect 4258 1278 4265 1281
rect 78 1268 89 1271
rect 158 1268 169 1271
rect 322 1268 342 1271
rect 372 1268 385 1271
rect 950 1271 953 1278
rect 882 1268 897 1271
rect 902 1268 913 1271
rect 918 1268 937 1271
rect 942 1268 953 1271
rect 966 1272 969 1278
rect 1062 1271 1065 1278
rect 3262 1277 3266 1278
rect 1070 1271 1074 1272
rect 1062 1268 1074 1271
rect 1090 1268 1097 1271
rect 1346 1268 1353 1271
rect 1454 1268 1462 1271
rect 1482 1268 1497 1271
rect 902 1262 905 1268
rect 1558 1262 1561 1271
rect 1582 1268 1590 1271
rect 1674 1268 1681 1271
rect 78 1258 89 1261
rect 410 1258 417 1261
rect 518 1258 526 1261
rect 946 1258 961 1261
rect 1210 1258 1217 1261
rect 1234 1258 1241 1261
rect 1314 1258 1321 1261
rect 1642 1258 1649 1261
rect 2042 1258 2049 1261
rect 2062 1261 2065 1271
rect 2098 1268 2105 1271
rect 2146 1268 2153 1271
rect 2306 1268 2313 1271
rect 2494 1271 2498 1274
rect 3366 1272 3370 1274
rect 2486 1268 2498 1271
rect 2758 1268 2769 1271
rect 2966 1268 2977 1271
rect 3130 1268 3137 1271
rect 3446 1268 3454 1271
rect 3558 1268 3566 1271
rect 3594 1268 3601 1271
rect 3606 1268 3617 1271
rect 3650 1268 3665 1271
rect 3682 1268 3689 1271
rect 3734 1271 3738 1274
rect 4094 1271 4097 1278
rect 4134 1277 4138 1278
rect 4646 1272 4649 1281
rect 4786 1278 4793 1282
rect 4790 1272 4793 1278
rect 3726 1268 3738 1271
rect 4078 1268 4097 1271
rect 4421 1268 4422 1272
rect 2062 1258 2070 1261
rect 2142 1258 2153 1261
rect 2314 1258 2321 1261
rect 2758 1262 2761 1268
rect 2710 1258 2737 1261
rect 2814 1261 2817 1268
rect 2966 1262 2969 1268
rect 2814 1258 2825 1261
rect 2830 1258 2841 1261
rect 3122 1258 3145 1261
rect 3614 1262 3617 1268
rect 3562 1258 3569 1261
rect 3678 1258 3686 1261
rect 4662 1262 4665 1271
rect 4850 1268 4857 1271
rect 5294 1268 5302 1271
rect 3950 1258 3958 1261
rect 4018 1258 4025 1261
rect 4110 1258 4121 1261
rect 4246 1258 4254 1261
rect 4266 1258 4281 1261
rect 4374 1258 4386 1261
rect 4514 1258 4521 1261
rect 5082 1258 5100 1261
rect 5186 1258 5193 1261
rect 5198 1258 5206 1261
rect 5262 1258 5270 1261
rect 78 1252 81 1258
rect 286 1248 294 1251
rect 706 1248 713 1251
rect 814 1248 825 1251
rect 894 1248 905 1251
rect 1166 1248 1185 1251
rect 1226 1248 1233 1251
rect 1518 1251 1521 1258
rect 4382 1257 4386 1258
rect 4150 1252 4154 1257
rect 1518 1248 1529 1251
rect 1554 1248 1561 1251
rect 2738 1248 2742 1252
rect 2986 1248 2993 1251
rect 3078 1248 3105 1251
rect 4830 1251 4833 1258
rect 4822 1248 4833 1251
rect 5258 1248 5262 1252
rect 346 1238 369 1241
rect 1110 1238 1142 1241
rect 2178 1238 2185 1241
rect 2218 1238 2220 1242
rect 2451 1238 2454 1242
rect 3158 1238 3169 1241
rect 4748 1238 4750 1242
rect 1197 1218 1198 1222
rect 1298 1218 1299 1222
rect 2922 1218 2937 1221
rect 344 1203 346 1207
rect 350 1203 353 1207
rect 357 1203 360 1207
rect 1368 1203 1370 1207
rect 1374 1203 1377 1207
rect 1381 1203 1384 1207
rect 2392 1203 2394 1207
rect 2398 1203 2401 1207
rect 2405 1203 2408 1207
rect 3416 1203 3418 1207
rect 3422 1203 3425 1207
rect 3429 1203 3432 1207
rect 4440 1203 4442 1207
rect 4446 1203 4449 1207
rect 4453 1203 4456 1207
rect 50 1188 54 1192
rect 213 1188 214 1192
rect 610 1188 611 1192
rect 714 1188 715 1192
rect 1756 1188 1758 1192
rect 2138 1188 2139 1192
rect 2290 1188 2292 1192
rect 2370 1188 2372 1192
rect 2522 1188 2524 1192
rect 2709 1188 2710 1192
rect 2906 1188 2921 1191
rect 3926 1188 3934 1191
rect 4844 1188 4846 1192
rect 4933 1188 4934 1192
rect 5205 1188 5206 1192
rect 2418 1178 2425 1181
rect 110 1168 142 1171
rect 174 1168 185 1171
rect 514 1168 516 1172
rect 762 1168 769 1171
rect 4878 1168 4894 1171
rect 174 1162 177 1168
rect 182 1158 201 1161
rect 658 1158 665 1161
rect 1890 1158 1902 1161
rect 2150 1158 2161 1161
rect 22 1148 57 1151
rect 90 1148 97 1151
rect 214 1148 238 1151
rect 462 1148 470 1151
rect 570 1148 577 1151
rect 678 1151 681 1158
rect 678 1148 689 1151
rect 774 1142 777 1151
rect 1414 1148 1438 1151
rect 1718 1148 1726 1151
rect 1994 1148 2012 1151
rect 2102 1148 2113 1151
rect 2578 1148 2601 1151
rect 2606 1148 2622 1151
rect 2662 1148 2673 1151
rect 1718 1146 1722 1148
rect 26 1138 33 1141
rect 222 1138 230 1141
rect 414 1138 425 1141
rect 542 1138 550 1141
rect 574 1138 585 1141
rect 590 1138 598 1141
rect 678 1138 689 1141
rect 830 1138 857 1141
rect 1426 1138 1433 1141
rect 1674 1138 1681 1141
rect 1774 1138 1777 1148
rect 2670 1142 2673 1148
rect 2820 1148 2822 1152
rect 2946 1148 2961 1151
rect 3146 1148 3161 1151
rect 2106 1138 2113 1141
rect 2118 1138 2126 1141
rect 2238 1138 2246 1141
rect 2318 1138 2326 1141
rect 2334 1138 2353 1141
rect 2402 1138 2425 1141
rect 2550 1138 2561 1141
rect 2582 1138 2590 1141
rect 2630 1138 2638 1141
rect 2686 1141 2689 1148
rect 3442 1148 3449 1151
rect 3494 1151 3497 1161
rect 4010 1158 4014 1162
rect 4022 1158 4030 1161
rect 4366 1158 4374 1161
rect 4910 1158 4921 1161
rect 5154 1158 5161 1161
rect 3494 1148 3513 1151
rect 3518 1148 3537 1151
rect 3598 1151 3601 1158
rect 3598 1148 3609 1151
rect 3726 1148 3737 1151
rect 3742 1148 3761 1151
rect 3806 1148 3817 1151
rect 3822 1148 3833 1151
rect 3726 1142 3729 1148
rect 3830 1142 3833 1148
rect 3986 1148 4009 1151
rect 4138 1148 4145 1151
rect 4262 1151 4265 1158
rect 4262 1148 4289 1151
rect 4894 1151 4898 1154
rect 4894 1148 4902 1151
rect 4934 1148 4969 1151
rect 5054 1148 5078 1151
rect 5174 1148 5190 1151
rect 5294 1148 5302 1151
rect 2678 1138 2689 1141
rect 2762 1138 2769 1141
rect 3045 1138 3046 1142
rect 3214 1138 3233 1141
rect 3590 1138 3606 1141
rect 3766 1138 3774 1141
rect 3790 1138 3809 1141
rect 4138 1138 4153 1141
rect 4302 1138 4337 1141
rect 4710 1138 4722 1141
rect 4966 1141 4969 1148
rect 4966 1138 4982 1141
rect 414 1132 417 1138
rect 574 1132 577 1138
rect 590 1128 593 1138
rect 1798 1132 1801 1138
rect 766 1128 777 1131
rect 1798 1128 1806 1132
rect 1878 1128 1886 1131
rect 2070 1128 2081 1131
rect 2118 1128 2121 1138
rect 2422 1128 2425 1138
rect 2454 1128 2457 1138
rect 3610 1128 3617 1131
rect 3790 1128 3793 1138
rect 4046 1132 4049 1138
rect 4042 1128 4049 1132
rect 4158 1128 4174 1131
rect 4230 1131 4233 1138
rect 4230 1128 4241 1131
rect 5146 1128 5153 1131
rect 378 1118 380 1122
rect 874 1118 876 1122
rect 930 1118 932 1122
rect 1101 1118 1102 1122
rect 1370 1118 1385 1121
rect 1492 1118 1494 1122
rect 1538 1118 1540 1122
rect 1610 1118 1612 1122
rect 2258 1118 2259 1122
rect 2338 1118 2339 1122
rect 4596 1118 4598 1122
rect 5306 1118 5313 1121
rect 5310 1108 5313 1118
rect 856 1103 858 1107
rect 862 1103 865 1107
rect 869 1103 872 1107
rect 1872 1103 1874 1107
rect 1878 1103 1881 1107
rect 1885 1103 1888 1107
rect 2904 1103 2906 1107
rect 2910 1103 2913 1107
rect 2917 1103 2920 1107
rect 3928 1103 3930 1107
rect 3934 1103 3937 1107
rect 3941 1103 3944 1107
rect 4952 1103 4954 1107
rect 4958 1103 4961 1107
rect 4965 1103 4968 1107
rect 85 1088 86 1092
rect 181 1088 182 1092
rect 908 1088 910 1092
rect 1389 1088 1390 1092
rect 2108 1088 2110 1092
rect 2386 1088 2388 1092
rect 2589 1088 2590 1092
rect 2717 1088 2718 1092
rect 4430 1088 4438 1091
rect 4636 1088 4638 1092
rect 4692 1088 4694 1092
rect 5157 1088 5158 1092
rect 5226 1088 5241 1091
rect 146 1078 161 1081
rect 734 1078 745 1081
rect 1242 1078 1249 1081
rect 3182 1078 3193 1081
rect 3614 1078 3622 1081
rect 3934 1078 3961 1081
rect 4354 1078 4361 1082
rect 4534 1078 4542 1081
rect 5178 1078 5185 1081
rect 5202 1078 5209 1081
rect 734 1072 737 1078
rect 94 1068 105 1071
rect 134 1068 150 1071
rect 190 1068 209 1071
rect 382 1061 385 1071
rect 430 1068 441 1071
rect 566 1068 577 1071
rect 614 1068 622 1071
rect 666 1068 673 1071
rect 766 1068 774 1071
rect 926 1068 934 1071
rect 958 1068 977 1071
rect 1102 1068 1110 1071
rect 1190 1068 1209 1071
rect 1294 1068 1321 1071
rect 1402 1068 1412 1071
rect 1934 1068 1961 1071
rect 2350 1071 2353 1078
rect 2340 1068 2353 1071
rect 566 1062 569 1068
rect 382 1058 414 1061
rect 582 1058 593 1061
rect 630 1058 638 1061
rect 662 1058 678 1061
rect 1106 1058 1113 1061
rect 1158 1058 1177 1061
rect 1198 1058 1206 1061
rect 1330 1058 1342 1061
rect 1350 1058 1385 1061
rect 1518 1058 1550 1061
rect 1594 1058 1609 1061
rect 1846 1058 1857 1061
rect 1918 1058 1937 1061
rect 1942 1058 1953 1061
rect 2198 1061 2201 1068
rect 2166 1058 2201 1061
rect 2242 1058 2250 1061
rect 2414 1061 2417 1071
rect 2518 1068 2529 1071
rect 2534 1068 2561 1071
rect 2622 1068 2633 1071
rect 2526 1062 2529 1068
rect 2622 1062 2625 1068
rect 2742 1071 2745 1078
rect 2742 1068 2756 1071
rect 3610 1068 3617 1071
rect 3878 1071 3882 1074
rect 4358 1072 4361 1078
rect 3878 1068 3889 1071
rect 3974 1068 3982 1071
rect 3998 1068 4006 1071
rect 4118 1068 4130 1071
rect 4486 1068 4494 1071
rect 4510 1068 4526 1071
rect 4806 1071 4810 1074
rect 4806 1068 4817 1071
rect 4910 1068 4918 1071
rect 4994 1068 5001 1071
rect 2414 1058 2449 1061
rect 2454 1058 2473 1061
rect 2834 1058 2841 1061
rect 2882 1058 2905 1061
rect 2930 1058 2937 1061
rect 3214 1058 3225 1061
rect 3738 1058 3753 1061
rect 3894 1058 3921 1061
rect 3982 1058 4009 1061
rect 4238 1061 4241 1068
rect 4230 1058 4241 1061
rect 4298 1058 4305 1061
rect 4374 1058 4382 1061
rect 4542 1058 4561 1061
rect 4566 1058 4585 1061
rect 4590 1058 4598 1061
rect 5002 1058 5025 1061
rect 582 1052 585 1058
rect 1054 1048 1081 1051
rect 1090 1048 1094 1052
rect 1382 1048 1385 1058
rect 1846 1052 1849 1058
rect 1942 1052 1945 1058
rect 2246 1056 2250 1058
rect 1862 1048 1873 1051
rect 2142 1048 2153 1051
rect 2162 1048 2166 1052
rect 2454 1048 2457 1058
rect 2822 1048 2830 1051
rect 242 1038 244 1042
rect 1474 1038 1481 1041
rect 4397 1038 4398 1042
rect 1014 1028 1017 1038
rect 1478 1028 1481 1038
rect 482 1018 483 1022
rect 682 1018 683 1022
rect 794 1018 796 1022
rect 1229 1018 1230 1022
rect 1450 1018 1451 1022
rect 2509 1018 2510 1022
rect 344 1003 346 1007
rect 350 1003 353 1007
rect 357 1003 360 1007
rect 1368 1003 1370 1007
rect 1374 1003 1377 1007
rect 1381 1003 1384 1007
rect 2392 1003 2394 1007
rect 2398 1003 2401 1007
rect 2405 1003 2408 1007
rect 3416 1003 3418 1007
rect 3422 1003 3425 1007
rect 3429 1003 3432 1007
rect 4440 1003 4442 1007
rect 4446 1003 4449 1007
rect 4453 1003 4456 1007
rect 290 988 291 992
rect 437 988 438 992
rect 2106 988 2107 992
rect 2740 988 2742 992
rect 3146 988 3147 992
rect 4669 988 4670 992
rect 4826 988 4830 992
rect 5020 988 5022 992
rect 845 978 846 982
rect 3122 978 3123 982
rect 242 968 244 972
rect 370 968 377 971
rect 466 968 489 971
rect 506 968 513 971
rect 994 968 1009 971
rect 1204 968 1206 972
rect 2882 968 2897 971
rect 3674 968 3689 971
rect 4602 968 4609 971
rect 4749 968 4750 972
rect 5100 968 5102 972
rect 142 951 145 961
rect 326 958 361 961
rect 614 961 617 968
rect 606 958 617 961
rect 902 958 929 961
rect 2398 958 2414 961
rect 2518 958 2526 961
rect 2990 956 2994 958
rect 126 948 145 951
rect 206 948 222 951
rect 294 948 313 951
rect 318 948 329 951
rect 442 948 457 951
rect 694 948 710 951
rect 718 948 726 951
rect 102 938 121 941
rect 182 938 190 941
rect 278 941 281 948
rect 278 938 289 941
rect 570 938 593 941
rect 598 938 609 941
rect 614 938 622 941
rect 642 938 652 941
rect 678 938 681 948
rect 846 948 886 951
rect 1126 948 1137 951
rect 1150 948 1161 951
rect 1250 948 1257 951
rect 702 938 710 941
rect 858 938 881 941
rect 902 938 905 948
rect 1134 942 1137 948
rect 1558 951 1562 954
rect 1558 948 1566 951
rect 1614 948 1622 951
rect 1634 948 1649 951
rect 1654 948 1681 951
rect 1686 948 1694 951
rect 938 938 948 941
rect 1030 938 1041 941
rect 1098 938 1105 941
rect 1414 941 1417 948
rect 1414 938 1428 941
rect 1622 938 1657 941
rect 1842 938 1857 941
rect 1934 941 1937 948
rect 2086 948 2102 951
rect 2122 948 2129 951
rect 2454 948 2489 951
rect 1934 938 1945 941
rect 1950 938 1962 941
rect 182 928 185 938
rect 614 928 617 938
rect 1038 932 1041 938
rect 1142 928 1150 931
rect 1494 928 1505 931
rect 1582 931 1585 938
rect 1574 928 1585 931
rect 1618 928 1625 931
rect 1758 931 1761 938
rect 1958 936 1962 938
rect 2430 941 2433 948
rect 2486 942 2489 948
rect 3086 948 3097 951
rect 3174 951 3177 961
rect 3434 958 3449 961
rect 3546 958 3550 962
rect 3174 948 3193 951
rect 3214 948 3222 951
rect 3286 948 3297 951
rect 3310 948 3321 951
rect 3526 948 3534 951
rect 3558 951 3561 961
rect 3662 958 3673 961
rect 3750 958 3758 961
rect 3918 958 3934 961
rect 4286 958 4297 961
rect 4442 958 4465 961
rect 4550 958 4558 961
rect 4954 958 4961 961
rect 3558 948 3569 951
rect 3606 948 3617 951
rect 4014 948 4033 951
rect 4038 948 4046 951
rect 4422 948 4433 951
rect 4466 948 4473 951
rect 4614 948 4625 951
rect 4718 948 4726 951
rect 4750 948 4774 951
rect 4982 948 4990 951
rect 3086 942 3089 948
rect 3294 942 3297 948
rect 2430 938 2441 941
rect 2530 938 2545 941
rect 3566 941 3569 948
rect 3614 942 3617 948
rect 3566 938 3577 941
rect 4046 938 4062 941
rect 4078 938 4086 941
rect 4146 938 4161 941
rect 4178 938 4185 941
rect 4358 938 4374 941
rect 4390 938 4409 941
rect 4494 938 4497 948
rect 4614 942 4617 948
rect 4590 938 4598 941
rect 4758 938 4766 941
rect 4790 938 4801 941
rect 5042 938 5057 941
rect 5118 938 5126 941
rect 5134 938 5146 941
rect 1746 928 1761 931
rect 2054 931 2057 938
rect 2054 928 2065 931
rect 2230 931 2234 936
rect 2218 928 2234 931
rect 2246 931 2250 933
rect 2246 928 2257 931
rect 2498 928 2505 931
rect 3346 928 3361 931
rect 3426 928 3441 931
rect 3446 928 3457 931
rect 4030 931 4033 938
rect 3918 928 3945 931
rect 4018 928 4033 931
rect 4046 928 4049 938
rect 4190 928 4198 931
rect 4406 928 4409 938
rect 5142 936 5146 938
rect 5262 932 5265 938
rect 4610 928 4625 931
rect 5262 928 5270 932
rect 526 918 534 921
rect 1237 918 1238 922
rect 1494 918 1497 928
rect 1642 918 1649 921
rect 1820 918 1822 922
rect 1916 918 1918 922
rect 4233 918 4246 921
rect 856 903 858 907
rect 862 903 865 907
rect 869 903 872 907
rect 1872 903 1874 907
rect 1878 903 1881 907
rect 1885 903 1888 907
rect 2904 903 2906 907
rect 2910 903 2913 907
rect 2917 903 2920 907
rect 3928 903 3930 907
rect 3934 903 3937 907
rect 3941 903 3944 907
rect 4952 903 4954 907
rect 4958 903 4961 907
rect 4965 903 4968 907
rect 394 888 395 892
rect 1484 888 1486 892
rect 1588 888 1590 892
rect 1884 888 1886 892
rect 1956 888 1958 892
rect 2092 888 2094 892
rect 2126 888 2134 891
rect 3054 888 3065 891
rect 3649 888 3670 891
rect 4325 888 4326 892
rect 4882 888 4883 892
rect 5005 888 5006 892
rect 5030 888 5041 891
rect 5146 888 5148 892
rect 5202 888 5204 892
rect 3054 882 3057 888
rect 518 878 529 881
rect 890 878 897 881
rect 902 878 910 881
rect 1074 878 1081 882
rect 3010 878 3017 881
rect 3710 878 3718 881
rect 3750 878 3769 881
rect 5030 882 5033 888
rect 4546 878 4553 881
rect 4682 878 4694 881
rect 4782 878 4790 881
rect 4806 878 4814 881
rect 1078 872 1081 878
rect 370 868 382 871
rect 450 868 481 871
rect 554 868 569 871
rect 574 868 601 871
rect 630 868 641 871
rect 678 868 686 871
rect 934 868 945 871
rect 958 868 966 871
rect 1106 868 1121 871
rect 1170 868 1185 871
rect 74 858 81 861
rect 534 861 537 868
rect 942 862 945 868
rect 534 858 545 861
rect 658 858 665 861
rect 670 858 686 861
rect 950 858 969 861
rect 990 858 993 868
rect 1262 861 1265 871
rect 1354 868 1369 871
rect 1554 868 1561 871
rect 1262 858 1281 861
rect 1438 858 1454 861
rect 1702 861 1705 871
rect 1846 871 1850 874
rect 1846 868 1857 871
rect 1922 868 1929 871
rect 1986 868 1993 871
rect 1998 868 2014 871
rect 2058 868 2065 871
rect 2178 868 2185 871
rect 2198 868 2214 871
rect 2278 868 2286 871
rect 2322 868 2329 871
rect 2350 868 2358 871
rect 2460 868 2481 871
rect 2506 868 2513 871
rect 3294 868 3302 871
rect 3414 868 3422 871
rect 3442 868 3449 871
rect 3482 868 3497 871
rect 4050 868 4060 871
rect 1670 858 1705 861
rect 2318 858 2337 861
rect 2342 858 2366 861
rect 2374 858 2382 861
rect 2794 858 2801 861
rect 2982 858 2990 861
rect 3210 858 3217 861
rect 3358 858 3377 861
rect 3386 858 3401 861
rect 3570 858 3577 861
rect 3674 858 3689 861
rect 3734 858 3753 861
rect 3858 858 3865 861
rect 3894 858 3910 861
rect 3958 858 3966 861
rect 4098 858 4105 861
rect 4178 858 4185 861
rect 4382 861 4385 871
rect 4412 868 4414 872
rect 4490 868 4497 871
rect 4510 868 4526 871
rect 4382 858 4394 861
rect 4478 861 4481 868
rect 4754 868 4761 871
rect 4774 868 4782 871
rect 4830 868 4857 871
rect 4470 858 4481 861
rect 4650 858 4657 861
rect 4782 858 4793 861
rect 4942 858 4977 861
rect 638 848 657 851
rect 1054 848 1062 851
rect 1386 848 1388 852
rect 2038 851 2041 858
rect 2030 848 2041 851
rect 2382 848 2406 851
rect 3302 851 3305 858
rect 3302 848 3313 851
rect 3398 848 3401 858
rect 3694 851 3697 858
rect 4390 856 4394 858
rect 3694 848 3705 851
rect 3926 851 3930 854
rect 3902 848 3930 851
rect 4558 848 4569 851
rect 4906 848 4910 852
rect 4974 848 4977 858
rect 5018 848 5025 851
rect 1827 838 1830 842
rect 2126 838 2134 841
rect 1330 828 1331 832
rect 1253 818 1254 822
rect 2620 818 2622 822
rect 2772 818 2774 822
rect 344 803 346 807
rect 350 803 353 807
rect 357 803 360 807
rect 1368 803 1370 807
rect 1374 803 1377 807
rect 1381 803 1384 807
rect 2392 803 2394 807
rect 2398 803 2401 807
rect 2405 803 2408 807
rect 3416 803 3418 807
rect 3422 803 3425 807
rect 3429 803 3432 807
rect 4440 803 4442 807
rect 4446 803 4449 807
rect 4453 803 4456 807
rect 636 788 638 792
rect 1098 788 1099 792
rect 1844 788 1846 792
rect 2357 788 2358 792
rect 2802 788 2804 792
rect 3612 788 3614 792
rect 4365 788 4366 792
rect 4770 788 4771 792
rect 5266 788 5268 792
rect 300 778 302 782
rect 2493 778 2494 782
rect 469 768 470 772
rect 692 768 694 772
rect 1122 768 1129 771
rect 1190 768 1201 771
rect 1502 768 1510 771
rect 1541 768 1542 772
rect 1788 768 1790 772
rect 2140 768 2142 772
rect 3556 768 3558 772
rect 3698 768 3705 771
rect 4262 768 4273 771
rect 4954 768 4990 771
rect 5170 768 5173 772
rect 1190 762 1193 768
rect 4270 762 4273 768
rect 154 748 161 751
rect 166 748 174 751
rect 206 751 209 761
rect 1110 758 1118 761
rect 1126 758 1137 761
rect 2230 758 2241 761
rect 2334 758 2345 761
rect 2434 758 2441 761
rect 3033 758 3038 762
rect 2238 752 2241 758
rect 3910 752 3913 761
rect 4326 758 4353 761
rect 4394 758 4398 762
rect 4498 758 4502 762
rect 4702 758 4729 761
rect 4934 758 4945 761
rect 5126 761 5129 768
rect 5118 758 5129 761
rect 5118 752 5122 754
rect 206 748 214 751
rect 254 748 270 751
rect 142 738 158 741
rect 270 738 273 748
rect 438 742 441 751
rect 454 748 465 751
rect 574 748 582 751
rect 714 748 721 751
rect 454 742 457 748
rect 334 738 348 741
rect 406 738 425 741
rect 582 738 585 748
rect 1046 748 1054 751
rect 1070 748 1094 751
rect 1302 748 1313 751
rect 1446 748 1454 751
rect 1686 748 1694 751
rect 1310 742 1313 748
rect 2078 748 2089 751
rect 2314 748 2321 751
rect 2382 748 2409 751
rect 2414 748 2422 751
rect 2494 748 2521 751
rect 2526 748 2534 751
rect 2542 748 2561 751
rect 2662 748 2681 751
rect 2686 748 2705 751
rect 2862 748 2894 751
rect 2086 742 2089 748
rect 594 738 609 741
rect 710 738 721 741
rect 726 738 738 741
rect 1078 738 1086 741
rect 1174 738 1185 741
rect 1378 738 1401 741
rect 1470 738 1478 741
rect 1602 738 1609 741
rect 1918 738 1934 741
rect 2198 738 2214 741
rect 2534 738 2545 741
rect 2558 738 2561 748
rect 3058 748 3065 751
rect 2606 738 2617 741
rect 2654 738 2665 741
rect 2998 738 3009 741
rect 3062 738 3065 748
rect 3330 748 3337 751
rect 3382 742 3385 751
rect 3426 748 3441 751
rect 3518 748 3526 751
rect 3634 748 3641 751
rect 3914 748 3921 751
rect 4366 748 4382 751
rect 4730 748 4737 751
rect 4746 748 4769 751
rect 4894 748 4921 751
rect 4926 748 4934 751
rect 5102 748 5113 751
rect 5110 742 5113 748
rect 3142 738 3150 741
rect 3322 738 3329 741
rect 3398 738 3406 741
rect 3630 738 3641 741
rect 3658 738 3673 741
rect 3678 738 3697 741
rect 3798 738 3806 741
rect 3854 738 3862 741
rect 4138 738 4145 741
rect 4482 738 4489 741
rect 4754 738 4761 741
rect 4862 738 4897 741
rect 4942 738 4950 741
rect 5086 738 5094 741
rect 5294 738 5302 741
rect 334 732 337 738
rect 150 728 161 731
rect 502 731 505 738
rect 734 736 738 738
rect 1182 732 1185 738
rect 494 728 505 731
rect 1438 731 1441 738
rect 1410 728 1425 731
rect 1430 728 1441 731
rect 1878 728 1886 731
rect 1974 731 1978 733
rect 2254 732 2257 738
rect 2662 732 2665 738
rect 2998 736 3002 738
rect 1966 728 1978 731
rect 2250 728 2257 732
rect 3350 728 3361 731
rect 3906 728 3918 731
rect 3934 728 3953 731
rect 4450 728 4462 731
rect 158 718 161 728
rect 900 718 902 722
rect 933 718 934 722
rect 2588 718 2590 722
rect 2756 718 2758 722
rect 3092 718 3094 722
rect 3950 721 3953 728
rect 3950 718 3961 721
rect 856 703 858 707
rect 862 703 865 707
rect 869 703 872 707
rect 1872 703 1874 707
rect 1878 703 1881 707
rect 1885 703 1888 707
rect 2904 703 2906 707
rect 2910 703 2913 707
rect 2917 703 2920 707
rect 3928 703 3930 707
rect 3934 703 3937 707
rect 3941 703 3944 707
rect 4952 703 4954 707
rect 4958 703 4961 707
rect 4965 703 4968 707
rect 362 688 369 691
rect 390 688 398 691
rect 628 688 630 692
rect 794 688 795 692
rect 1189 688 1190 692
rect 1690 688 1692 692
rect 1756 688 1758 692
rect 1858 688 1860 692
rect 1930 688 1932 692
rect 2108 688 2110 692
rect 2154 688 2156 692
rect 2322 688 2324 692
rect 2834 688 2835 692
rect 2938 688 2939 692
rect 3058 688 3060 692
rect 3124 688 3126 692
rect 3325 688 3326 692
rect 3450 688 3457 691
rect 4796 688 4798 692
rect 4966 688 4974 691
rect 4994 688 5015 691
rect 206 672 209 681
rect 862 678 870 681
rect 2758 678 2774 681
rect 2834 678 2849 681
rect 3638 678 3649 681
rect 4370 678 4377 681
rect 4746 678 4753 681
rect 4934 678 4942 681
rect 142 668 158 671
rect 234 668 249 671
rect 446 671 449 678
rect 3638 677 3642 678
rect 438 668 449 671
rect 462 668 478 671
rect 562 668 569 671
rect 906 668 913 671
rect 994 668 1001 671
rect 1038 668 1046 671
rect 46 658 54 661
rect 158 661 161 668
rect 158 658 177 661
rect 194 658 201 661
rect 218 658 225 661
rect 518 658 534 661
rect 554 658 577 661
rect 874 658 897 661
rect 1062 658 1089 661
rect 1782 661 1785 671
rect 1886 668 1894 671
rect 2358 668 2366 671
rect 2478 668 2489 671
rect 2522 668 2529 671
rect 2610 668 2625 671
rect 2730 668 2745 671
rect 2750 668 2758 671
rect 2486 662 2489 668
rect 1778 658 1785 661
rect 1802 658 1809 661
rect 2034 658 2041 661
rect 2350 658 2361 661
rect 2514 658 2537 661
rect 2542 658 2550 661
rect 2622 658 2625 668
rect 2914 668 2929 671
rect 2974 668 2993 671
rect 2702 658 2713 661
rect 2942 658 2961 661
rect 3006 661 3009 671
rect 3030 662 3033 671
rect 3542 668 3554 671
rect 3782 671 3785 678
rect 3782 668 3793 671
rect 4434 668 4446 671
rect 4818 668 4825 671
rect 2990 658 3009 661
rect 3394 658 3401 661
rect 3830 662 3834 664
rect 3722 658 3729 661
rect 3946 658 3961 661
rect 3978 658 3985 661
rect 4246 658 4254 661
rect 4598 658 4622 661
rect 4894 658 4910 661
rect 5030 661 5033 668
rect 5030 658 5065 661
rect 1422 652 1425 658
rect 2350 652 2353 658
rect 2710 652 2713 658
rect 190 648 201 651
rect 346 648 353 651
rect 362 648 370 651
rect 426 648 430 652
rect 546 648 550 652
rect 1417 648 1425 652
rect 2398 648 2430 651
rect 2822 651 2825 658
rect 2814 648 2825 651
rect 2942 648 2945 658
rect 3926 648 3950 651
rect 4150 648 4169 651
rect 5078 648 5089 651
rect 366 646 370 648
rect 326 638 369 641
rect 798 641 802 644
rect 2942 642 2946 644
rect 798 638 825 641
rect 981 638 982 642
rect 2509 638 2510 642
rect 4010 638 4011 642
rect 4290 638 4294 642
rect 2390 628 2393 638
rect 2886 628 2889 638
rect 4221 628 4222 632
rect 1346 618 1350 622
rect 3765 618 3766 622
rect 4189 618 4190 622
rect 344 603 346 607
rect 350 603 353 607
rect 357 603 360 607
rect 1368 603 1370 607
rect 1374 603 1377 607
rect 1381 603 1384 607
rect 2392 603 2394 607
rect 2398 603 2401 607
rect 2405 603 2408 607
rect 3416 603 3418 607
rect 3422 603 3425 607
rect 3429 603 3432 607
rect 4440 603 4442 607
rect 4446 603 4449 607
rect 4453 603 4456 607
rect 269 588 270 592
rect 413 588 414 592
rect 442 588 443 592
rect 1042 588 1043 592
rect 1130 588 1134 592
rect 1444 588 1446 592
rect 1604 588 1606 592
rect 1660 588 1662 592
rect 1730 588 1732 592
rect 2466 588 2467 592
rect 2741 588 2742 592
rect 2818 588 2819 592
rect 3372 588 3374 592
rect 174 568 185 571
rect 374 568 402 571
rect 490 568 497 571
rect 778 568 793 571
rect 1898 568 1905 571
rect 2434 568 2435 572
rect 2590 568 2606 571
rect 3236 568 3238 572
rect 3262 568 3273 571
rect 3316 568 3318 572
rect 3514 568 3516 572
rect 3734 568 3750 571
rect 3894 568 3902 571
rect 3906 568 3926 571
rect 4510 568 4521 571
rect 182 562 185 568
rect 246 558 257 561
rect 454 558 481 561
rect 770 558 777 561
rect 1054 558 1065 561
rect 1926 561 1929 568
rect 2358 561 2361 568
rect 3262 562 3265 568
rect 4518 562 4521 568
rect 1926 558 1937 561
rect 2350 558 2361 561
rect 2478 558 2505 561
rect 2689 558 2697 562
rect 3078 558 3086 561
rect 3686 558 3697 561
rect 3706 558 3718 561
rect 4238 558 4249 561
rect 4606 558 4617 561
rect 230 551 234 554
rect 230 548 238 551
rect 418 548 441 551
rect 822 548 833 551
rect 1022 548 1041 551
rect 198 541 201 548
rect 1542 548 1550 551
rect 1806 548 1838 551
rect 1866 548 1873 551
rect 2054 548 2062 551
rect 190 538 201 541
rect 422 538 430 541
rect 722 538 729 541
rect 926 538 945 541
rect 950 538 966 541
rect 1390 538 1406 541
rect 1542 538 1545 548
rect 1694 538 1713 541
rect 1806 538 1809 548
rect 2290 548 2297 551
rect 2374 551 2377 558
rect 2694 552 2697 558
rect 5174 556 5178 558
rect 2374 548 2385 551
rect 2390 548 2430 551
rect 2722 548 2729 551
rect 2946 548 2953 551
rect 2990 548 3001 551
rect 3142 548 3166 551
rect 3542 548 3553 551
rect 3778 548 3785 551
rect 4014 548 4022 551
rect 2322 538 2329 541
rect 2418 538 2425 541
rect 2774 538 2793 541
rect 2902 538 2953 541
rect 2962 538 2969 541
rect 2998 538 3001 548
rect 3542 542 3545 548
rect 3190 538 3198 541
rect 3270 538 3289 541
rect 3574 538 3582 541
rect 3598 538 3606 541
rect 3622 538 3638 541
rect 3930 538 3945 541
rect 4030 541 4033 548
rect 4134 542 4137 551
rect 4274 548 4281 551
rect 4522 548 4529 551
rect 3974 538 3993 541
rect 4022 538 4033 541
rect 4046 538 4065 541
rect 4214 538 4241 541
rect 4278 538 4289 541
rect 4574 541 4577 551
rect 4582 548 4593 551
rect 4634 548 4665 551
rect 4706 548 4713 551
rect 4886 548 4894 551
rect 4566 538 4577 541
rect 4590 542 4593 548
rect 4662 538 4665 548
rect 5046 546 5050 548
rect 4738 538 4742 541
rect 4870 538 4878 541
rect 4918 538 4937 541
rect 910 532 913 538
rect 754 528 758 532
rect 886 528 894 531
rect 910 528 918 532
rect 2326 528 2329 538
rect 3078 532 3081 538
rect 3830 532 3833 538
rect 4046 532 4049 538
rect 2754 528 2761 531
rect 2910 528 2926 531
rect 3074 528 3081 532
rect 3830 528 3838 532
rect 4178 528 4188 531
rect 4214 528 4217 538
rect 4278 532 4281 538
rect 4226 528 4233 531
rect 4806 528 4814 531
rect 4934 531 4937 538
rect 4926 528 4953 531
rect 1292 518 1294 522
rect 1362 518 1364 522
rect 1524 518 1526 522
rect 1698 518 1699 522
rect 2268 518 2270 522
rect 2874 518 2887 521
rect 3458 518 3460 522
rect 3722 518 3729 521
rect 4444 518 4446 522
rect 4550 518 4558 521
rect 4854 518 4862 521
rect 856 503 858 507
rect 862 503 865 507
rect 869 503 872 507
rect 1872 503 1874 507
rect 1878 503 1881 507
rect 1885 503 1888 507
rect 2904 503 2906 507
rect 2910 503 2913 507
rect 2917 503 2920 507
rect 3928 503 3930 507
rect 3934 503 3937 507
rect 3941 503 3944 507
rect 4952 503 4954 507
rect 4958 503 4961 507
rect 4965 503 4968 507
rect 108 488 110 492
rect 281 488 294 491
rect 622 488 630 491
rect 700 488 702 492
rect 1322 488 1324 492
rect 1404 488 1406 492
rect 1772 488 1774 492
rect 1874 488 1875 492
rect 2100 488 2102 492
rect 2882 488 2889 491
rect 3970 488 3977 491
rect 250 478 257 481
rect 874 478 881 481
rect 1206 472 1209 481
rect 1518 478 1529 481
rect 2750 478 2758 481
rect 3574 478 3582 482
rect 4518 478 4526 482
rect 4790 478 4798 481
rect 4812 478 4841 481
rect 5174 478 5186 481
rect 1518 477 1522 478
rect 126 468 134 471
rect 230 468 265 471
rect 454 468 462 471
rect 650 468 657 471
rect 862 468 889 471
rect 1214 468 1225 471
rect 1238 468 1257 471
rect 1266 468 1281 471
rect 1294 468 1305 471
rect 1534 468 1545 471
rect 1562 468 1577 471
rect 1790 468 1801 471
rect 2126 471 2130 474
rect 2118 468 2130 471
rect 2165 468 2166 472
rect 2342 468 2350 471
rect 2634 468 2641 471
rect 2742 468 2750 471
rect 3054 468 3066 471
rect 3150 471 3154 474
rect 3574 472 3577 478
rect 4518 472 4521 478
rect 5182 477 5186 478
rect 3150 468 3161 471
rect 3494 468 3502 471
rect 3550 468 3558 471
rect 3726 468 3737 471
rect 3878 468 3886 471
rect 3926 468 3934 471
rect 4194 468 4206 471
rect 4350 468 4358 471
rect 4366 468 4382 471
rect 4430 468 4438 471
rect 4450 468 4465 471
rect 4786 468 4793 471
rect 5098 468 5105 471
rect 862 462 865 468
rect 46 458 54 461
rect 750 458 774 461
rect 942 461 945 468
rect 934 458 945 461
rect 1222 462 1225 468
rect 1542 462 1545 468
rect 1814 458 1833 461
rect 1890 458 1913 461
rect 1998 458 2006 461
rect 2414 458 2422 461
rect 2774 461 2777 468
rect 3726 462 3729 468
rect 2766 458 2777 461
rect 3538 458 3545 461
rect 3678 458 3686 461
rect 3702 458 3713 461
rect 3870 458 3878 461
rect 3882 458 3897 461
rect 3902 458 3910 461
rect 4018 458 4025 461
rect 4038 458 4054 461
rect 4082 458 4089 461
rect 4098 458 4113 461
rect 4214 458 4222 461
rect 4782 461 4785 468
rect 4758 458 4785 461
rect 4794 458 4801 461
rect 5090 458 5113 461
rect 5118 458 5138 461
rect 5174 461 5177 468
rect 5174 458 5186 461
rect 1982 456 1986 458
rect 2870 456 2874 458
rect 377 448 382 452
rect 634 448 641 451
rect 886 448 897 451
rect 1878 448 1886 451
rect 1898 448 1905 451
rect 2034 448 2039 452
rect 3594 448 3601 451
rect 3686 448 3694 451
rect 4022 448 4025 458
rect 5134 456 5138 458
rect 5182 457 5186 458
rect 4510 448 4518 451
rect 5166 448 5174 451
rect 626 438 638 441
rect 690 438 697 441
rect 1686 438 1702 441
rect 2146 438 2149 442
rect 2986 438 2989 442
rect 3131 438 3134 442
rect 3514 438 3515 442
rect 3869 438 3870 442
rect 4757 438 4758 442
rect 4150 428 4153 438
rect 2250 418 2254 422
rect 3266 418 3270 422
rect 3645 418 3646 422
rect 4970 418 4985 421
rect 344 403 346 407
rect 350 403 353 407
rect 357 403 360 407
rect 1368 403 1370 407
rect 1374 403 1377 407
rect 1381 403 1384 407
rect 2392 403 2394 407
rect 2398 403 2401 407
rect 2405 403 2408 407
rect 3416 403 3418 407
rect 3422 403 3425 407
rect 3429 403 3432 407
rect 4440 403 4442 407
rect 4446 403 4449 407
rect 4453 403 4456 407
rect 172 388 174 392
rect 653 388 654 392
rect 685 388 686 392
rect 954 388 956 392
rect 1020 388 1022 392
rect 1172 388 1174 392
rect 1218 388 1220 392
rect 1898 388 1899 392
rect 2546 388 2547 392
rect 2578 388 2579 392
rect 5154 388 5155 392
rect 5294 388 5310 391
rect 2442 378 2444 382
rect 2750 372 2753 381
rect 340 368 342 372
rect 402 368 404 372
rect 1558 368 1586 371
rect 1741 368 1742 372
rect 1850 368 1851 372
rect 1942 368 1966 371
rect 2090 368 2091 372
rect 2174 368 2182 371
rect 2274 368 2277 372
rect 2682 368 2689 371
rect 2834 368 2849 371
rect 3650 368 3657 371
rect 4682 368 4683 372
rect 566 361 569 368
rect 1582 366 1586 368
rect 558 358 569 361
rect 614 358 641 361
rect 1286 358 1297 361
rect 1942 358 1945 368
rect 2590 358 2601 361
rect 3434 358 3441 361
rect 3634 358 3641 361
rect 3838 358 3846 361
rect 3918 358 3926 361
rect 4086 361 4089 368
rect 4086 358 4097 361
rect 5062 358 5089 361
rect 5166 358 5178 361
rect 190 348 209 351
rect 190 342 193 348
rect 1246 348 1265 351
rect 1298 348 1305 351
rect 1310 348 1329 351
rect 1406 348 1425 351
rect 1534 348 1542 351
rect 1630 348 1641 351
rect 1662 348 1673 351
rect 1682 348 1689 351
rect 1742 348 1750 351
rect 2182 351 2185 358
rect 5174 356 5178 358
rect 2114 348 2137 351
rect 2182 348 2193 351
rect 2306 348 2313 351
rect 2370 348 2377 351
rect 2410 348 2425 351
rect 2502 348 2513 351
rect 2526 348 2534 351
rect 2622 348 2633 351
rect 118 338 129 341
rect 1246 338 1249 348
rect 1346 338 1353 341
rect 1434 338 1441 341
rect 1666 338 1673 341
rect 1774 338 1801 341
rect 1822 338 1830 341
rect 2122 338 2129 341
rect 2422 338 2425 348
rect 2510 342 2513 348
rect 2630 342 2633 348
rect 3494 348 3502 351
rect 3874 348 3881 351
rect 4026 348 4049 351
rect 4502 348 4510 351
rect 2966 338 2978 341
rect 3462 338 3473 341
rect 3574 338 3593 341
rect 3598 338 3614 341
rect 3818 338 3820 342
rect 3886 338 3900 341
rect 4158 338 4166 341
rect 4542 341 4545 348
rect 4662 342 4665 351
rect 4978 348 4985 351
rect 5018 348 5025 351
rect 5130 348 5153 351
rect 5206 348 5214 351
rect 4542 338 4553 341
rect 4574 338 4593 341
rect 4630 338 4649 341
rect 4690 338 4705 341
rect 5274 338 5281 341
rect 118 336 122 338
rect 582 332 585 338
rect 1582 332 1585 338
rect 578 328 585 332
rect 806 328 814 331
rect 1386 328 1393 331
rect 1582 328 1590 332
rect 2182 328 2190 331
rect 2230 331 2233 338
rect 3462 332 3465 338
rect 2230 328 2241 331
rect 3502 328 3513 331
rect 3518 328 3526 331
rect 3998 331 4001 338
rect 5174 336 5178 338
rect 3998 328 4009 331
rect 4662 328 4670 331
rect 770 318 771 322
rect 2874 318 2881 321
rect 3274 318 3276 322
rect 3362 318 3364 322
rect 3650 318 3657 321
rect 3690 318 3692 322
rect 3746 318 3748 322
rect 4186 318 4188 322
rect 4298 318 4300 322
rect 856 303 858 307
rect 862 303 865 307
rect 869 303 872 307
rect 1872 303 1874 307
rect 1878 303 1881 307
rect 1885 303 1888 307
rect 2904 303 2906 307
rect 2910 303 2913 307
rect 2917 303 2920 307
rect 3928 303 3930 307
rect 3934 303 3937 307
rect 3941 303 3944 307
rect 4952 303 4954 307
rect 4958 303 4961 307
rect 4965 303 4968 307
rect 450 288 452 292
rect 602 288 604 292
rect 882 288 884 292
rect 1106 288 1108 292
rect 1172 288 1174 292
rect 1469 288 1470 292
rect 1516 288 1518 292
rect 2406 288 2422 291
rect 2674 288 2676 292
rect 2733 288 2734 292
rect 3546 288 3548 292
rect 4138 288 4145 291
rect 4210 288 4212 292
rect 4346 288 4348 292
rect 5034 288 5041 291
rect 5286 288 5294 291
rect 230 278 238 281
rect 1370 278 1382 281
rect 1678 272 1681 281
rect 2974 272 2977 281
rect 4398 274 4402 278
rect 5166 272 5169 281
rect 174 268 204 271
rect 334 268 358 271
rect 426 268 433 271
rect 810 268 817 271
rect 234 258 257 261
rect 274 258 281 261
rect 298 258 305 261
rect 518 258 526 261
rect 798 258 822 261
rect 954 258 961 261
rect 974 261 977 271
rect 1006 268 1014 271
rect 1602 268 1617 271
rect 1686 262 1689 271
rect 1746 268 1753 271
rect 1962 268 1969 271
rect 2470 268 2486 271
rect 2718 268 2726 271
rect 3154 268 3161 271
rect 3286 268 3294 271
rect 3634 268 3641 271
rect 3742 268 3753 271
rect 4186 268 4193 271
rect 4238 268 4246 271
rect 4262 268 4281 271
rect 4286 268 4302 271
rect 4318 268 4329 271
rect 4654 268 4665 271
rect 4798 268 4809 271
rect 4914 268 4921 271
rect 5046 268 5057 271
rect 974 258 985 261
rect 1070 258 1086 261
rect 1230 258 1238 261
rect 1342 258 1369 261
rect 1770 258 1793 261
rect 1798 258 1809 261
rect 1814 258 1822 261
rect 1926 258 1950 261
rect 2274 258 2281 261
rect 2526 261 2529 268
rect 2526 258 2561 261
rect 2830 261 2833 268
rect 3750 262 3753 268
rect 4662 262 4665 268
rect 5046 262 5049 268
rect 2810 258 2825 261
rect 2830 258 2841 261
rect 3034 258 3057 261
rect 3098 258 3113 261
rect 3118 258 3129 261
rect 3162 258 3185 261
rect 3266 258 3273 261
rect 3278 258 3305 261
rect 3322 258 3329 261
rect 3590 258 3609 261
rect 3614 258 3633 261
rect 1806 252 1809 258
rect 3118 252 3121 258
rect 354 248 369 251
rect 758 248 785 251
rect 794 248 798 252
rect 1062 248 1073 251
rect 1198 248 1217 251
rect 1374 248 1398 251
rect 1662 248 1689 251
rect 2574 248 2585 251
rect 2958 248 2985 251
rect 3254 248 3265 251
rect 3330 248 3334 252
rect 3630 248 3633 258
rect 4058 258 4065 261
rect 4106 258 4113 261
rect 4318 258 4326 261
rect 4434 258 4441 261
rect 4730 258 4745 261
rect 4810 258 4817 261
rect 4822 258 4830 261
rect 4846 258 4857 261
rect 5094 258 5102 261
rect 5154 258 5177 261
rect 3646 251 3649 258
rect 3646 248 3657 251
rect 4126 248 4134 251
rect 4926 248 4937 251
rect 5070 248 5078 251
rect 4926 242 4929 248
rect 94 238 118 241
rect 362 238 382 241
rect 658 238 673 241
rect 1229 238 1230 242
rect 2291 238 2294 242
rect 4402 238 4405 242
rect 5046 241 5050 244
rect 5034 238 5050 241
rect 165 218 166 222
rect 826 218 827 222
rect 2090 218 2092 222
rect 2628 218 2630 222
rect 2997 218 2998 222
rect 3029 218 3030 222
rect 3277 218 3278 222
rect 3690 218 3692 222
rect 4770 218 4771 222
rect 344 203 346 207
rect 350 203 353 207
rect 357 203 360 207
rect 1368 203 1370 207
rect 1374 203 1377 207
rect 1381 203 1384 207
rect 2392 203 2394 207
rect 2398 203 2401 207
rect 2405 203 2408 207
rect 3416 203 3418 207
rect 3422 203 3425 207
rect 3429 203 3432 207
rect 4440 203 4442 207
rect 4446 203 4449 207
rect 4453 203 4456 207
rect 149 188 150 192
rect 274 188 276 192
rect 730 188 732 192
rect 1477 188 1478 192
rect 1773 188 1774 192
rect 1834 188 1835 192
rect 1978 188 1980 192
rect 2082 188 2084 192
rect 2354 188 2356 192
rect 2618 188 2620 192
rect 4506 188 4508 192
rect 1546 168 1562 171
rect 1590 168 1598 171
rect 1874 168 1897 171
rect 2562 168 2564 172
rect 2718 168 2742 171
rect 3194 168 3196 172
rect 3326 168 3337 171
rect 3746 168 3753 171
rect 3830 168 3841 171
rect 4762 168 4769 171
rect 5278 168 5294 171
rect 1558 166 1562 168
rect 3326 162 3329 168
rect 3830 162 3833 168
rect 126 158 137 161
rect 110 151 114 154
rect 110 148 118 151
rect 150 148 169 151
rect 326 151 329 161
rect 338 158 353 161
rect 1734 158 1761 161
rect 186 148 193 151
rect 302 148 321 151
rect 326 148 361 151
rect 370 148 382 151
rect 666 148 689 151
rect 694 148 702 151
rect 758 148 769 151
rect 894 148 902 151
rect 950 148 958 151
rect 974 148 985 151
rect 1054 151 1058 154
rect 1054 148 1065 151
rect 1190 151 1193 158
rect 1190 148 1201 151
rect 166 142 169 148
rect 170 138 185 141
rect 302 138 305 148
rect 318 138 334 141
rect 390 138 417 141
rect 530 138 540 141
rect 674 138 681 141
rect 758 138 761 148
rect 858 138 881 141
rect 930 138 937 141
rect 1014 138 1022 141
rect 1062 138 1065 148
rect 1806 148 1833 151
rect 2402 148 2409 151
rect 2758 151 2761 161
rect 2810 158 2814 162
rect 2874 158 2881 161
rect 3698 158 3702 162
rect 4810 158 4814 162
rect 4822 158 4833 161
rect 4954 158 4961 161
rect 5126 158 5137 161
rect 2758 148 2777 151
rect 2910 148 2926 151
rect 3014 148 3022 151
rect 3038 148 3073 151
rect 3166 148 3174 151
rect 3258 148 3265 151
rect 3270 148 3289 151
rect 3294 148 3302 151
rect 3306 148 3321 151
rect 3414 148 3438 151
rect 3510 148 3521 151
rect 3670 148 3694 151
rect 3714 148 3729 151
rect 3890 148 3897 151
rect 1178 138 1185 141
rect 1430 138 1438 141
rect 1486 138 1505 141
rect 2166 138 2174 141
rect 2190 141 2193 148
rect 2190 138 2201 141
rect 2678 141 2681 148
rect 3070 142 3073 148
rect 3166 146 3170 148
rect 2646 138 2665 141
rect 2670 138 2681 141
rect 2716 138 2718 142
rect 2862 138 2873 141
rect 2910 138 2934 141
rect 2938 138 2945 141
rect 3018 138 3025 141
rect 3114 138 3129 141
rect 3302 138 3310 141
rect 3530 138 3545 141
rect 3654 138 3657 148
rect 3994 148 4009 151
rect 4438 148 4473 151
rect 3678 138 3686 141
rect 622 128 630 131
rect 994 128 1001 131
rect 1486 128 1489 138
rect 1558 132 1561 138
rect 1558 128 1566 132
rect 1742 128 1745 138
rect 2042 128 2046 132
rect 2166 128 2169 138
rect 2178 128 2182 132
rect 2214 131 2218 133
rect 2870 132 2873 138
rect 2206 128 2218 131
rect 2910 128 2913 138
rect 2922 128 2937 131
rect 3230 131 3233 138
rect 3982 132 3985 142
rect 4470 141 4473 148
rect 4838 151 4841 158
rect 4802 148 4809 151
rect 4838 148 4849 151
rect 5142 151 5145 158
rect 5142 148 5161 151
rect 4470 138 4489 141
rect 4646 138 4649 148
rect 5074 138 5076 142
rect 4918 132 4921 138
rect 5174 132 5178 133
rect 3230 128 3241 131
rect 4694 128 4702 131
rect 4750 128 4758 131
rect 4918 128 4926 132
rect 237 118 238 122
rect 460 118 462 122
rect 820 118 822 122
rect 2450 118 2452 122
rect 2506 118 2508 122
rect 2661 118 2662 122
rect 2973 118 2974 122
rect 3814 118 3822 121
rect 4292 118 4294 122
rect 4378 118 4380 122
rect 4562 118 4564 122
rect 4618 118 4620 122
rect 856 103 858 107
rect 862 103 865 107
rect 869 103 872 107
rect 1872 103 1874 107
rect 1878 103 1881 107
rect 1885 103 1888 107
rect 2904 103 2906 107
rect 2910 103 2913 107
rect 2917 103 2920 107
rect 3928 103 3930 107
rect 3934 103 3937 107
rect 3941 103 3944 107
rect 4952 103 4954 107
rect 4958 103 4961 107
rect 4965 103 4968 107
rect 562 88 563 92
rect 850 88 852 92
rect 1090 88 1091 92
rect 1340 88 1342 92
rect 1402 88 1404 92
rect 1574 88 1582 91
rect 1606 88 1614 91
rect 1834 88 1835 92
rect 1858 88 1865 91
rect 2338 88 2340 92
rect 2466 88 2468 92
rect 2618 88 2620 92
rect 2700 88 2702 92
rect 2749 88 2750 92
rect 3034 88 3036 92
rect 3386 88 3388 92
rect 3934 88 3942 91
rect 4610 88 4612 92
rect 4874 88 4876 92
rect 442 78 449 81
rect 666 78 673 81
rect 178 68 185 71
rect 306 68 313 71
rect 430 68 438 71
rect 502 68 518 71
rect 570 68 577 71
rect 822 68 833 71
rect 22 58 30 61
rect 186 58 209 61
rect 266 58 281 61
rect 342 58 390 61
rect 470 61 473 68
rect 462 58 473 61
rect 626 58 633 61
rect 750 58 777 61
rect 878 61 881 71
rect 910 68 921 71
rect 1030 71 1033 81
rect 2118 78 2130 81
rect 2666 78 2673 82
rect 2126 77 2130 78
rect 1010 68 1033 71
rect 1140 68 1142 72
rect 1226 68 1233 71
rect 1250 68 1257 71
rect 1522 68 1545 71
rect 1682 68 1697 71
rect 2310 71 2314 74
rect 2670 72 2673 78
rect 2106 68 2113 71
rect 2214 68 2226 71
rect 2310 68 2321 71
rect 2846 71 2849 78
rect 2846 68 2889 71
rect 2974 68 2985 71
rect 3062 68 3073 71
rect 3098 68 3105 71
rect 3166 68 3177 71
rect 3182 68 3201 71
rect 3356 68 3358 72
rect 3462 68 3473 71
rect 878 58 913 61
rect 934 58 961 61
rect 1158 58 1166 61
rect 1174 58 1193 61
rect 1198 58 1206 61
rect 1238 58 1270 61
rect 1630 58 1641 61
rect 1754 58 1777 61
rect 3174 62 3177 68
rect 2922 58 2953 61
rect 3090 58 3113 61
rect 3226 58 3249 61
rect 3518 61 3521 71
rect 3534 68 3545 71
rect 3622 68 3630 71
rect 3730 68 3732 72
rect 3910 71 3913 78
rect 4270 72 4273 81
rect 5166 78 5178 81
rect 5174 77 5178 78
rect 3850 68 3865 71
rect 3902 68 3913 71
rect 4070 68 4082 71
rect 4278 68 4289 71
rect 4358 68 4369 71
rect 4734 71 4738 74
rect 4734 68 4745 71
rect 3434 58 3449 61
rect 3518 58 3537 61
rect 3558 58 3585 61
rect 3638 58 3646 61
rect 3670 58 3689 61
rect 3694 58 3702 61
rect 4026 58 4041 61
rect 4286 62 4289 68
rect 4110 58 4118 61
rect 4206 58 4214 61
rect 4294 58 4302 61
rect 4538 58 4553 61
rect 4678 58 4686 61
rect 4854 61 4857 71
rect 5206 68 5209 78
rect 4762 58 4769 61
rect 4830 58 4857 61
rect 4978 58 4985 61
rect 5218 58 5233 61
rect 1158 56 1162 58
rect 1630 52 1633 58
rect 2678 56 2682 58
rect 1206 48 1217 51
rect 1281 48 1286 52
rect 1694 48 1705 51
rect 2758 51 2761 58
rect 2758 48 2769 51
rect 2806 48 2817 51
rect 3330 48 3337 51
rect 3686 48 3689 58
rect 3822 51 3825 58
rect 3822 48 3833 51
rect 5038 51 5041 58
rect 5038 48 5049 51
rect 5122 48 5124 52
rect 282 38 283 42
rect 702 41 706 44
rect 702 38 729 41
rect 962 38 963 42
rect 2410 38 2412 42
rect 3490 38 3492 42
rect 3702 41 3705 48
rect 3702 38 3713 41
rect 4386 38 4388 42
rect 344 3 346 7
rect 350 3 353 7
rect 357 3 360 7
rect 1368 3 1370 7
rect 1374 3 1377 7
rect 1381 3 1384 7
rect 2392 3 2394 7
rect 2398 3 2401 7
rect 2405 3 2408 7
rect 3416 3 3418 7
rect 3422 3 3425 7
rect 3429 3 3432 7
rect 4440 3 4442 7
rect 4446 3 4449 7
rect 4453 3 4456 7
<< m2contact >>
rect 858 3703 862 3707
rect 865 3703 869 3707
rect 1874 3703 1878 3707
rect 1881 3703 1885 3707
rect 2906 3703 2910 3707
rect 2913 3703 2917 3707
rect 3930 3703 3934 3707
rect 3937 3703 3941 3707
rect 4954 3703 4958 3707
rect 4961 3703 4965 3707
rect 1446 3698 1450 3702
rect 1806 3698 1810 3702
rect 494 3688 498 3692
rect 694 3688 698 3692
rect 1110 3688 1114 3692
rect 1198 3688 1202 3692
rect 1574 3688 1578 3692
rect 1734 3688 1738 3692
rect 1782 3688 1786 3692
rect 1966 3688 1970 3692
rect 1982 3688 1986 3692
rect 2270 3688 2274 3692
rect 2750 3688 2754 3692
rect 2942 3688 2946 3692
rect 2974 3688 2978 3692
rect 3110 3688 3114 3692
rect 3158 3688 3162 3692
rect 3302 3688 3306 3692
rect 3318 3688 3322 3692
rect 3382 3688 3386 3692
rect 3390 3688 3394 3692
rect 3622 3688 3626 3692
rect 3662 3688 3666 3692
rect 3686 3688 3690 3692
rect 3854 3688 3858 3692
rect 3982 3688 3986 3692
rect 4102 3688 4106 3692
rect 4302 3688 4306 3692
rect 4438 3688 4442 3692
rect 4590 3688 4594 3692
rect 4710 3688 4714 3692
rect 4774 3688 4778 3692
rect 4894 3688 4898 3692
rect 5158 3688 5162 3692
rect 5182 3688 5186 3692
rect 14 3679 18 3683
rect 38 3679 42 3683
rect 62 3679 66 3683
rect 86 3679 90 3683
rect 110 3679 114 3683
rect 134 3679 138 3683
rect 158 3679 162 3683
rect 206 3679 210 3683
rect 230 3679 234 3683
rect 294 3678 298 3682
rect 318 3678 322 3682
rect 286 3668 290 3672
rect 366 3668 370 3672
rect 406 3678 410 3682
rect 534 3678 538 3682
rect 630 3678 634 3682
rect 742 3678 746 3682
rect 406 3668 410 3672
rect 414 3668 418 3672
rect 454 3668 458 3672
rect 462 3668 466 3672
rect 566 3668 570 3672
rect 598 3668 602 3672
rect 614 3668 618 3672
rect 622 3668 626 3672
rect 670 3668 674 3672
rect 702 3668 706 3672
rect 734 3668 738 3672
rect 838 3678 842 3682
rect 910 3678 914 3682
rect 934 3678 938 3682
rect 990 3678 994 3682
rect 1214 3678 1218 3682
rect 1222 3678 1226 3682
rect 1270 3678 1274 3682
rect 1318 3678 1322 3682
rect 1446 3678 1450 3682
rect 1606 3678 1610 3682
rect 1630 3678 1634 3682
rect 1686 3678 1690 3682
rect 1806 3678 1810 3682
rect 1998 3678 2002 3682
rect 2038 3679 2042 3683
rect 2054 3678 2058 3682
rect 2078 3679 2082 3683
rect 2094 3678 2098 3682
rect 2214 3679 2218 3683
rect 2230 3678 2234 3682
rect 2310 3678 2314 3682
rect 2318 3678 2322 3682
rect 2358 3678 2362 3682
rect 2446 3678 2450 3682
rect 2494 3678 2498 3682
rect 2550 3678 2554 3682
rect 2558 3678 2562 3682
rect 2598 3679 2602 3683
rect 2622 3679 2626 3683
rect 2638 3678 2642 3682
rect 2918 3678 2922 3682
rect 3118 3678 3122 3682
rect 3326 3678 3330 3682
rect 3846 3678 3850 3682
rect 4086 3678 4090 3682
rect 4182 3678 4186 3682
rect 4310 3678 4314 3682
rect 4414 3678 4418 3682
rect 4718 3678 4722 3682
rect 4886 3678 4890 3682
rect 5006 3678 5010 3682
rect 5038 3678 5042 3682
rect 5198 3679 5202 3683
rect 774 3668 778 3672
rect 790 3668 794 3672
rect 846 3668 850 3672
rect 950 3668 954 3672
rect 966 3668 970 3672
rect 998 3668 1002 3672
rect 1046 3668 1050 3672
rect 1078 3668 1082 3672
rect 1126 3668 1130 3672
rect 1158 3668 1162 3672
rect 1206 3668 1210 3672
rect 1230 3668 1234 3672
rect 1422 3668 1426 3672
rect 1454 3668 1458 3672
rect 6 3658 10 3662
rect 30 3658 34 3662
rect 54 3658 58 3662
rect 78 3658 82 3662
rect 102 3658 106 3662
rect 142 3658 146 3662
rect 166 3658 170 3662
rect 198 3658 202 3662
rect 222 3658 226 3662
rect 262 3658 266 3662
rect 342 3658 346 3662
rect 374 3658 378 3662
rect 398 3658 402 3662
rect 422 3658 426 3662
rect 446 3658 450 3662
rect 518 3658 522 3662
rect 558 3658 562 3662
rect 590 3658 594 3662
rect 606 3658 610 3662
rect 646 3658 650 3662
rect 1566 3668 1570 3672
rect 1598 3668 1602 3672
rect 1606 3668 1610 3672
rect 1638 3668 1642 3672
rect 1670 3668 1674 3672
rect 1694 3668 1698 3672
rect 726 3658 730 3662
rect 806 3658 810 3662
rect 886 3658 890 3662
rect 942 3658 946 3662
rect 958 3658 962 3662
rect 974 3658 978 3662
rect 990 3658 994 3662
rect 1054 3658 1058 3662
rect 1158 3658 1162 3662
rect 1238 3658 1242 3662
rect 1294 3658 1298 3662
rect 1310 3658 1314 3662
rect 1342 3658 1346 3662
rect 1430 3658 1434 3662
rect 1446 3658 1450 3662
rect 1478 3658 1482 3662
rect 1502 3658 1506 3662
rect 1526 3658 1530 3662
rect 1574 3658 1578 3662
rect 1590 3658 1594 3662
rect 1662 3658 1666 3662
rect 1726 3658 1730 3662
rect 1750 3668 1754 3672
rect 1798 3668 1802 3672
rect 1862 3668 1866 3672
rect 1878 3668 1882 3672
rect 1902 3668 1906 3672
rect 1950 3668 1954 3672
rect 1958 3668 1962 3672
rect 2198 3668 2202 3672
rect 2246 3668 2250 3672
rect 2278 3668 2282 3672
rect 2430 3668 2434 3672
rect 2446 3668 2450 3672
rect 2542 3668 2546 3672
rect 2694 3668 2698 3672
rect 2742 3668 2746 3672
rect 2854 3668 2858 3672
rect 2910 3668 2914 3672
rect 3078 3668 3082 3672
rect 3110 3668 3114 3672
rect 3222 3668 3226 3672
rect 3318 3668 3322 3672
rect 3726 3668 3730 3672
rect 3734 3668 3738 3672
rect 3822 3668 3826 3672
rect 3854 3668 3858 3672
rect 3950 3668 3954 3672
rect 4070 3668 4074 3672
rect 4102 3668 4106 3672
rect 4174 3668 4178 3672
rect 4190 3668 4194 3672
rect 4246 3668 4250 3672
rect 4326 3668 4330 3672
rect 4334 3668 4338 3672
rect 4350 3668 4354 3672
rect 4366 3668 4370 3672
rect 4446 3668 4450 3672
rect 4510 3668 4514 3672
rect 4566 3668 4570 3672
rect 4678 3668 4682 3672
rect 4710 3668 4714 3672
rect 4894 3668 4898 3672
rect 4982 3668 4986 3672
rect 4998 3668 5002 3672
rect 5078 3668 5082 3672
rect 1750 3658 1754 3662
rect 1822 3658 1826 3662
rect 1838 3658 1842 3662
rect 1910 3658 1914 3662
rect 1950 3658 1954 3662
rect 1966 3658 1970 3662
rect 1982 3658 1986 3662
rect 2006 3658 2010 3662
rect 2046 3658 2050 3662
rect 2070 3658 2074 3662
rect 2094 3658 2098 3662
rect 2126 3658 2130 3662
rect 2150 3658 2154 3662
rect 2174 3658 2178 3662
rect 2182 3658 2186 3662
rect 2190 3658 2194 3662
rect 2206 3658 2210 3662
rect 2254 3658 2258 3662
rect 2286 3658 2290 3662
rect 2342 3658 2346 3662
rect 2390 3658 2394 3662
rect 2422 3658 2426 3662
rect 2462 3658 2466 3662
rect 2518 3658 2522 3662
rect 2534 3658 2538 3662
rect 2590 3658 2594 3662
rect 2614 3658 2618 3662
rect 2638 3658 2642 3662
rect 2654 3658 2658 3662
rect 2678 3658 2682 3662
rect 2838 3659 2842 3663
rect 2902 3658 2906 3662
rect 2966 3658 2970 3662
rect 2990 3658 2994 3662
rect 3062 3659 3066 3663
rect 3118 3658 3122 3662
rect 3174 3658 3178 3662
rect 3214 3658 3218 3662
rect 3326 3658 3330 3662
rect 3366 3658 3370 3662
rect 3494 3659 3498 3663
rect 3558 3658 3562 3662
rect 3582 3658 3586 3662
rect 3638 3658 3642 3662
rect 3646 3658 3650 3662
rect 3670 3658 3674 3662
rect 3694 3658 3698 3662
rect 3702 3658 3706 3662
rect 3806 3659 3810 3663
rect 3862 3658 3866 3662
rect 3902 3658 3906 3662
rect 3910 3658 3914 3662
rect 3966 3658 3970 3662
rect 4054 3659 4058 3663
rect 4110 3658 4114 3662
rect 4182 3658 4186 3662
rect 4238 3659 4242 3663
rect 4358 3658 4362 3662
rect 4374 3658 4378 3662
rect 4390 3658 4394 3662
rect 4398 3658 4402 3662
rect 4422 3658 4426 3662
rect 4454 3658 4458 3662
rect 4494 3658 4498 3662
rect 4502 3658 4506 3662
rect 4526 3658 4530 3662
rect 4534 3658 4538 3662
rect 4574 3658 4578 3662
rect 4662 3659 4666 3663
rect 4718 3658 4722 3662
rect 4758 3658 4762 3662
rect 4814 3658 4818 3662
rect 4846 3659 4850 3663
rect 4902 3658 4906 3662
rect 4990 3658 4994 3662
rect 5022 3658 5026 3662
rect 5030 3658 5034 3662
rect 5062 3658 5066 3662
rect 5094 3659 5098 3663
rect 5190 3658 5194 3662
rect 5246 3658 5250 3662
rect 5278 3659 5282 3663
rect 270 3648 274 3652
rect 310 3648 314 3652
rect 350 3648 354 3652
rect 430 3648 434 3652
rect 542 3648 546 3652
rect 574 3648 578 3652
rect 638 3648 642 3652
rect 670 3648 674 3652
rect 766 3648 770 3652
rect 790 3648 794 3652
rect 798 3648 802 3652
rect 822 3648 826 3652
rect 830 3648 834 3652
rect 942 3648 946 3652
rect 1270 3648 1274 3652
rect 1358 3648 1362 3652
rect 1406 3648 1410 3652
rect 1438 3648 1442 3652
rect 1478 3648 1482 3652
rect 1510 3648 1514 3652
rect 1526 3648 1530 3652
rect 1630 3648 1634 3652
rect 1654 3648 1658 3652
rect 1830 3648 1834 3652
rect 1862 3648 1866 3652
rect 1934 3648 1938 3652
rect 1982 3648 1986 3652
rect 2134 3648 2138 3652
rect 2142 3648 2146 3652
rect 2230 3648 2234 3652
rect 2270 3648 2274 3652
rect 2302 3648 2306 3652
rect 2318 3648 2322 3652
rect 2366 3648 2370 3652
rect 2398 3648 2402 3652
rect 2454 3648 2458 3652
rect 2526 3648 2530 3652
rect 2662 3648 2666 3652
rect 2870 3648 2874 3652
rect 254 3638 258 3642
rect 334 3638 338 3642
rect 366 3638 370 3642
rect 654 3638 658 3642
rect 814 3638 818 3642
rect 878 3638 882 3642
rect 1286 3638 1290 3642
rect 1334 3638 1338 3642
rect 1494 3638 1498 3642
rect 1550 3638 1554 3642
rect 1838 3638 1842 3642
rect 1846 3638 1850 3642
rect 2062 3638 2066 3642
rect 2118 3638 2122 3642
rect 2150 3638 2154 3642
rect 2158 3638 2162 3642
rect 2334 3638 2338 3642
rect 2382 3638 2386 3642
rect 2470 3638 2474 3642
rect 2494 3638 2498 3642
rect 2510 3638 2514 3642
rect 3758 3638 3762 3642
rect 3990 3638 3994 3642
rect 4006 3638 4010 3642
rect 4598 3638 4602 3642
rect 5142 3638 5146 3642
rect 2342 3628 2346 3632
rect 2478 3628 2482 3632
rect 2774 3628 2778 3632
rect 262 3618 266 3622
rect 326 3618 330 3622
rect 446 3618 450 3622
rect 558 3618 562 3622
rect 646 3618 650 3622
rect 854 3618 858 3622
rect 1030 3618 1034 3622
rect 1190 3618 1194 3622
rect 1238 3618 1242 3622
rect 1294 3618 1298 3622
rect 1342 3618 1346 3622
rect 1502 3618 1506 3622
rect 1558 3618 1562 3622
rect 1646 3618 1650 3622
rect 1686 3618 1690 3622
rect 1838 3618 1842 3622
rect 1926 3618 1930 3622
rect 2126 3618 2130 3622
rect 2150 3618 2154 3622
rect 2286 3618 2290 3622
rect 2390 3618 2394 3622
rect 2518 3618 2522 3622
rect 2678 3618 2682 3622
rect 2726 3618 2730 3622
rect 2998 3618 3002 3622
rect 3270 3618 3274 3622
rect 3430 3618 3434 3622
rect 3614 3618 3618 3622
rect 4350 3618 4354 3622
rect 4390 3618 4394 3622
rect 4518 3618 4522 3622
rect 4782 3618 4786 3622
rect 5214 3618 5218 3622
rect 346 3603 350 3607
rect 353 3603 357 3607
rect 1370 3603 1374 3607
rect 1377 3603 1381 3607
rect 2394 3603 2398 3607
rect 2401 3603 2405 3607
rect 3418 3603 3422 3607
rect 3425 3603 3429 3607
rect 4442 3603 4446 3607
rect 4449 3603 4453 3607
rect 174 3588 178 3592
rect 222 3588 226 3592
rect 286 3588 290 3592
rect 326 3588 330 3592
rect 622 3588 626 3592
rect 702 3588 706 3592
rect 830 3588 834 3592
rect 1158 3588 1162 3592
rect 1222 3588 1226 3592
rect 1478 3588 1482 3592
rect 1494 3588 1498 3592
rect 2270 3588 2274 3592
rect 2294 3588 2298 3592
rect 3094 3588 3098 3592
rect 3318 3588 3322 3592
rect 4118 3588 4122 3592
rect 4246 3588 4250 3592
rect 4734 3588 4738 3592
rect 4830 3588 4834 3592
rect 5246 3588 5250 3592
rect 758 3578 762 3582
rect 1574 3578 1578 3582
rect 4046 3578 4050 3582
rect 4134 3578 4138 3582
rect 166 3568 170 3572
rect 254 3568 258 3572
rect 670 3568 674 3572
rect 686 3568 690 3572
rect 750 3568 754 3572
rect 1046 3568 1050 3572
rect 1270 3568 1274 3572
rect 1318 3568 1322 3572
rect 1382 3568 1386 3572
rect 1518 3568 1522 3572
rect 1566 3568 1570 3572
rect 1758 3568 1762 3572
rect 1766 3568 1770 3572
rect 2166 3568 2170 3572
rect 2278 3568 2282 3572
rect 2454 3568 2458 3572
rect 2630 3568 2634 3572
rect 2670 3568 2674 3572
rect 2702 3568 2706 3572
rect 2718 3568 2722 3572
rect 3206 3568 3210 3572
rect 3222 3568 3226 3572
rect 4382 3568 4386 3572
rect 5222 3568 5226 3572
rect 5294 3568 5298 3572
rect 14 3558 18 3562
rect 94 3558 98 3562
rect 118 3558 122 3562
rect 198 3558 202 3562
rect 222 3558 226 3562
rect 230 3558 234 3562
rect 302 3558 306 3562
rect 390 3558 394 3562
rect 470 3558 474 3562
rect 638 3558 642 3562
rect 38 3548 42 3552
rect 54 3548 58 3552
rect 126 3548 130 3552
rect 174 3548 178 3552
rect 222 3548 226 3552
rect 286 3548 290 3552
rect 22 3538 26 3542
rect 398 3548 402 3552
rect 414 3548 418 3552
rect 470 3548 474 3552
rect 558 3548 562 3552
rect 574 3548 578 3552
rect 622 3548 626 3552
rect 646 3548 650 3552
rect 766 3558 770 3562
rect 942 3558 946 3562
rect 974 3558 978 3562
rect 1062 3558 1066 3562
rect 1070 3558 1074 3562
rect 1102 3558 1106 3562
rect 1134 3558 1138 3562
rect 1150 3558 1154 3562
rect 1166 3558 1170 3562
rect 1334 3558 1338 3562
rect 1398 3558 1402 3562
rect 1470 3558 1474 3562
rect 1550 3558 1554 3562
rect 1582 3558 1586 3562
rect 1686 3558 1690 3562
rect 1742 3558 1746 3562
rect 1750 3558 1754 3562
rect 1846 3558 1850 3562
rect 1886 3558 1890 3562
rect 1934 3558 1938 3562
rect 2030 3558 2034 3562
rect 2142 3558 2146 3562
rect 2150 3558 2154 3562
rect 2238 3558 2242 3562
rect 2254 3558 2258 3562
rect 2262 3558 2266 3562
rect 2366 3558 2370 3562
rect 2438 3558 2442 3562
rect 2494 3558 2498 3562
rect 2518 3558 2522 3562
rect 2550 3558 2554 3562
rect 2590 3558 2594 3562
rect 2614 3558 2618 3562
rect 2638 3558 2642 3562
rect 2654 3558 2658 3562
rect 2686 3558 2690 3562
rect 2734 3558 2738 3562
rect 2798 3558 2802 3562
rect 2854 3558 2858 3562
rect 2950 3558 2954 3562
rect 2966 3558 2970 3562
rect 3046 3558 3050 3562
rect 3070 3558 3074 3562
rect 710 3548 714 3552
rect 726 3548 730 3552
rect 758 3548 762 3552
rect 822 3548 826 3552
rect 878 3548 882 3552
rect 910 3548 914 3552
rect 926 3548 930 3552
rect 934 3548 938 3552
rect 958 3548 962 3552
rect 990 3548 994 3552
rect 1030 3548 1034 3552
rect 1038 3548 1042 3552
rect 1054 3548 1058 3552
rect 1086 3548 1090 3552
rect 1150 3548 1154 3552
rect 1246 3548 1250 3552
rect 1278 3548 1282 3552
rect 1326 3548 1330 3552
rect 1390 3548 1394 3552
rect 1406 3548 1410 3552
rect 1446 3548 1450 3552
rect 1510 3548 1514 3552
rect 118 3538 122 3542
rect 134 3538 138 3542
rect 294 3538 298 3542
rect 318 3538 322 3542
rect 342 3538 346 3542
rect 374 3538 378 3542
rect 446 3538 450 3542
rect 454 3538 458 3542
rect 1590 3548 1594 3552
rect 1662 3548 1666 3552
rect 1710 3548 1714 3552
rect 1758 3548 1762 3552
rect 1782 3548 1786 3552
rect 1814 3548 1818 3552
rect 1862 3548 1866 3552
rect 1918 3548 1922 3552
rect 1942 3548 1946 3552
rect 2014 3548 2018 3552
rect 2046 3548 2050 3552
rect 2158 3548 2162 3552
rect 2182 3548 2186 3552
rect 2222 3548 2226 3552
rect 2270 3548 2274 3552
rect 2310 3548 2314 3552
rect 2350 3548 2354 3552
rect 2366 3548 2370 3552
rect 2406 3548 2410 3552
rect 2446 3548 2450 3552
rect 2470 3548 2474 3552
rect 3750 3557 3754 3561
rect 3894 3557 3898 3561
rect 4230 3558 4234 3562
rect 4358 3558 4362 3562
rect 4398 3558 4402 3562
rect 4662 3558 4666 3562
rect 4694 3558 4698 3562
rect 4710 3558 4714 3562
rect 4766 3558 4770 3562
rect 5126 3558 5130 3562
rect 5286 3558 5290 3562
rect 2574 3548 2578 3552
rect 2590 3548 2594 3552
rect 2678 3548 2682 3552
rect 2694 3548 2698 3552
rect 2726 3548 2730 3552
rect 2742 3548 2746 3552
rect 2774 3548 2778 3552
rect 2830 3548 2834 3552
rect 2958 3548 2962 3552
rect 2990 3548 2994 3552
rect 3078 3548 3082 3552
rect 3110 3548 3114 3552
rect 3118 3548 3122 3552
rect 3126 3548 3130 3552
rect 3158 3548 3162 3552
rect 3190 3548 3194 3552
rect 3198 3548 3202 3552
rect 478 3538 482 3542
rect 526 3538 530 3542
rect 550 3538 554 3542
rect 566 3538 570 3542
rect 614 3538 618 3542
rect 686 3538 690 3542
rect 734 3538 738 3542
rect 790 3538 794 3542
rect 822 3538 826 3542
rect 910 3538 914 3542
rect 918 3538 922 3542
rect 950 3538 954 3542
rect 1102 3538 1106 3542
rect 1118 3538 1122 3542
rect 1166 3538 1170 3542
rect 1190 3538 1194 3542
rect 1238 3538 1242 3542
rect 1286 3538 1290 3542
rect 1414 3538 1418 3542
rect 1438 3538 1442 3542
rect 1454 3538 1458 3542
rect 1486 3538 1490 3542
rect 1534 3538 1538 3542
rect 1550 3538 1554 3542
rect 1574 3538 1578 3542
rect 1598 3538 1602 3542
rect 1614 3538 1618 3542
rect 1654 3538 1658 3542
rect 3270 3547 3274 3551
rect 3302 3548 3306 3552
rect 3334 3548 3338 3552
rect 3350 3548 3354 3552
rect 3358 3548 3362 3552
rect 3398 3548 3402 3552
rect 3446 3548 3450 3552
rect 3494 3548 3498 3552
rect 3566 3547 3570 3551
rect 3598 3548 3602 3552
rect 3630 3548 3634 3552
rect 3638 3548 3642 3552
rect 3670 3548 3674 3552
rect 3718 3548 3722 3552
rect 3758 3548 3762 3552
rect 3806 3548 3810 3552
rect 3814 3548 3818 3552
rect 3846 3548 3850 3552
rect 3854 3548 3858 3552
rect 3950 3548 3954 3552
rect 3982 3547 3986 3551
rect 4006 3548 4010 3552
rect 4086 3548 4090 3552
rect 4094 3548 4098 3552
rect 4102 3548 4106 3552
rect 4174 3548 4178 3552
rect 4190 3548 4194 3552
rect 4206 3548 4210 3552
rect 4310 3548 4314 3552
rect 4374 3548 4378 3552
rect 4510 3548 4514 3552
rect 4526 3548 4530 3552
rect 4542 3548 4546 3552
rect 4558 3548 4562 3552
rect 4590 3548 4594 3552
rect 4614 3548 4618 3552
rect 4646 3548 4650 3552
rect 4670 3548 4674 3552
rect 4718 3548 4722 3552
rect 4750 3548 4754 3552
rect 4774 3548 4778 3552
rect 4838 3548 4842 3552
rect 4846 3548 4850 3552
rect 4862 3548 4866 3552
rect 4878 3548 4882 3552
rect 4950 3548 4954 3552
rect 5022 3548 5026 3552
rect 5030 3548 5034 3552
rect 5062 3548 5066 3552
rect 5094 3548 5098 3552
rect 1718 3538 1722 3542
rect 1726 3538 1730 3542
rect 1742 3538 1746 3542
rect 1822 3538 1826 3542
rect 1854 3538 1858 3542
rect 1870 3538 1874 3542
rect 1902 3538 1906 3542
rect 1910 3538 1914 3542
rect 1926 3538 1930 3542
rect 1958 3538 1962 3542
rect 2006 3538 2010 3542
rect 2070 3538 2074 3542
rect 2118 3538 2122 3542
rect 2126 3538 2130 3542
rect 2190 3538 2194 3542
rect 2214 3538 2218 3542
rect 2318 3538 2322 3542
rect 2342 3538 2346 3542
rect 2414 3538 2418 3542
rect 2486 3538 2490 3542
rect 2510 3538 2514 3542
rect 2534 3538 2538 3542
rect 2566 3538 2570 3542
rect 2598 3538 2602 3542
rect 2630 3538 2634 3542
rect 2654 3538 2658 3542
rect 2718 3538 2722 3542
rect 2750 3538 2754 3542
rect 2766 3538 2770 3542
rect 2782 3538 2786 3542
rect 2822 3538 2826 3542
rect 2830 3538 2834 3542
rect 2854 3538 2858 3542
rect 2862 3538 2866 3542
rect 2910 3538 2914 3542
rect 2974 3538 2978 3542
rect 2998 3538 3002 3542
rect 3014 3538 3018 3542
rect 3030 3538 3034 3542
rect 3054 3538 3058 3542
rect 3070 3538 3074 3542
rect 3134 3538 3138 3542
rect 3150 3538 3154 3542
rect 3254 3538 3258 3542
rect 3414 3538 3418 3542
rect 3454 3538 3458 3542
rect 3534 3538 3538 3542
rect 3582 3538 3586 3542
rect 3662 3538 3666 3542
rect 3726 3538 3730 3542
rect 3766 3538 3770 3542
rect 3822 3538 3826 3542
rect 3918 3538 3922 3542
rect 3966 3538 3970 3542
rect 4054 3538 4058 3542
rect 4150 3538 4154 3542
rect 4166 3538 4170 3542
rect 4182 3538 4186 3542
rect 4302 3538 4306 3542
rect 4318 3538 4322 3542
rect 4342 3538 4346 3542
rect 4398 3538 4402 3542
rect 4414 3538 4418 3542
rect 4422 3538 4426 3542
rect 4446 3538 4450 3542
rect 4462 3538 4466 3542
rect 4486 3538 4490 3542
rect 4502 3538 4506 3542
rect 4518 3538 4522 3542
rect 4558 3538 4562 3542
rect 4582 3538 4586 3542
rect 5158 3547 5162 3551
rect 5254 3548 5258 3552
rect 5286 3548 5290 3552
rect 4614 3538 4618 3542
rect 4630 3538 4634 3542
rect 4638 3538 4642 3542
rect 4710 3538 4714 3542
rect 4806 3538 4810 3542
rect 4854 3538 4858 3542
rect 4894 3538 4898 3542
rect 4918 3538 4922 3542
rect 4942 3538 4946 3542
rect 5014 3538 5018 3542
rect 5142 3538 5146 3542
rect 6 3528 10 3532
rect 70 3528 74 3532
rect 150 3528 154 3532
rect 198 3528 202 3532
rect 246 3528 250 3532
rect 254 3528 258 3532
rect 310 3528 314 3532
rect 326 3528 330 3532
rect 534 3528 538 3532
rect 542 3528 546 3532
rect 606 3528 610 3532
rect 662 3528 666 3532
rect 774 3528 778 3532
rect 870 3528 874 3532
rect 1102 3528 1106 3532
rect 1126 3528 1130 3532
rect 1182 3528 1186 3532
rect 1302 3528 1306 3532
rect 1350 3528 1354 3532
rect 1430 3528 1434 3532
rect 1470 3528 1474 3532
rect 1478 3528 1482 3532
rect 1526 3528 1530 3532
rect 1614 3528 1618 3532
rect 1622 3528 1626 3532
rect 1758 3528 1762 3532
rect 1838 3528 1842 3532
rect 1950 3528 1954 3532
rect 2206 3528 2210 3532
rect 2238 3528 2242 3532
rect 2254 3528 2258 3532
rect 2302 3528 2306 3532
rect 2334 3528 2338 3532
rect 2374 3528 2378 3532
rect 2390 3528 2394 3532
rect 2430 3528 2434 3532
rect 2486 3528 2490 3532
rect 2542 3528 2546 3532
rect 2678 3528 2682 3532
rect 2694 3528 2698 3532
rect 2974 3528 2978 3532
rect 3142 3528 3146 3532
rect 3150 3528 3154 3532
rect 3462 3528 3466 3532
rect 3486 3527 3490 3531
rect 3622 3528 3626 3532
rect 3670 3528 3674 3532
rect 3726 3528 3730 3532
rect 3862 3527 3866 3531
rect 3918 3528 3922 3532
rect 4126 3528 4130 3532
rect 4230 3528 4234 3532
rect 4334 3528 4338 3532
rect 4670 3528 4674 3532
rect 4774 3528 4778 3532
rect 5070 3528 5074 3532
rect 5270 3528 5274 3532
rect 22 3518 26 3522
rect 94 3518 98 3522
rect 142 3518 146 3522
rect 510 3518 514 3522
rect 590 3518 594 3522
rect 726 3518 730 3522
rect 1006 3518 1010 3522
rect 1294 3518 1298 3522
rect 1326 3518 1330 3522
rect 1390 3518 1394 3522
rect 1422 3518 1426 3522
rect 1646 3518 1650 3522
rect 1686 3518 1690 3522
rect 1694 3518 1698 3522
rect 1782 3518 1786 3522
rect 1958 3518 1962 3522
rect 2094 3518 2098 3522
rect 2134 3518 2138 3522
rect 2158 3518 2162 3522
rect 2198 3518 2202 3522
rect 2326 3518 2330 3522
rect 2350 3518 2354 3522
rect 2422 3518 2426 3522
rect 2454 3518 2458 3522
rect 2518 3518 2522 3522
rect 2614 3518 2618 3522
rect 2766 3518 2770 3522
rect 2814 3518 2818 3522
rect 2894 3518 2898 3522
rect 2950 3518 2954 3522
rect 3038 3518 3042 3522
rect 3454 3518 3458 3522
rect 3502 3518 3506 3522
rect 3662 3518 3666 3522
rect 4158 3518 4162 3522
rect 4190 3518 4194 3522
rect 4326 3518 4330 3522
rect 4382 3518 4386 3522
rect 4470 3518 4474 3522
rect 4494 3518 4498 3522
rect 4526 3518 4530 3522
rect 4574 3518 4578 3522
rect 4662 3518 4666 3522
rect 4878 3518 4882 3522
rect 4918 3518 4922 3522
rect 4998 3518 5002 3522
rect 5262 3518 5266 3522
rect 5286 3518 5290 3522
rect 6 3508 10 3512
rect 438 3508 442 3512
rect 662 3508 666 3512
rect 1126 3508 1130 3512
rect 1166 3508 1170 3512
rect 1254 3508 1258 3512
rect 1526 3508 1530 3512
rect 2078 3508 2082 3512
rect 2486 3508 2490 3512
rect 2630 3508 2634 3512
rect 2782 3508 2786 3512
rect 2838 3508 2842 3512
rect 2974 3508 2978 3512
rect 5254 3508 5258 3512
rect 858 3503 862 3507
rect 865 3503 869 3507
rect 1874 3503 1878 3507
rect 1881 3503 1885 3507
rect 2906 3503 2910 3507
rect 2913 3503 2917 3507
rect 3930 3503 3934 3507
rect 3937 3503 3941 3507
rect 4954 3503 4958 3507
rect 4961 3503 4965 3507
rect 614 3498 618 3502
rect 806 3498 810 3502
rect 1086 3498 1090 3502
rect 1438 3498 1442 3502
rect 1846 3498 1850 3502
rect 38 3488 42 3492
rect 70 3488 74 3492
rect 270 3488 274 3492
rect 414 3488 418 3492
rect 494 3488 498 3492
rect 582 3488 586 3492
rect 710 3488 714 3492
rect 718 3488 722 3492
rect 790 3488 794 3492
rect 814 3488 818 3492
rect 862 3488 866 3492
rect 926 3488 930 3492
rect 998 3488 1002 3492
rect 1014 3488 1018 3492
rect 1054 3488 1058 3492
rect 1118 3488 1122 3492
rect 1190 3488 1194 3492
rect 1214 3488 1218 3492
rect 1238 3488 1242 3492
rect 1286 3488 1290 3492
rect 1638 3488 1642 3492
rect 1806 3488 1810 3492
rect 1918 3488 1922 3492
rect 2062 3488 2066 3492
rect 2158 3488 2162 3492
rect 2262 3488 2266 3492
rect 2598 3488 2602 3492
rect 2662 3488 2666 3492
rect 2822 3488 2826 3492
rect 2902 3488 2906 3492
rect 2990 3488 2994 3492
rect 3022 3488 3026 3492
rect 3078 3488 3082 3492
rect 3190 3488 3194 3492
rect 3374 3488 3378 3492
rect 3398 3488 3402 3492
rect 3606 3488 3610 3492
rect 3630 3488 3634 3492
rect 3782 3488 3786 3492
rect 3870 3488 3874 3492
rect 3910 3488 3914 3492
rect 4070 3488 4074 3492
rect 4110 3488 4114 3492
rect 4174 3488 4178 3492
rect 4710 3488 4714 3492
rect 4734 3488 4738 3492
rect 4766 3488 4770 3492
rect 4894 3488 4898 3492
rect 5206 3488 5210 3492
rect 5230 3488 5234 3492
rect 174 3478 178 3482
rect 182 3478 186 3482
rect 326 3478 330 3482
rect 462 3478 466 3482
rect 518 3478 522 3482
rect 534 3478 538 3482
rect 550 3478 554 3482
rect 590 3478 594 3482
rect 662 3478 666 3482
rect 806 3478 810 3482
rect 846 3478 850 3482
rect 934 3478 938 3482
rect 950 3478 954 3482
rect 1086 3478 1090 3482
rect 1134 3478 1138 3482
rect 1406 3478 1410 3482
rect 1430 3478 1434 3482
rect 1438 3478 1442 3482
rect 1662 3478 1666 3482
rect 1694 3478 1698 3482
rect 1814 3478 1818 3482
rect 1846 3478 1850 3482
rect 1854 3478 1858 3482
rect 1926 3478 1930 3482
rect 1966 3478 1970 3482
rect 2134 3478 2138 3482
rect 2302 3478 2306 3482
rect 2366 3478 2370 3482
rect 2462 3478 2466 3482
rect 2542 3478 2546 3482
rect 2590 3478 2594 3482
rect 2718 3478 2722 3482
rect 2878 3478 2882 3482
rect 2894 3478 2898 3482
rect 2966 3478 2970 3482
rect 3102 3478 3106 3482
rect 3150 3478 3154 3482
rect 3158 3478 3162 3482
rect 3254 3478 3258 3482
rect 3502 3479 3506 3483
rect 3630 3478 3634 3482
rect 3686 3478 3690 3482
rect 3830 3478 3834 3482
rect 4054 3478 4058 3482
rect 4142 3478 4146 3482
rect 4294 3478 4298 3482
rect 4358 3478 4362 3482
rect 4406 3478 4410 3482
rect 4422 3478 4426 3482
rect 4478 3478 4482 3482
rect 4494 3478 4498 3482
rect 4526 3478 4530 3482
rect 4574 3478 4578 3482
rect 4774 3478 4778 3482
rect 5070 3478 5074 3482
rect 5142 3478 5146 3482
rect 6 3468 10 3472
rect 54 3468 58 3472
rect 62 3468 66 3472
rect 94 3468 98 3472
rect 102 3468 106 3472
rect 150 3468 154 3472
rect 230 3468 234 3472
rect 246 3468 250 3472
rect 318 3468 322 3472
rect 358 3468 362 3472
rect 446 3468 450 3472
rect 478 3468 482 3472
rect 566 3468 570 3472
rect 614 3468 618 3472
rect 630 3468 634 3472
rect 638 3468 642 3472
rect 702 3468 706 3472
rect 750 3468 754 3472
rect 766 3468 770 3472
rect 790 3468 794 3472
rect 830 3468 834 3472
rect 854 3468 858 3472
rect 862 3468 866 3472
rect 918 3468 922 3472
rect 958 3468 962 3472
rect 1006 3468 1010 3472
rect 1038 3468 1042 3472
rect 1046 3468 1050 3472
rect 1086 3468 1090 3472
rect 1126 3468 1130 3472
rect 1166 3468 1170 3472
rect 1198 3468 1202 3472
rect 1246 3468 1250 3472
rect 1254 3468 1258 3472
rect 1302 3468 1306 3472
rect 1390 3468 1394 3472
rect 1454 3468 1458 3472
rect 1486 3468 1490 3472
rect 1518 3468 1522 3472
rect 1526 3468 1530 3472
rect 1574 3468 1578 3472
rect 1606 3468 1610 3472
rect 1662 3468 1666 3472
rect 1678 3468 1682 3472
rect 1686 3468 1690 3472
rect 1742 3468 1746 3472
rect 1854 3468 1858 3472
rect 1870 3468 1874 3472
rect 1894 3468 1898 3472
rect 22 3458 26 3462
rect 70 3458 74 3462
rect 126 3458 130 3462
rect 150 3458 154 3462
rect 206 3458 210 3462
rect 254 3458 258 3462
rect 310 3458 314 3462
rect 318 3458 322 3462
rect 398 3458 402 3462
rect 438 3458 442 3462
rect 446 3458 450 3462
rect 478 3458 482 3462
rect 494 3458 498 3462
rect 550 3458 554 3462
rect 614 3458 618 3462
rect 638 3458 642 3462
rect 678 3458 682 3462
rect 790 3458 794 3462
rect 854 3458 858 3462
rect 1006 3458 1010 3462
rect 1030 3458 1034 3462
rect 1070 3458 1074 3462
rect 1102 3458 1106 3462
rect 1158 3458 1162 3462
rect 1174 3458 1178 3462
rect 1318 3458 1322 3462
rect 1326 3458 1330 3462
rect 1350 3458 1354 3462
rect 1414 3458 1418 3462
rect 1462 3458 1466 3462
rect 1510 3458 1514 3462
rect 1598 3458 1602 3462
rect 1686 3458 1690 3462
rect 1710 3458 1714 3462
rect 1734 3458 1738 3462
rect 1766 3458 1770 3462
rect 1790 3458 1794 3462
rect 1814 3458 1818 3462
rect 1830 3458 1834 3462
rect 1902 3466 1906 3470
rect 1966 3468 1970 3472
rect 2022 3468 2026 3472
rect 2030 3468 2034 3472
rect 2078 3468 2082 3472
rect 2086 3468 2090 3472
rect 2102 3468 2106 3472
rect 2118 3468 2122 3472
rect 2142 3468 2146 3472
rect 2222 3468 2226 3472
rect 2230 3468 2234 3472
rect 2278 3468 2282 3472
rect 2310 3468 2314 3472
rect 2358 3468 2362 3472
rect 2390 3468 2394 3472
rect 2406 3468 2410 3472
rect 1942 3458 1946 3462
rect 2110 3458 2114 3462
rect 2214 3458 2218 3462
rect 2286 3458 2290 3462
rect 2350 3458 2354 3462
rect 2382 3458 2386 3462
rect 2494 3468 2498 3472
rect 2534 3468 2538 3472
rect 2630 3468 2634 3472
rect 2638 3468 2642 3472
rect 2734 3468 2738 3472
rect 2782 3468 2786 3472
rect 2790 3468 2794 3472
rect 2838 3468 2842 3472
rect 2870 3468 2874 3472
rect 2958 3468 2962 3472
rect 2966 3468 2970 3472
rect 2982 3468 2986 3472
rect 2990 3468 2994 3472
rect 3070 3468 3074 3472
rect 3182 3468 3186 3472
rect 3478 3468 3482 3472
rect 3630 3468 3634 3472
rect 3710 3468 3714 3472
rect 3774 3468 3778 3472
rect 3838 3468 3842 3472
rect 3966 3468 3970 3472
rect 4054 3468 4058 3472
rect 4190 3468 4194 3472
rect 4214 3468 4218 3472
rect 4246 3468 4250 3472
rect 2462 3458 2466 3462
rect 2478 3458 2482 3462
rect 2494 3458 2498 3462
rect 2526 3458 2530 3462
rect 2574 3458 2578 3462
rect 2606 3458 2610 3462
rect 2622 3458 2626 3462
rect 2646 3458 2650 3462
rect 2686 3458 2690 3462
rect 2694 3458 2698 3462
rect 2878 3458 2882 3462
rect 2894 3458 2898 3462
rect 2910 3458 2914 3462
rect 2958 3458 2962 3462
rect 2990 3458 2994 3462
rect 3006 3458 3010 3462
rect 3014 3458 3018 3462
rect 3046 3458 3050 3462
rect 3062 3458 3066 3462
rect 3118 3458 3122 3462
rect 3174 3458 3178 3462
rect 3254 3459 3258 3463
rect 3326 3458 3330 3462
rect 3342 3458 3346 3462
rect 3454 3458 3458 3462
rect 3494 3458 3498 3462
rect 3542 3459 3546 3463
rect 3574 3458 3578 3462
rect 3638 3458 3642 3462
rect 3702 3458 3706 3462
rect 3798 3458 3802 3462
rect 3830 3458 3834 3462
rect 3854 3458 3858 3462
rect 3886 3458 3890 3462
rect 3974 3459 3978 3463
rect 4038 3458 4042 3462
rect 4086 3458 4090 3462
rect 4094 3458 4098 3462
rect 4118 3458 4122 3462
rect 4174 3458 4178 3462
rect 4190 3458 4194 3462
rect 4222 3458 4226 3462
rect 4230 3458 4234 3462
rect 4238 3458 4242 3462
rect 4310 3468 4314 3472
rect 4326 3468 4330 3472
rect 4350 3468 4354 3472
rect 4374 3468 4378 3472
rect 4414 3468 4418 3472
rect 4462 3468 4466 3472
rect 4486 3468 4490 3472
rect 4518 3468 4522 3472
rect 4566 3468 4570 3472
rect 4614 3468 4618 3472
rect 4646 3468 4650 3472
rect 4654 3468 4658 3472
rect 4798 3468 4802 3472
rect 4830 3468 4834 3472
rect 4270 3458 4274 3462
rect 4278 3458 4282 3462
rect 4302 3458 4306 3462
rect 4334 3458 4338 3462
rect 4382 3458 4386 3462
rect 4390 3458 4394 3462
rect 4406 3458 4410 3462
rect 4438 3458 4442 3462
rect 4494 3458 4498 3462
rect 4510 3458 4514 3462
rect 4542 3458 4546 3462
rect 4590 3458 4594 3462
rect 4750 3458 4754 3462
rect 4758 3458 4762 3462
rect 4790 3458 4794 3462
rect 4798 3458 4802 3462
rect 4822 3458 4826 3462
rect 4862 3468 4866 3472
rect 4878 3468 4882 3472
rect 4910 3468 4914 3472
rect 4918 3468 4922 3472
rect 4934 3468 4938 3472
rect 4942 3468 4946 3472
rect 4998 3468 5002 3472
rect 4854 3458 4858 3462
rect 4886 3458 4890 3462
rect 5006 3458 5010 3462
rect 5014 3458 5018 3462
rect 5062 3458 5066 3462
rect 5078 3458 5082 3462
rect 5142 3459 5146 3463
rect 5254 3458 5258 3462
rect 5270 3458 5274 3462
rect 86 3448 90 3452
rect 110 3448 114 3452
rect 118 3448 122 3452
rect 238 3448 242 3452
rect 278 3448 282 3452
rect 390 3448 394 3452
rect 486 3448 490 3452
rect 566 3448 570 3452
rect 582 3448 586 3452
rect 630 3448 634 3452
rect 670 3448 674 3452
rect 814 3448 818 3452
rect 838 3448 842 3452
rect 902 3448 906 3452
rect 942 3448 946 3452
rect 1062 3448 1066 3452
rect 1118 3448 1122 3452
rect 1190 3448 1194 3452
rect 1334 3448 1338 3452
rect 1342 3448 1346 3452
rect 1406 3448 1410 3452
rect 1422 3448 1426 3452
rect 1486 3448 1490 3452
rect 1494 3448 1498 3452
rect 1510 3448 1514 3452
rect 1598 3448 1602 3452
rect 1718 3448 1722 3452
rect 1750 3448 1754 3452
rect 1774 3448 1778 3452
rect 2102 3448 2106 3452
rect 2198 3448 2202 3452
rect 2294 3448 2298 3452
rect 2326 3448 2330 3452
rect 2334 3448 2338 3452
rect 2462 3448 2466 3452
rect 2582 3448 2586 3452
rect 2662 3448 2666 3452
rect 2846 3448 2850 3452
rect 2934 3448 2938 3452
rect 3022 3448 3026 3452
rect 3054 3448 3058 3452
rect 3110 3448 3114 3452
rect 3142 3448 3146 3452
rect 3158 3448 3162 3452
rect 4182 3448 4186 3452
rect 4206 3448 4210 3452
rect 4270 3448 4274 3452
rect 4286 3448 4290 3452
rect 4326 3448 4330 3452
rect 4366 3448 4370 3452
rect 4478 3448 4482 3452
rect 4550 3448 4554 3452
rect 4630 3448 4634 3452
rect 4774 3448 4778 3452
rect 4806 3448 4810 3452
rect 4878 3448 4882 3452
rect 4894 3448 4898 3452
rect 5110 3448 5114 3452
rect 5262 3448 5266 3452
rect 134 3438 138 3442
rect 182 3438 186 3442
rect 214 3438 218 3442
rect 286 3438 290 3442
rect 502 3438 506 3442
rect 534 3438 538 3442
rect 686 3438 690 3442
rect 758 3438 762 3442
rect 1358 3438 1362 3442
rect 1438 3438 1442 3442
rect 1558 3438 1562 3442
rect 1758 3438 1762 3442
rect 1814 3438 1818 3442
rect 2134 3438 2138 3442
rect 2566 3438 2570 3442
rect 3038 3438 3042 3442
rect 3046 3438 3050 3442
rect 3126 3438 3130 3442
rect 4166 3438 4170 3442
rect 4254 3438 4258 3442
rect 4342 3438 4346 3442
rect 4454 3438 4458 3442
rect 4566 3438 4570 3442
rect 5190 3438 5194 3442
rect 5278 3438 5282 3442
rect 1374 3428 1378 3432
rect 3134 3428 3138 3432
rect 126 3418 130 3422
rect 190 3418 194 3422
rect 206 3418 210 3422
rect 606 3418 610 3422
rect 662 3418 666 3422
rect 694 3418 698 3422
rect 1662 3418 1666 3422
rect 1734 3418 1738 3422
rect 1958 3418 1962 3422
rect 2006 3418 2010 3422
rect 2318 3418 2322 3422
rect 2350 3418 2354 3422
rect 2438 3418 2442 3422
rect 2574 3418 2578 3422
rect 2726 3418 2730 3422
rect 2766 3418 2770 3422
rect 2862 3418 2866 3422
rect 2950 3418 2954 3422
rect 4014 3418 4018 3422
rect 4542 3418 4546 3422
rect 4598 3418 4602 3422
rect 4710 3418 4714 3422
rect 4926 3418 4930 3422
rect 4982 3418 4986 3422
rect 5270 3418 5274 3422
rect 346 3403 350 3407
rect 353 3403 357 3407
rect 1370 3403 1374 3407
rect 1377 3403 1381 3407
rect 2394 3403 2398 3407
rect 2401 3403 2405 3407
rect 3418 3403 3422 3407
rect 3425 3403 3429 3407
rect 4442 3403 4446 3407
rect 4449 3403 4453 3407
rect 142 3388 146 3392
rect 174 3388 178 3392
rect 422 3388 426 3392
rect 526 3388 530 3392
rect 582 3388 586 3392
rect 670 3388 674 3392
rect 854 3388 858 3392
rect 1462 3388 1466 3392
rect 1558 3388 1562 3392
rect 1870 3388 1874 3392
rect 2086 3388 2090 3392
rect 2126 3388 2130 3392
rect 2622 3388 2626 3392
rect 2630 3388 2634 3392
rect 3030 3388 3034 3392
rect 3198 3388 3202 3392
rect 3342 3388 3346 3392
rect 3398 3388 3402 3392
rect 3574 3388 3578 3392
rect 3686 3388 3690 3392
rect 4222 3388 4226 3392
rect 4502 3388 4506 3392
rect 4798 3388 4802 3392
rect 5246 3388 5250 3392
rect 446 3378 450 3382
rect 558 3378 562 3382
rect 1166 3378 1170 3382
rect 1182 3378 1186 3382
rect 1518 3378 1522 3382
rect 2318 3378 2322 3382
rect 2582 3378 2586 3382
rect 78 3368 82 3372
rect 134 3368 138 3372
rect 166 3368 170 3372
rect 430 3368 434 3372
rect 534 3368 538 3372
rect 630 3368 634 3372
rect 782 3368 786 3372
rect 1078 3368 1082 3372
rect 1158 3368 1162 3372
rect 1566 3368 1570 3372
rect 1774 3368 1778 3372
rect 1846 3368 1850 3372
rect 2094 3368 2098 3372
rect 2134 3368 2138 3372
rect 2158 3368 2162 3372
rect 2318 3368 2322 3372
rect 2326 3368 2330 3372
rect 2614 3368 2618 3372
rect 2638 3368 2642 3372
rect 2814 3368 2818 3372
rect 2958 3368 2962 3372
rect 3206 3368 3210 3372
rect 3550 3368 3554 3372
rect 3590 3368 3594 3372
rect 3966 3368 3970 3372
rect 4118 3368 4122 3372
rect 4790 3368 4794 3372
rect 4806 3368 4810 3372
rect 4838 3368 4842 3372
rect 5110 3368 5114 3372
rect 5118 3368 5122 3372
rect 5134 3368 5138 3372
rect 54 3358 58 3362
rect 62 3358 66 3362
rect 118 3358 122 3362
rect 150 3358 154 3362
rect 286 3358 290 3362
rect 382 3358 386 3362
rect 414 3358 418 3362
rect 478 3358 482 3362
rect 518 3358 522 3362
rect 550 3358 554 3362
rect 574 3358 578 3362
rect 710 3358 714 3362
rect 766 3358 770 3362
rect 798 3358 802 3362
rect 814 3358 818 3362
rect 1006 3358 1010 3362
rect 1014 3358 1018 3362
rect 1030 3358 1034 3362
rect 1062 3358 1066 3362
rect 1094 3358 1098 3362
rect 1110 3358 1114 3362
rect 1454 3358 1458 3362
rect 1510 3358 1514 3362
rect 1542 3358 1546 3362
rect 1550 3358 1554 3362
rect 1582 3358 1586 3362
rect 1830 3358 1834 3362
rect 6 3348 10 3352
rect 30 3348 34 3352
rect 110 3348 114 3352
rect 126 3348 130 3352
rect 182 3348 186 3352
rect 254 3348 258 3352
rect 302 3348 306 3352
rect 22 3338 26 3342
rect 166 3338 170 3342
rect 198 3338 202 3342
rect 262 3338 266 3342
rect 294 3338 298 3342
rect 310 3338 314 3342
rect 358 3348 362 3352
rect 406 3348 410 3352
rect 422 3348 426 3352
rect 406 3338 410 3342
rect 462 3340 466 3344
rect 526 3348 530 3352
rect 630 3348 634 3352
rect 646 3348 650 3352
rect 686 3348 690 3352
rect 774 3348 778 3352
rect 894 3348 898 3352
rect 950 3348 954 3352
rect 1030 3348 1034 3352
rect 1054 3348 1058 3352
rect 1070 3348 1074 3352
rect 1142 3348 1146 3352
rect 1166 3348 1170 3352
rect 1230 3348 1234 3352
rect 1254 3348 1258 3352
rect 1278 3348 1282 3352
rect 1422 3348 1426 3352
rect 1446 3348 1450 3352
rect 1486 3348 1490 3352
rect 1502 3348 1506 3352
rect 1542 3348 1546 3352
rect 1558 3348 1562 3352
rect 1598 3348 1602 3352
rect 1630 3348 1634 3352
rect 1710 3348 1714 3352
rect 1774 3348 1778 3352
rect 1838 3348 1842 3352
rect 1862 3348 1866 3352
rect 1902 3348 1906 3352
rect 1926 3348 1930 3352
rect 2006 3348 2010 3352
rect 2078 3358 2082 3362
rect 2110 3358 2114 3362
rect 2126 3358 2130 3362
rect 2590 3358 2594 3362
rect 2598 3358 2602 3362
rect 2654 3358 2658 3362
rect 2678 3358 2682 3362
rect 2694 3358 2698 3362
rect 2726 3358 2730 3362
rect 2958 3358 2962 3362
rect 2974 3358 2978 3362
rect 3062 3358 3066 3362
rect 3094 3358 3098 3362
rect 3134 3358 3138 3362
rect 3190 3358 3194 3362
rect 3222 3358 3226 3362
rect 3286 3358 3290 3362
rect 4086 3358 4090 3362
rect 4238 3358 4242 3362
rect 4390 3358 4394 3362
rect 2062 3348 2066 3352
rect 2078 3348 2082 3352
rect 2102 3348 2106 3352
rect 2134 3348 2138 3352
rect 2166 3348 2170 3352
rect 2198 3348 2202 3352
rect 2278 3348 2282 3352
rect 2318 3348 2322 3352
rect 2342 3348 2346 3352
rect 2422 3348 2426 3352
rect 2518 3348 2522 3352
rect 2566 3348 2570 3352
rect 2606 3348 2610 3352
rect 2646 3348 2650 3352
rect 2742 3348 2746 3352
rect 2758 3348 2762 3352
rect 2838 3348 2842 3352
rect 2862 3348 2866 3352
rect 2966 3348 2970 3352
rect 2990 3348 2994 3352
rect 3046 3348 3050 3352
rect 3086 3348 3090 3352
rect 3142 3348 3146 3352
rect 3214 3348 3218 3352
rect 3246 3348 3250 3352
rect 3318 3348 3322 3352
rect 3358 3348 3362 3352
rect 3494 3348 3498 3352
rect 3630 3348 3634 3352
rect 3670 3348 3674 3352
rect 3702 3348 3706 3352
rect 3710 3348 3714 3352
rect 3774 3348 3778 3352
rect 3814 3348 3818 3352
rect 3822 3348 3826 3352
rect 3846 3348 3850 3352
rect 3886 3348 3890 3352
rect 3918 3348 3922 3352
rect 4030 3348 4034 3352
rect 4078 3348 4082 3352
rect 4102 3348 4106 3352
rect 4110 3348 4114 3352
rect 4174 3348 4178 3352
rect 494 3340 498 3344
rect 566 3338 570 3342
rect 638 3338 642 3342
rect 686 3338 690 3342
rect 718 3338 722 3342
rect 726 3340 730 3344
rect 750 3338 754 3342
rect 798 3338 802 3342
rect 814 3338 818 3342
rect 822 3338 826 3342
rect 870 3338 874 3342
rect 918 3338 922 3342
rect 966 3338 970 3342
rect 974 3338 978 3342
rect 990 3338 994 3342
rect 1038 3338 1042 3342
rect 1094 3338 1098 3342
rect 1118 3338 1122 3342
rect 1134 3338 1138 3342
rect 1222 3338 1226 3342
rect 1238 3338 1242 3342
rect 1246 3338 1250 3342
rect 1302 3338 1306 3342
rect 1350 3338 1354 3342
rect 1374 3338 1378 3342
rect 1430 3338 1434 3342
rect 1454 3338 1458 3342
rect 1470 3338 1474 3342
rect 1478 3338 1482 3342
rect 1590 3338 1594 3342
rect 1622 3338 1626 3342
rect 1654 3338 1658 3342
rect 1702 3338 1706 3342
rect 1750 3338 1754 3342
rect 1782 3338 1786 3342
rect 1798 3338 1802 3342
rect 1894 3338 1898 3342
rect 1950 3338 1954 3342
rect 1998 3338 2002 3342
rect 2046 3338 2050 3342
rect 2054 3338 2058 3342
rect 2174 3338 2178 3342
rect 2190 3338 2194 3342
rect 2206 3338 2210 3342
rect 4278 3347 4282 3351
rect 4390 3348 4394 3352
rect 4446 3358 4450 3362
rect 4614 3358 4618 3362
rect 4670 3358 4674 3362
rect 4822 3358 4826 3362
rect 4894 3358 4898 3362
rect 4910 3358 4914 3362
rect 5014 3358 5018 3362
rect 5094 3358 5098 3362
rect 5102 3358 5106 3362
rect 5270 3358 5274 3362
rect 4462 3348 4466 3352
rect 4478 3348 4482 3352
rect 4558 3348 4562 3352
rect 4654 3348 4658 3352
rect 4694 3348 4698 3352
rect 4734 3348 4738 3352
rect 4814 3348 4818 3352
rect 4846 3348 4850 3352
rect 4862 3348 4866 3352
rect 4878 3348 4882 3352
rect 4982 3348 4986 3352
rect 4990 3348 4994 3352
rect 5022 3348 5026 3352
rect 5070 3348 5074 3352
rect 5110 3348 5114 3352
rect 5134 3348 5138 3352
rect 5182 3347 5186 3351
rect 5294 3348 5298 3352
rect 2286 3338 2290 3342
rect 2350 3338 2354 3342
rect 2430 3338 2434 3342
rect 2438 3338 2442 3342
rect 2486 3338 2490 3342
rect 2494 3338 2498 3342
rect 2510 3338 2514 3342
rect 2542 3338 2546 3342
rect 2558 3338 2562 3342
rect 2574 3338 2578 3342
rect 2662 3338 2666 3342
rect 2678 3338 2682 3342
rect 2702 3338 2706 3342
rect 2734 3338 2738 3342
rect 2750 3338 2754 3342
rect 2782 3338 2786 3342
rect 2830 3338 2834 3342
rect 2902 3338 2906 3342
rect 2990 3338 2994 3342
rect 3038 3338 3042 3342
rect 3054 3338 3058 3342
rect 3094 3338 3098 3342
rect 3134 3338 3138 3342
rect 3166 3338 3170 3342
rect 3270 3338 3274 3342
rect 3310 3338 3314 3342
rect 3382 3338 3386 3342
rect 3430 3338 3434 3342
rect 3486 3338 3490 3342
rect 3566 3338 3570 3342
rect 3654 3338 3658 3342
rect 3798 3338 3802 3342
rect 3846 3338 3850 3342
rect 3854 3338 3858 3342
rect 3910 3338 3914 3342
rect 4198 3338 4202 3342
rect 4214 3338 4218 3342
rect 4262 3338 4266 3342
rect 4350 3338 4354 3342
rect 4358 3338 4362 3342
rect 4366 3338 4370 3342
rect 4398 3338 4402 3342
rect 4470 3338 4474 3342
rect 4582 3338 4586 3342
rect 4598 3338 4602 3342
rect 4622 3338 4626 3342
rect 4638 3338 4642 3342
rect 4654 3338 4658 3342
rect 4710 3338 4714 3342
rect 4854 3338 4858 3342
rect 4870 3338 4874 3342
rect 4886 3338 4890 3342
rect 4894 3338 4898 3342
rect 4966 3338 4970 3342
rect 5038 3338 5042 3342
rect 5062 3338 5066 3342
rect 5078 3338 5082 3342
rect 5094 3338 5098 3342
rect 5190 3338 5194 3342
rect 5254 3338 5258 3342
rect 5310 3338 5314 3342
rect 6 3328 10 3332
rect 54 3328 58 3332
rect 94 3328 98 3332
rect 110 3328 114 3332
rect 182 3328 186 3332
rect 214 3328 218 3332
rect 270 3328 274 3332
rect 318 3328 322 3332
rect 478 3328 482 3332
rect 510 3328 514 3332
rect 598 3328 602 3332
rect 678 3328 682 3332
rect 710 3328 714 3332
rect 750 3328 754 3332
rect 1006 3328 1010 3332
rect 1046 3328 1050 3332
rect 1118 3328 1122 3332
rect 1190 3328 1194 3332
rect 1198 3328 1202 3332
rect 1510 3328 1514 3332
rect 1590 3328 1594 3332
rect 1614 3328 1618 3332
rect 1638 3328 1642 3332
rect 1734 3328 1738 3332
rect 1774 3328 1778 3332
rect 1822 3328 1826 3332
rect 1862 3328 1866 3332
rect 2022 3328 2026 3332
rect 2158 3328 2162 3332
rect 2190 3328 2194 3332
rect 2294 3328 2298 3332
rect 2366 3328 2370 3332
rect 2494 3328 2498 3332
rect 2526 3328 2530 3332
rect 2686 3328 2690 3332
rect 2718 3328 2722 3332
rect 2774 3328 2778 3332
rect 3006 3328 3010 3332
rect 3014 3328 3018 3332
rect 3070 3328 3074 3332
rect 3118 3328 3122 3332
rect 3190 3328 3194 3332
rect 3230 3328 3234 3332
rect 3246 3328 3250 3332
rect 3262 3328 3266 3332
rect 3302 3328 3306 3332
rect 3462 3328 3466 3332
rect 3510 3328 3514 3332
rect 3910 3328 3914 3332
rect 4038 3328 4042 3332
rect 4246 3328 4250 3332
rect 4430 3328 4434 3332
rect 4622 3328 4626 3332
rect 4678 3328 4682 3332
rect 4830 3328 4834 3332
rect 4934 3328 4938 3332
rect 5006 3328 5010 3332
rect 5046 3328 5050 3332
rect 5150 3328 5154 3332
rect 22 3318 26 3322
rect 70 3318 74 3322
rect 102 3318 106 3322
rect 142 3318 146 3322
rect 206 3318 210 3322
rect 222 3318 226 3322
rect 326 3318 330 3322
rect 742 3318 746 3322
rect 830 3318 834 3322
rect 1110 3318 1114 3322
rect 1270 3318 1274 3322
rect 1286 3318 1290 3322
rect 1334 3318 1338 3322
rect 1646 3318 1650 3322
rect 1686 3318 1690 3322
rect 1742 3318 1746 3322
rect 1918 3318 1922 3322
rect 1958 3318 1962 3322
rect 1982 3318 1986 3322
rect 2038 3318 2042 3322
rect 2238 3318 2242 3322
rect 2358 3318 2362 3322
rect 2390 3318 2394 3322
rect 2454 3318 2458 3322
rect 2766 3318 2770 3322
rect 2934 3318 2938 3322
rect 2974 3318 2978 3322
rect 3094 3318 3098 3322
rect 3158 3318 3162 3322
rect 3294 3318 3298 3322
rect 3718 3318 3722 3322
rect 3910 3318 3914 3322
rect 4390 3318 4394 3322
rect 4630 3318 4634 3322
rect 4670 3318 4674 3322
rect 4686 3318 4690 3322
rect 5262 3318 5266 3322
rect 5278 3318 5282 3322
rect 6 3308 10 3312
rect 318 3308 322 3312
rect 2366 3308 2370 3312
rect 3070 3308 3074 3312
rect 5238 3308 5242 3312
rect 5310 3308 5314 3312
rect 858 3303 862 3307
rect 865 3303 869 3307
rect 1874 3303 1878 3307
rect 1881 3303 1885 3307
rect 2906 3303 2910 3307
rect 2913 3303 2917 3307
rect 3930 3303 3934 3307
rect 3937 3303 3941 3307
rect 4954 3303 4958 3307
rect 4961 3303 4965 3307
rect 414 3298 418 3302
rect 2414 3298 2418 3302
rect 2926 3298 2930 3302
rect 3038 3298 3042 3302
rect 4478 3298 4482 3302
rect 5286 3298 5290 3302
rect 14 3288 18 3292
rect 54 3288 58 3292
rect 358 3288 362 3292
rect 406 3288 410 3292
rect 454 3288 458 3292
rect 494 3288 498 3292
rect 646 3288 650 3292
rect 798 3288 802 3292
rect 822 3288 826 3292
rect 942 3288 946 3292
rect 966 3288 970 3292
rect 1038 3288 1042 3292
rect 1046 3288 1050 3292
rect 1134 3288 1138 3292
rect 1246 3288 1250 3292
rect 1262 3288 1266 3292
rect 1350 3288 1354 3292
rect 1454 3288 1458 3292
rect 1710 3288 1714 3292
rect 2038 3288 2042 3292
rect 2046 3288 2050 3292
rect 2086 3288 2090 3292
rect 2150 3288 2154 3292
rect 2166 3288 2170 3292
rect 2190 3288 2194 3292
rect 2230 3288 2234 3292
rect 2262 3288 2266 3292
rect 2430 3288 2434 3292
rect 2502 3288 2506 3292
rect 2550 3288 2554 3292
rect 2622 3288 2626 3292
rect 2646 3288 2650 3292
rect 2774 3288 2778 3292
rect 2998 3288 3002 3292
rect 3030 3288 3034 3292
rect 3174 3288 3178 3292
rect 3422 3288 3426 3292
rect 3606 3288 3610 3292
rect 3774 3288 3778 3292
rect 3846 3288 3850 3292
rect 3974 3288 3978 3292
rect 3998 3288 4002 3292
rect 4022 3288 4026 3292
rect 4046 3288 4050 3292
rect 4230 3288 4234 3292
rect 4326 3288 4330 3292
rect 4366 3288 4370 3292
rect 4494 3288 4498 3292
rect 4542 3288 4546 3292
rect 4670 3288 4674 3292
rect 4726 3288 4730 3292
rect 4838 3288 4842 3292
rect 4854 3288 4858 3292
rect 4894 3288 4898 3292
rect 4926 3288 4930 3292
rect 5054 3288 5058 3292
rect 5070 3288 5074 3292
rect 5102 3288 5106 3292
rect 5190 3288 5194 3292
rect 62 3278 66 3282
rect 134 3278 138 3282
rect 414 3278 418 3282
rect 446 3278 450 3282
rect 574 3278 578 3282
rect 726 3278 730 3282
rect 830 3278 834 3282
rect 862 3278 866 3282
rect 902 3278 906 3282
rect 990 3278 994 3282
rect 1078 3278 1082 3282
rect 1206 3278 1210 3282
rect 1254 3278 1258 3282
rect 1446 3278 1450 3282
rect 1470 3278 1474 3282
rect 1526 3278 1530 3282
rect 1686 3278 1690 3282
rect 1718 3278 1722 3282
rect 1766 3278 1770 3282
rect 1830 3278 1834 3282
rect 2054 3278 2058 3282
rect 2078 3278 2082 3282
rect 2142 3278 2146 3282
rect 2222 3278 2226 3282
rect 2270 3278 2274 3282
rect 2318 3278 2322 3282
rect 2414 3278 2418 3282
rect 2462 3278 2466 3282
rect 2478 3278 2482 3282
rect 6 3268 10 3272
rect 46 3268 50 3272
rect 110 3268 114 3272
rect 126 3268 130 3272
rect 158 3268 162 3272
rect 206 3268 210 3272
rect 14 3258 18 3262
rect 38 3258 42 3262
rect 78 3258 82 3262
rect 102 3258 106 3262
rect 118 3258 122 3262
rect 134 3258 138 3262
rect 166 3258 170 3262
rect 262 3268 266 3272
rect 318 3268 322 3272
rect 350 3268 354 3272
rect 470 3268 474 3272
rect 502 3268 506 3272
rect 550 3268 554 3272
rect 614 3268 618 3272
rect 662 3268 666 3272
rect 670 3268 674 3272
rect 734 3268 738 3272
rect 782 3268 786 3272
rect 806 3268 810 3272
rect 838 3268 842 3272
rect 886 3268 890 3272
rect 902 3268 906 3272
rect 910 3268 914 3272
rect 958 3268 962 3272
rect 982 3268 986 3272
rect 1014 3268 1018 3272
rect 1022 3268 1026 3272
rect 1150 3268 1154 3272
rect 1198 3268 1202 3272
rect 1222 3268 1226 3272
rect 1270 3268 1274 3272
rect 1286 3268 1290 3272
rect 1366 3268 1370 3272
rect 1390 3268 1394 3272
rect 1438 3268 1442 3272
rect 1446 3268 1450 3272
rect 1534 3268 1538 3272
rect 1582 3268 1586 3272
rect 1638 3268 1642 3272
rect 1646 3268 1650 3272
rect 1662 3268 1666 3272
rect 1694 3268 1698 3272
rect 1734 3268 1738 3272
rect 1838 3268 1842 3272
rect 1886 3268 1890 3272
rect 1934 3268 1938 3272
rect 1982 3268 1986 3272
rect 1990 3268 1994 3272
rect 2102 3268 2106 3272
rect 2110 3268 2114 3272
rect 2126 3268 2130 3272
rect 2222 3268 2226 3272
rect 2238 3268 2242 3272
rect 2310 3268 2314 3272
rect 2366 3268 2370 3272
rect 2382 3268 2386 3272
rect 2430 3268 2434 3272
rect 2510 3268 2514 3272
rect 2630 3278 2634 3282
rect 2726 3278 2730 3282
rect 2790 3278 2794 3282
rect 2926 3278 2930 3282
rect 3030 3278 3034 3282
rect 3062 3278 3066 3282
rect 3166 3278 3170 3282
rect 3254 3278 3258 3282
rect 3766 3278 3770 3282
rect 3830 3279 3834 3283
rect 2566 3268 2570 3272
rect 2582 3268 2586 3272
rect 2622 3268 2626 3272
rect 2670 3268 2674 3272
rect 2678 3268 2682 3272
rect 2710 3268 2714 3272
rect 2822 3268 2826 3272
rect 2862 3268 2866 3272
rect 2950 3268 2954 3272
rect 2958 3268 2962 3272
rect 270 3258 274 3262
rect 310 3258 314 3262
rect 326 3258 330 3262
rect 374 3258 378 3262
rect 390 3258 394 3262
rect 398 3258 402 3262
rect 422 3258 426 3262
rect 462 3258 466 3262
rect 558 3258 562 3262
rect 590 3258 594 3262
rect 790 3258 794 3262
rect 814 3258 818 3262
rect 878 3258 882 3262
rect 1006 3258 1010 3262
rect 1062 3258 1066 3262
rect 1094 3258 1098 3262
rect 1222 3258 1226 3262
rect 1230 3258 1234 3262
rect 1278 3258 1282 3262
rect 1294 3258 1298 3262
rect 1462 3258 1466 3262
rect 1486 3258 1490 3262
rect 1510 3258 1514 3262
rect 1542 3258 1546 3262
rect 1566 3258 1570 3262
rect 1582 3258 1586 3262
rect 1742 3258 1746 3262
rect 1750 3258 1754 3262
rect 1774 3258 1778 3262
rect 1790 3258 1794 3262
rect 1814 3258 1818 3262
rect 1838 3258 1842 3262
rect 1926 3258 1930 3262
rect 1998 3258 2002 3262
rect 2062 3258 2066 3262
rect 2118 3258 2122 3262
rect 2238 3258 2242 3262
rect 2286 3258 2290 3262
rect 2302 3258 2306 3262
rect 2326 3258 2330 3262
rect 2342 3258 2346 3262
rect 2374 3258 2378 3262
rect 2446 3258 2450 3262
rect 2534 3258 2538 3262
rect 2614 3258 2618 3262
rect 2678 3258 2682 3262
rect 2686 3258 2690 3262
rect 2710 3258 2714 3262
rect 2790 3258 2794 3262
rect 2814 3258 2818 3262
rect 2838 3258 2842 3262
rect 2870 3258 2874 3262
rect 2894 3258 2898 3262
rect 2966 3258 2970 3262
rect 3022 3258 3026 3262
rect 3054 3268 3058 3272
rect 3094 3268 3098 3272
rect 3102 3268 3106 3272
rect 3182 3268 3186 3272
rect 3078 3258 3082 3262
rect 3110 3258 3114 3262
rect 3142 3258 3146 3262
rect 3190 3258 3194 3262
rect 3214 3258 3218 3262
rect 3286 3268 3290 3272
rect 3302 3268 3306 3272
rect 3310 3268 3314 3272
rect 3358 3268 3362 3272
rect 3390 3268 3394 3272
rect 3414 3268 3418 3272
rect 3454 3268 3458 3272
rect 3486 3268 3490 3272
rect 3510 3268 3514 3272
rect 3654 3268 3658 3272
rect 3894 3268 3898 3272
rect 4262 3278 4266 3282
rect 4502 3278 4506 3282
rect 4510 3278 4514 3282
rect 4550 3278 4554 3282
rect 4558 3278 4562 3282
rect 4574 3278 4578 3282
rect 4702 3278 4706 3282
rect 4734 3278 4738 3282
rect 4758 3278 4762 3282
rect 4806 3278 4810 3282
rect 4846 3278 4850 3282
rect 4886 3278 4890 3282
rect 4958 3278 4962 3282
rect 4990 3278 4994 3282
rect 5038 3278 5042 3282
rect 4078 3268 4082 3272
rect 4246 3268 4250 3272
rect 4334 3268 4338 3272
rect 4382 3268 4386 3272
rect 3246 3258 3250 3262
rect 3294 3258 3298 3262
rect 3382 3258 3386 3262
rect 3446 3258 3450 3262
rect 3478 3258 3482 3262
rect 3494 3258 3498 3262
rect 3542 3259 3546 3263
rect 3574 3258 3578 3262
rect 3638 3259 3642 3263
rect 3710 3258 3714 3262
rect 3718 3258 3722 3262
rect 3742 3258 3746 3262
rect 3782 3258 3786 3262
rect 3838 3258 3842 3262
rect 3910 3259 3914 3263
rect 3950 3258 3954 3262
rect 4038 3258 4042 3262
rect 4110 3259 4114 3263
rect 4166 3259 4170 3263
rect 4486 3268 4490 3272
rect 4534 3268 4538 3272
rect 4606 3268 4610 3272
rect 4678 3268 4682 3272
rect 4830 3268 4834 3272
rect 4870 3266 4874 3270
rect 4886 3268 4890 3272
rect 4902 3268 4906 3272
rect 4918 3268 4922 3272
rect 4942 3268 4946 3272
rect 4982 3268 4986 3272
rect 4998 3268 5002 3272
rect 5022 3268 5026 3272
rect 5062 3268 5066 3272
rect 5086 3268 5090 3272
rect 5094 3268 5098 3272
rect 5126 3268 5130 3272
rect 4198 3258 4202 3262
rect 4270 3258 4274 3262
rect 4390 3258 4394 3262
rect 4462 3258 4466 3262
rect 4558 3258 4562 3262
rect 4614 3258 4618 3262
rect 4678 3258 4682 3262
rect 4710 3258 4714 3262
rect 4742 3258 4746 3262
rect 4774 3258 4778 3262
rect 4910 3258 4914 3262
rect 4958 3258 4962 3262
rect 5046 3258 5050 3262
rect 5102 3258 5106 3262
rect 5118 3258 5122 3262
rect 5150 3278 5154 3282
rect 5254 3279 5258 3283
rect 5286 3278 5290 3282
rect 5150 3268 5154 3272
rect 5166 3268 5170 3272
rect 5198 3268 5202 3272
rect 5206 3268 5210 3272
rect 5214 3268 5218 3272
rect 5174 3258 5178 3262
rect 5190 3258 5194 3262
rect 5238 3258 5242 3262
rect 5262 3258 5266 3262
rect 5270 3258 5274 3262
rect 30 3248 34 3252
rect 70 3248 74 3252
rect 182 3248 186 3252
rect 190 3248 194 3252
rect 494 3248 498 3252
rect 566 3248 570 3252
rect 606 3248 610 3252
rect 670 3248 674 3252
rect 790 3248 794 3252
rect 854 3248 858 3252
rect 966 3248 970 3252
rect 990 3248 994 3252
rect 1038 3248 1042 3252
rect 1046 3248 1050 3252
rect 1158 3248 1162 3252
rect 1246 3248 1250 3252
rect 1310 3248 1314 3252
rect 1566 3248 1570 3252
rect 1662 3248 1666 3252
rect 1694 3248 1698 3252
rect 1726 3248 1730 3252
rect 1758 3248 1762 3252
rect 1782 3248 1786 3252
rect 1966 3248 1970 3252
rect 1998 3248 2002 3252
rect 2022 3248 2026 3252
rect 2038 3248 2042 3252
rect 2142 3248 2146 3252
rect 2174 3248 2178 3252
rect 2214 3248 2218 3252
rect 2286 3248 2290 3252
rect 2334 3248 2338 3252
rect 2406 3248 2410 3252
rect 2502 3248 2506 3252
rect 2526 3248 2530 3252
rect 2646 3248 2650 3252
rect 2702 3248 2706 3252
rect 2750 3248 2754 3252
rect 2798 3248 2802 3252
rect 2830 3248 2834 3252
rect 2926 3248 2930 3252
rect 3070 3248 3074 3252
rect 3126 3248 3130 3252
rect 3198 3248 3202 3252
rect 3222 3248 3226 3252
rect 3246 3248 3250 3252
rect 3278 3248 3282 3252
rect 3422 3248 3426 3252
rect 3430 3248 3434 3252
rect 3462 3248 3466 3252
rect 3478 3248 3482 3252
rect 3494 3248 3498 3252
rect 4462 3248 4466 3252
rect 4934 3248 4938 3252
rect 5014 3248 5018 3252
rect 5046 3248 5050 3252
rect 5070 3248 5074 3252
rect 5158 3248 5162 3252
rect 86 3238 90 3242
rect 246 3238 250 3242
rect 358 3238 362 3242
rect 694 3238 698 3242
rect 1558 3238 1562 3242
rect 1622 3238 1626 3242
rect 1798 3238 1802 3242
rect 1870 3238 1874 3242
rect 2086 3238 2090 3242
rect 2350 3238 2354 3242
rect 2430 3238 2434 3242
rect 2846 3238 2850 3242
rect 3086 3238 3090 3242
rect 3206 3238 3210 3242
rect 3702 3238 3706 3242
rect 4422 3238 4426 3242
rect 14 3218 18 3222
rect 166 3218 170 3222
rect 1806 3218 1810 3222
rect 2302 3218 2306 3222
rect 2342 3218 2346 3222
rect 2686 3218 2690 3222
rect 2814 3218 2818 3222
rect 2854 3218 2858 3222
rect 2886 3218 2890 3222
rect 2942 3218 2946 3222
rect 3158 3218 3162 3222
rect 3254 3218 3258 3222
rect 3342 3218 3346 3222
rect 4758 3218 4762 3222
rect 4790 3218 4794 3222
rect 5278 3218 5282 3222
rect 346 3203 350 3207
rect 353 3203 357 3207
rect 1370 3203 1374 3207
rect 1377 3203 1381 3207
rect 2394 3203 2398 3207
rect 2401 3203 2405 3207
rect 3418 3203 3422 3207
rect 3425 3203 3429 3207
rect 4442 3203 4446 3207
rect 4449 3203 4453 3207
rect 206 3188 210 3192
rect 286 3188 290 3192
rect 374 3188 378 3192
rect 566 3188 570 3192
rect 734 3188 738 3192
rect 862 3188 866 3192
rect 886 3188 890 3192
rect 926 3188 930 3192
rect 1134 3188 1138 3192
rect 1142 3188 1146 3192
rect 1262 3188 1266 3192
rect 1318 3188 1322 3192
rect 1358 3188 1362 3192
rect 1422 3188 1426 3192
rect 1470 3188 1474 3192
rect 1494 3188 1498 3192
rect 1686 3188 1690 3192
rect 2438 3188 2442 3192
rect 2766 3188 2770 3192
rect 2814 3188 2818 3192
rect 2974 3188 2978 3192
rect 3174 3188 3178 3192
rect 3198 3188 3202 3192
rect 3246 3188 3250 3192
rect 3510 3188 3514 3192
rect 3550 3188 3554 3192
rect 3614 3188 3618 3192
rect 3758 3188 3762 3192
rect 3926 3188 3930 3192
rect 4038 3188 4042 3192
rect 4150 3188 4154 3192
rect 4214 3188 4218 3192
rect 4470 3188 4474 3192
rect 4606 3188 4610 3192
rect 4726 3188 4730 3192
rect 4854 3188 4858 3192
rect 478 3178 482 3182
rect 1182 3178 1186 3182
rect 4414 3178 4418 3182
rect 6 3168 10 3172
rect 30 3168 34 3172
rect 38 3168 42 3172
rect 326 3168 330 3172
rect 366 3168 370 3172
rect 454 3168 458 3172
rect 470 3168 474 3172
rect 894 3168 898 3172
rect 934 3168 938 3172
rect 958 3168 962 3172
rect 1190 3168 1194 3172
rect 1214 3168 1218 3172
rect 1270 3168 1274 3172
rect 1294 3168 1298 3172
rect 1430 3168 1434 3172
rect 1478 3168 1482 3172
rect 2662 3168 2666 3172
rect 3502 3168 3506 3172
rect 4838 3168 4842 3172
rect 5078 3168 5082 3172
rect 5246 3168 5250 3172
rect 46 3158 50 3162
rect 94 3158 98 3162
rect 110 3158 114 3162
rect 214 3158 218 3162
rect 302 3158 306 3162
rect 310 3158 314 3162
rect 382 3158 386 3162
rect 478 3158 482 3162
rect 526 3158 530 3162
rect 558 3158 562 3162
rect 910 3158 914 3162
rect 918 3158 922 3162
rect 1174 3158 1178 3162
rect 1254 3158 1258 3162
rect 1350 3158 1354 3162
rect 1406 3158 1410 3162
rect 1414 3158 1418 3162
rect 38 3148 42 3152
rect 62 3148 66 3152
rect 78 3148 82 3152
rect 102 3148 106 3152
rect 126 3148 130 3152
rect 238 3148 242 3152
rect 286 3148 290 3152
rect 374 3148 378 3152
rect 478 3148 482 3152
rect 526 3148 530 3152
rect 534 3148 538 3152
rect 774 3148 778 3152
rect 902 3148 906 3152
rect 926 3148 930 3152
rect 966 3148 970 3152
rect 982 3148 986 3152
rect 998 3148 1002 3152
rect 1166 3148 1170 3152
rect 1182 3148 1186 3152
rect 1214 3148 1218 3152
rect 1238 3148 1242 3152
rect 1262 3148 1266 3152
rect 1342 3148 1346 3152
rect 1390 3148 1394 3152
rect 1422 3148 1426 3152
rect 1462 3148 1466 3152
rect 1470 3148 1474 3152
rect 1494 3148 1498 3152
rect 1654 3158 1658 3162
rect 1718 3158 1722 3162
rect 1742 3158 1746 3162
rect 1806 3158 1810 3162
rect 2294 3158 2298 3162
rect 1550 3148 1554 3152
rect 1638 3148 1642 3152
rect 1670 3148 1674 3152
rect 1694 3148 1698 3152
rect 70 3138 74 3142
rect 118 3138 122 3142
rect 134 3138 138 3142
rect 142 3138 146 3142
rect 190 3138 194 3142
rect 214 3138 218 3142
rect 270 3138 274 3142
rect 278 3138 282 3142
rect 398 3138 402 3142
rect 422 3138 426 3142
rect 502 3138 506 3142
rect 510 3138 514 3142
rect 1766 3148 1770 3152
rect 1806 3148 1810 3152
rect 1870 3148 1874 3152
rect 1942 3148 1946 3152
rect 2094 3148 2098 3152
rect 2158 3148 2162 3152
rect 2254 3148 2258 3152
rect 2318 3158 2322 3162
rect 2398 3158 2402 3162
rect 2638 3158 2642 3162
rect 2646 3158 2650 3162
rect 2358 3148 2362 3152
rect 2494 3148 2498 3152
rect 2534 3148 2538 3152
rect 2622 3148 2626 3152
rect 2742 3158 2746 3162
rect 2838 3158 2842 3162
rect 3014 3158 3018 3162
rect 3038 3158 3042 3162
rect 3158 3158 3162 3162
rect 2654 3148 2658 3152
rect 2670 3148 2674 3152
rect 2678 3148 2682 3152
rect 2702 3148 2706 3152
rect 2750 3148 2754 3152
rect 2782 3148 2786 3152
rect 2998 3148 3002 3152
rect 3134 3148 3138 3152
rect 3174 3148 3178 3152
rect 3238 3158 3242 3162
rect 3230 3148 3234 3152
rect 3278 3148 3282 3152
rect 3294 3148 3298 3152
rect 3326 3148 3330 3152
rect 3422 3158 3426 3162
rect 3470 3158 3474 3162
rect 3534 3158 3538 3162
rect 3382 3148 3386 3152
rect 3446 3148 3450 3152
rect 3462 3148 3466 3152
rect 3486 3148 3490 3152
rect 3494 3148 3498 3152
rect 3558 3158 3562 3162
rect 3574 3158 3578 3162
rect 3606 3158 3610 3162
rect 3630 3158 3634 3162
rect 4262 3158 4266 3162
rect 5294 3158 5298 3162
rect 3582 3148 3586 3152
rect 3654 3148 3658 3152
rect 574 3138 578 3142
rect 582 3138 586 3142
rect 630 3138 634 3142
rect 638 3138 642 3142
rect 686 3138 690 3142
rect 766 3138 770 3142
rect 798 3138 802 3142
rect 846 3138 850 3142
rect 974 3138 978 3142
rect 990 3138 994 3142
rect 1006 3138 1010 3142
rect 1054 3138 1058 3142
rect 1062 3138 1066 3142
rect 1110 3138 1114 3142
rect 1158 3138 1162 3142
rect 1230 3138 1234 3142
rect 1334 3138 1338 3142
rect 1366 3138 1370 3142
rect 1374 3138 1378 3142
rect 1406 3138 1410 3142
rect 1510 3138 1514 3142
rect 1526 3138 1530 3142
rect 1534 3138 1538 3142
rect 1582 3138 1586 3142
rect 1622 3138 1626 3142
rect 1710 3138 1714 3142
rect 1734 3140 1738 3144
rect 1742 3138 1746 3142
rect 1782 3138 1786 3142
rect 3694 3147 3698 3151
rect 3726 3148 3730 3152
rect 3766 3148 3770 3152
rect 3870 3148 3874 3152
rect 3894 3148 3898 3152
rect 3942 3148 3946 3152
rect 4078 3148 4082 3152
rect 4102 3148 4106 3152
rect 4286 3148 4290 3152
rect 4350 3147 4354 3151
rect 4622 3148 4626 3152
rect 4662 3147 4666 3151
rect 4734 3148 4738 3152
rect 4798 3148 4802 3152
rect 4862 3148 4866 3152
rect 4870 3148 4874 3152
rect 4918 3148 4922 3152
rect 4942 3148 4946 3152
rect 5022 3148 5026 3152
rect 5086 3148 5090 3152
rect 5094 3148 5098 3152
rect 5126 3148 5130 3152
rect 5134 3148 5138 3152
rect 5198 3148 5202 3152
rect 5238 3148 5242 3152
rect 5262 3148 5266 3152
rect 5278 3148 5282 3152
rect 1814 3138 1818 3142
rect 1862 3138 1866 3142
rect 1910 3138 1914 3142
rect 1958 3138 1962 3142
rect 1966 3138 1970 3142
rect 2014 3138 2018 3142
rect 2022 3138 2026 3142
rect 2094 3138 2098 3142
rect 2150 3138 2154 3142
rect 2230 3138 2234 3142
rect 2318 3138 2322 3142
rect 2350 3138 2354 3142
rect 2358 3138 2362 3142
rect 2382 3138 2386 3142
rect 2390 3138 2394 3142
rect 2398 3138 2402 3142
rect 2502 3138 2506 3142
rect 2550 3138 2554 3142
rect 2558 3138 2562 3142
rect 2606 3138 2610 3142
rect 2742 3138 2746 3142
rect 2774 3138 2778 3142
rect 2822 3138 2826 3142
rect 2894 3138 2898 3142
rect 2918 3138 2922 3142
rect 2966 3138 2970 3142
rect 2990 3138 2994 3142
rect 3046 3138 3050 3142
rect 3094 3138 3098 3142
rect 3102 3138 3106 3142
rect 3150 3138 3154 3142
rect 3182 3138 3186 3142
rect 3190 3138 3194 3142
rect 3238 3138 3242 3142
rect 3302 3138 3306 3142
rect 3334 3138 3338 3142
rect 3358 3138 3362 3142
rect 3438 3138 3442 3142
rect 3518 3138 3522 3142
rect 3558 3138 3562 3142
rect 3646 3138 3650 3142
rect 3830 3138 3834 3142
rect 4014 3138 4018 3142
rect 4022 3138 4026 3142
rect 4070 3138 4074 3142
rect 4126 3138 4130 3142
rect 4134 3140 4138 3144
rect 4158 3138 4162 3142
rect 4238 3138 4242 3142
rect 4254 3138 4258 3142
rect 4270 3138 4274 3142
rect 4318 3138 4322 3142
rect 4334 3138 4338 3142
rect 4438 3138 4442 3142
rect 4494 3138 4498 3142
rect 4542 3138 4546 3142
rect 4550 3138 4554 3142
rect 4646 3138 4650 3142
rect 14 3128 18 3132
rect 54 3128 58 3132
rect 86 3128 90 3132
rect 310 3128 314 3132
rect 342 3128 346 3132
rect 414 3128 418 3132
rect 430 3128 434 3132
rect 454 3128 458 3132
rect 502 3128 506 3132
rect 710 3128 714 3132
rect 878 3128 882 3132
rect 958 3128 962 3132
rect 1118 3128 1122 3132
rect 1142 3128 1146 3132
rect 1214 3128 1218 3132
rect 1246 3128 1250 3132
rect 1278 3128 1282 3132
rect 1294 3128 1298 3132
rect 1302 3128 1306 3132
rect 1446 3128 1450 3132
rect 1510 3128 1514 3132
rect 1590 3128 1594 3132
rect 1710 3128 1714 3132
rect 1782 3128 1786 3132
rect 2078 3128 2082 3132
rect 2174 3128 2178 3132
rect 2262 3128 2266 3132
rect 2374 3128 2378 3132
rect 2478 3128 2482 3132
rect 2694 3128 2698 3132
rect 2726 3128 2730 3132
rect 2806 3128 2810 3132
rect 2982 3128 2986 3132
rect 3214 3128 3218 3132
rect 3262 3128 3266 3132
rect 3366 3128 3370 3132
rect 3406 3128 3410 3132
rect 3470 3128 3474 3132
rect 3598 3128 3602 3132
rect 4774 3138 4778 3142
rect 4950 3138 4954 3142
rect 5030 3138 5034 3142
rect 5214 3138 5218 3142
rect 5270 3138 5274 3142
rect 4086 3127 4090 3131
rect 4110 3127 4114 3131
rect 4622 3128 4626 3132
rect 4694 3128 4698 3132
rect 4918 3128 4922 3132
rect 4942 3128 4946 3132
rect 5142 3128 5146 3132
rect 174 3118 178 3122
rect 406 3118 410 3122
rect 614 3118 618 3122
rect 830 3118 834 3122
rect 1038 3118 1042 3122
rect 1046 3118 1050 3122
rect 1094 3118 1098 3122
rect 1262 3118 1266 3122
rect 1582 3118 1586 3122
rect 1750 3118 1754 3122
rect 1822 3118 1826 3122
rect 1830 3118 1834 3122
rect 1998 3118 2002 3122
rect 2038 3118 2042 3122
rect 2086 3118 2090 3122
rect 2094 3118 2098 3122
rect 2118 3118 2122 3122
rect 2214 3118 2218 3122
rect 2302 3118 2306 3122
rect 2702 3118 2706 3122
rect 2798 3118 2802 3122
rect 2862 3118 2866 3122
rect 2950 3118 2954 3122
rect 3038 3118 3042 3122
rect 3070 3118 3074 3122
rect 3142 3118 3146 3122
rect 3174 3118 3178 3122
rect 3294 3118 3298 3122
rect 3310 3118 3314 3122
rect 3342 3118 3346 3122
rect 4230 3118 4234 3122
rect 4510 3118 4514 3122
rect 4606 3118 4610 3122
rect 4750 3118 4754 3122
rect 4950 3118 4954 3122
rect 5182 3118 5186 3122
rect 5302 3118 5306 3122
rect 1142 3108 1146 3112
rect 1710 3108 1714 3112
rect 2598 3108 2602 3112
rect 2694 3108 2698 3112
rect 3214 3108 3218 3112
rect 4238 3108 4242 3112
rect 4870 3108 4874 3112
rect 4942 3108 4946 3112
rect 858 3103 862 3107
rect 865 3103 869 3107
rect 1874 3103 1878 3107
rect 1881 3103 1885 3107
rect 2906 3103 2910 3107
rect 2913 3103 2917 3107
rect 3930 3103 3934 3107
rect 3937 3103 3941 3107
rect 4954 3103 4958 3107
rect 4961 3103 4965 3107
rect 510 3098 514 3102
rect 846 3098 850 3102
rect 1174 3098 1178 3102
rect 1454 3098 1458 3102
rect 1854 3098 1858 3102
rect 2022 3098 2026 3102
rect 2590 3098 2594 3102
rect 2606 3098 2610 3102
rect 2990 3098 2994 3102
rect 3286 3098 3290 3102
rect 4494 3098 4498 3102
rect 4694 3098 4698 3102
rect 5238 3098 5242 3102
rect 62 3088 66 3092
rect 150 3088 154 3092
rect 190 3088 194 3092
rect 262 3088 266 3092
rect 310 3088 314 3092
rect 334 3088 338 3092
rect 414 3088 418 3092
rect 470 3088 474 3092
rect 478 3088 482 3092
rect 542 3088 546 3092
rect 574 3088 578 3092
rect 670 3088 674 3092
rect 718 3088 722 3092
rect 878 3088 882 3092
rect 894 3088 898 3092
rect 942 3088 946 3092
rect 1006 3088 1010 3092
rect 1078 3088 1082 3092
rect 1110 3088 1114 3092
rect 1126 3088 1130 3092
rect 1214 3088 1218 3092
rect 1350 3088 1354 3092
rect 1398 3088 1402 3092
rect 1510 3088 1514 3092
rect 1534 3088 1538 3092
rect 1590 3088 1594 3092
rect 1646 3088 1650 3092
rect 1662 3088 1666 3092
rect 1758 3088 1762 3092
rect 1982 3088 1986 3092
rect 2446 3088 2450 3092
rect 2486 3088 2490 3092
rect 2574 3088 2578 3092
rect 2654 3088 2658 3092
rect 2718 3088 2722 3092
rect 2742 3088 2746 3092
rect 2894 3088 2898 3092
rect 3222 3088 3226 3092
rect 3262 3088 3266 3092
rect 3278 3088 3282 3092
rect 3822 3088 3826 3092
rect 3878 3088 3882 3092
rect 3990 3088 3994 3092
rect 4070 3088 4074 3092
rect 4222 3088 4226 3092
rect 4270 3088 4274 3092
rect 4398 3088 4402 3092
rect 4462 3088 4466 3092
rect 4574 3088 4578 3092
rect 4686 3088 4690 3092
rect 4742 3088 4746 3092
rect 4790 3088 4794 3092
rect 4830 3088 4834 3092
rect 4854 3088 4858 3092
rect 4910 3088 4914 3092
rect 5150 3088 5154 3092
rect 5246 3088 5250 3092
rect 14 3079 18 3083
rect 54 3078 58 3082
rect 198 3078 202 3082
rect 286 3078 290 3082
rect 422 3078 426 3082
rect 510 3078 514 3082
rect 70 3068 74 3072
rect 158 3068 162 3072
rect 174 3068 178 3072
rect 254 3068 258 3072
rect 270 3068 274 3072
rect 294 3068 298 3072
rect 302 3068 306 3072
rect 350 3068 354 3072
rect 398 3068 402 3072
rect 446 3068 450 3072
rect 534 3068 538 3072
rect 550 3068 554 3072
rect 558 3068 562 3072
rect 606 3068 610 3072
rect 614 3068 618 3072
rect 670 3068 674 3072
rect 686 3068 690 3072
rect 694 3068 698 3072
rect 742 3068 746 3072
rect 838 3078 842 3082
rect 846 3078 850 3082
rect 950 3078 954 3082
rect 1038 3078 1042 3082
rect 1134 3078 1138 3082
rect 1174 3078 1178 3082
rect 1302 3078 1306 3082
rect 1358 3078 1362 3082
rect 1454 3078 1458 3082
rect 1854 3078 1858 3082
rect 2022 3078 2026 3082
rect 2230 3078 2234 3082
rect 2374 3078 2378 3082
rect 2382 3078 2386 3082
rect 2590 3078 2594 3082
rect 2678 3078 2682 3082
rect 2830 3078 2834 3082
rect 3006 3078 3010 3082
rect 3062 3078 3066 3082
rect 3286 3078 3290 3082
rect 3294 3078 3298 3082
rect 3350 3078 3354 3082
rect 3366 3078 3370 3082
rect 3454 3078 3458 3082
rect 3462 3078 3466 3082
rect 3534 3078 3538 3082
rect 3582 3078 3586 3082
rect 3646 3078 3650 3082
rect 774 3068 778 3072
rect 790 3068 794 3072
rect 806 3068 810 3072
rect 822 3068 826 3072
rect 910 3068 914 3072
rect 918 3068 922 3072
rect 966 3068 970 3072
rect 1038 3068 1042 3072
rect 1118 3068 1122 3072
rect 1142 3068 1146 3072
rect 1174 3068 1178 3072
rect 1262 3068 1266 3072
rect 1302 3068 1306 3072
rect 1382 3068 1386 3072
rect 1406 3068 1410 3072
rect 1422 3068 1426 3072
rect 1462 3068 1466 3072
rect 1478 3068 1482 3072
rect 22 3058 26 3062
rect 78 3058 82 3062
rect 94 3058 98 3062
rect 174 3058 178 3062
rect 230 3058 234 3062
rect 246 3058 250 3062
rect 278 3058 282 3062
rect 398 3058 402 3062
rect 422 3058 426 3062
rect 438 3058 442 3062
rect 454 3058 458 3062
rect 494 3058 498 3062
rect 526 3058 530 3062
rect 662 3058 666 3062
rect 750 3058 754 3062
rect 782 3058 786 3062
rect 814 3058 818 3062
rect 926 3058 930 3062
rect 966 3058 970 3062
rect 974 3058 978 3062
rect 990 3058 994 3062
rect 1014 3058 1018 3062
rect 1494 3066 1498 3070
rect 1550 3068 1554 3072
rect 1598 3068 1602 3072
rect 1726 3068 1730 3072
rect 1902 3068 1906 3072
rect 1990 3068 1994 3072
rect 2094 3068 2098 3072
rect 2126 3068 2130 3072
rect 2182 3068 2186 3072
rect 2270 3068 2274 3072
rect 2318 3068 2322 3072
rect 2326 3068 2330 3072
rect 2350 3068 2354 3072
rect 2454 3068 2458 3072
rect 2510 3068 2514 3072
rect 2518 3068 2522 3072
rect 2574 3068 2578 3072
rect 2598 3068 2602 3072
rect 2694 3068 2698 3072
rect 2726 3068 2730 3072
rect 2774 3068 2778 3072
rect 2854 3068 2858 3072
rect 2902 3068 2906 3072
rect 2950 3068 2954 3072
rect 2958 3068 2962 3072
rect 2974 3068 2978 3072
rect 3014 3068 3018 3072
rect 3078 3068 3082 3072
rect 3126 3068 3130 3072
rect 3158 3068 3162 3072
rect 3206 3068 3210 3072
rect 3214 3068 3218 3072
rect 3318 3068 3322 3072
rect 3366 3068 3370 3072
rect 3502 3068 3506 3072
rect 3518 3068 3522 3072
rect 3534 3068 3538 3072
rect 3630 3068 3634 3072
rect 4038 3078 4042 3082
rect 4166 3078 4170 3082
rect 4182 3078 4186 3082
rect 4366 3078 4370 3082
rect 4510 3078 4514 3082
rect 3686 3068 3690 3072
rect 3710 3068 3714 3072
rect 3726 3068 3730 3072
rect 3782 3068 3786 3072
rect 3790 3068 3794 3072
rect 3838 3068 3842 3072
rect 3846 3068 3850 3072
rect 3894 3068 3898 3072
rect 3902 3068 3906 3072
rect 3950 3068 3954 3072
rect 4006 3068 4010 3072
rect 1062 3058 1066 3062
rect 1094 3058 1098 3062
rect 1110 3058 1114 3062
rect 1150 3058 1154 3062
rect 1190 3058 1194 3062
rect 1214 3058 1218 3062
rect 1238 3058 1242 3062
rect 1270 3058 1274 3062
rect 1286 3058 1290 3062
rect 1326 3058 1330 3062
rect 1414 3058 1418 3062
rect 1438 3058 1442 3062
rect 1534 3058 1538 3062
rect 1614 3058 1618 3062
rect 1718 3058 1722 3062
rect 1790 3058 1794 3062
rect 1822 3059 1826 3063
rect 1870 3058 1874 3062
rect 1918 3059 1922 3063
rect 2046 3058 2050 3062
rect 2102 3058 2106 3062
rect 2246 3058 2250 3062
rect 2334 3058 2338 3062
rect 2358 3058 2362 3062
rect 2574 3058 2578 3062
rect 2606 3058 2610 3062
rect 2702 3058 2706 3062
rect 2750 3058 2754 3062
rect 2846 3058 2850 3062
rect 2862 3058 2866 3062
rect 2966 3058 2970 3062
rect 2982 3058 2986 3062
rect 3094 3058 3098 3062
rect 3134 3058 3138 3062
rect 3222 3058 3226 3062
rect 3270 3058 3274 3062
rect 3310 3058 3314 3062
rect 3326 3058 3330 3062
rect 3398 3058 3402 3062
rect 3438 3058 3442 3062
rect 3494 3058 3498 3062
rect 3502 3058 3506 3062
rect 4014 3066 4018 3070
rect 4126 3068 4130 3072
rect 4142 3068 4146 3072
rect 4166 3068 4170 3072
rect 4190 3068 4194 3072
rect 4238 3068 4242 3072
rect 4246 3068 4250 3072
rect 4294 3068 4298 3072
rect 4334 3068 4338 3072
rect 4438 3068 4442 3072
rect 4486 3068 4490 3072
rect 4694 3078 4698 3082
rect 4846 3078 4850 3082
rect 5038 3078 5042 3082
rect 4526 3068 4530 3072
rect 4542 3068 4546 3072
rect 4590 3068 4594 3072
rect 4606 3068 4610 3072
rect 4646 3068 4650 3072
rect 4710 3068 4714 3072
rect 4742 3068 4746 3072
rect 4830 3068 4834 3072
rect 4854 3068 4858 3072
rect 4942 3068 4946 3072
rect 4990 3068 4994 3072
rect 5022 3068 5026 3072
rect 5038 3068 5042 3072
rect 5070 3068 5074 3072
rect 5270 3068 5274 3072
rect 3558 3058 3562 3062
rect 3606 3058 3610 3062
rect 3622 3058 3626 3062
rect 3670 3058 3674 3062
rect 3694 3058 3698 3062
rect 3750 3058 3754 3062
rect 3918 3058 3922 3062
rect 3974 3058 3978 3062
rect 4030 3058 4034 3062
rect 4062 3058 4066 3062
rect 4094 3058 4098 3062
rect 4150 3058 4154 3062
rect 4318 3058 4322 3062
rect 4342 3058 4346 3062
rect 4366 3058 4370 3062
rect 4390 3058 4394 3062
rect 4406 3058 4410 3062
rect 4414 3058 4418 3062
rect 4430 3058 4434 3062
rect 4478 3058 4482 3062
rect 4494 3058 4498 3062
rect 4534 3058 4538 3062
rect 4622 3059 4626 3063
rect 4726 3058 4730 3062
rect 4830 3058 4834 3062
rect 4846 3058 4850 3062
rect 4950 3058 4954 3062
rect 4958 3058 4962 3062
rect 5006 3058 5010 3062
rect 5030 3058 5034 3062
rect 5086 3059 5090 3063
rect 5182 3059 5186 3063
rect 5206 3058 5210 3062
rect 5254 3058 5258 3062
rect 5286 3058 5290 3062
rect 86 3048 90 3052
rect 134 3048 138 3052
rect 190 3048 194 3052
rect 214 3048 218 3052
rect 238 3048 242 3052
rect 414 3048 418 3052
rect 470 3048 474 3052
rect 534 3048 538 3052
rect 670 3048 674 3052
rect 798 3048 802 3052
rect 830 3048 834 3052
rect 886 3048 890 3052
rect 990 3048 994 3052
rect 1070 3048 1074 3052
rect 1102 3048 1106 3052
rect 1166 3048 1170 3052
rect 1222 3048 1226 3052
rect 1238 3048 1242 3052
rect 1254 3048 1258 3052
rect 1310 3048 1314 3052
rect 1326 3048 1330 3052
rect 1398 3048 1402 3052
rect 1446 3048 1450 3052
rect 1478 3048 1482 3052
rect 1542 3048 1546 3052
rect 1630 3048 1634 3052
rect 1654 3048 1658 3052
rect 2006 3048 2010 3052
rect 2054 3048 2058 3052
rect 2062 3048 2066 3052
rect 2102 3048 2106 3052
rect 2158 3048 2162 3052
rect 2198 3048 2202 3052
rect 2222 3048 2226 3052
rect 2350 3048 2354 3052
rect 2366 3048 2370 3052
rect 2430 3048 2434 3052
rect 2582 3048 2586 3052
rect 2622 3048 2626 3052
rect 2654 3048 2658 3052
rect 2694 3048 2698 3052
rect 2742 3048 2746 3052
rect 2982 3048 2986 3052
rect 2998 3048 3002 3052
rect 3038 3048 3042 3052
rect 3190 3048 3194 3052
rect 3238 3048 3242 3052
rect 3262 3048 3266 3052
rect 3366 3048 3370 3052
rect 3406 3048 3410 3052
rect 3430 3048 3434 3052
rect 3462 3048 3466 3052
rect 3494 3048 3498 3052
rect 3550 3048 3554 3052
rect 3566 3048 3570 3052
rect 3614 3048 3618 3052
rect 3678 3048 3682 3052
rect 3710 3048 3714 3052
rect 4038 3048 4042 3052
rect 4054 3048 4058 3052
rect 4086 3048 4090 3052
rect 4118 3048 4122 3052
rect 4326 3048 4330 3052
rect 4814 3048 4818 3052
rect 4870 3048 4874 3052
rect 5278 3048 5282 3052
rect 94 3038 98 3042
rect 222 3038 226 3042
rect 758 3038 762 3042
rect 942 3038 946 3042
rect 1006 3038 1010 3042
rect 1054 3038 1058 3042
rect 1086 3038 1090 3042
rect 1190 3038 1194 3042
rect 1214 3038 1218 3042
rect 1430 3038 1434 3042
rect 1470 3038 1474 3042
rect 1526 3038 1530 3042
rect 2038 3038 2042 3042
rect 2254 3038 2258 3042
rect 2806 3038 2810 3042
rect 3350 3038 3354 3042
rect 3390 3038 3394 3042
rect 3446 3038 3450 3042
rect 3598 3038 3602 3042
rect 3670 3038 3674 3042
rect 4070 3038 4074 3042
rect 4102 3038 4106 3042
rect 4150 3038 4154 3042
rect 4334 3038 4338 3042
rect 5294 3038 5298 3042
rect 206 3028 210 3032
rect 1062 3028 1066 3032
rect 1998 3028 2002 3032
rect 3398 3028 3402 3032
rect 1862 3018 1866 3022
rect 2014 3018 2018 3022
rect 2030 3018 2034 3022
rect 2078 3018 2082 3022
rect 2150 3018 2154 3022
rect 2214 3018 2218 3022
rect 2238 3018 2242 3022
rect 2286 3018 2290 3022
rect 2638 3018 2642 3022
rect 2934 3018 2938 3022
rect 3022 3018 3026 3022
rect 3302 3018 3306 3022
rect 3326 3018 3330 3022
rect 3558 3018 3562 3022
rect 3606 3018 3610 3022
rect 3718 3018 3722 3022
rect 4094 3018 4098 3022
rect 4302 3018 4306 3022
rect 5286 3018 5290 3022
rect 346 3003 350 3007
rect 353 3003 357 3007
rect 1370 3003 1374 3007
rect 1377 3003 1381 3007
rect 2394 3003 2398 3007
rect 2401 3003 2405 3007
rect 3418 3003 3422 3007
rect 3425 3003 3429 3007
rect 4442 3003 4446 3007
rect 4449 3003 4453 3007
rect 46 2988 50 2992
rect 94 2988 98 2992
rect 238 2988 242 2992
rect 406 2988 410 2992
rect 438 2988 442 2992
rect 510 2988 514 2992
rect 550 2988 554 2992
rect 574 2988 578 2992
rect 598 2988 602 2992
rect 702 2988 706 2992
rect 790 2988 794 2992
rect 902 2988 906 2992
rect 1006 2988 1010 2992
rect 1014 2988 1018 2992
rect 1118 2988 1122 2992
rect 1214 2988 1218 2992
rect 1230 2988 1234 2992
rect 1462 2988 1466 2992
rect 1470 2988 1474 2992
rect 1582 2988 1586 2992
rect 2414 2988 2418 2992
rect 2710 2988 2714 2992
rect 2750 2988 2754 2992
rect 2838 2988 2842 2992
rect 2878 2988 2882 2992
rect 2974 2988 2978 2992
rect 3118 2988 3122 2992
rect 3206 2988 3210 2992
rect 3726 2988 3730 2992
rect 3838 2988 3842 2992
rect 3870 2988 3874 2992
rect 4110 2988 4114 2992
rect 4158 2988 4162 2992
rect 4182 2988 4186 2992
rect 4278 2988 4282 2992
rect 4382 2988 4386 2992
rect 4846 2988 4850 2992
rect 742 2978 746 2982
rect 2118 2978 2122 2982
rect 3310 2978 3314 2982
rect 3502 2978 3506 2982
rect 54 2968 58 2972
rect 246 2968 250 2972
rect 270 2968 274 2972
rect 766 2968 770 2972
rect 1166 2968 1170 2972
rect 1342 2968 1346 2972
rect 1790 2968 1794 2972
rect 2014 2968 2018 2972
rect 2086 2968 2090 2972
rect 2150 2968 2154 2972
rect 2270 2968 2274 2972
rect 2286 2968 2290 2972
rect 2566 2968 2570 2972
rect 2686 2968 2690 2972
rect 2758 2968 2762 2972
rect 2886 2968 2890 2972
rect 3230 2968 3234 2972
rect 3358 2968 3362 2972
rect 3518 2968 3522 2972
rect 3526 2968 3530 2972
rect 3702 2968 3706 2972
rect 3766 2968 3770 2972
rect 4502 2968 4506 2972
rect 5054 2968 5058 2972
rect 70 2958 74 2962
rect 94 2958 98 2962
rect 102 2958 106 2962
rect 126 2958 130 2962
rect 158 2958 162 2962
rect 166 2958 170 2962
rect 190 2958 194 2962
rect 230 2958 234 2962
rect 262 2958 266 2962
rect 286 2958 290 2962
rect 382 2958 386 2962
rect 422 2958 426 2962
rect 6 2948 10 2952
rect 46 2948 50 2952
rect 94 2948 98 2952
rect 118 2948 122 2952
rect 142 2948 146 2952
rect 190 2948 194 2952
rect 206 2948 210 2952
rect 238 2948 242 2952
rect 278 2948 282 2952
rect 326 2948 330 2952
rect 342 2948 346 2952
rect 390 2948 394 2952
rect 454 2958 458 2962
rect 590 2958 594 2962
rect 694 2958 698 2962
rect 782 2958 786 2962
rect 1134 2958 1138 2962
rect 1198 2958 1202 2962
rect 1574 2958 1578 2962
rect 1806 2958 1810 2962
rect 1814 2958 1818 2962
rect 1846 2958 1850 2962
rect 1862 2958 1866 2962
rect 1942 2958 1946 2962
rect 1950 2958 1954 2962
rect 2030 2958 2034 2962
rect 2102 2958 2106 2962
rect 2134 2958 2138 2962
rect 2166 2958 2170 2962
rect 2230 2958 2234 2962
rect 2254 2958 2258 2962
rect 574 2948 578 2952
rect 662 2947 666 2951
rect 718 2948 722 2952
rect 734 2948 738 2952
rect 766 2948 770 2952
rect 854 2947 858 2951
rect 966 2947 970 2951
rect 1078 2947 1082 2951
rect 1118 2948 1122 2952
rect 1142 2948 1146 2952
rect 1206 2948 1210 2952
rect 1294 2947 1298 2951
rect 1406 2947 1410 2951
rect 1502 2948 1506 2952
rect 1510 2948 1514 2952
rect 1614 2948 1618 2952
rect 1646 2947 1650 2951
rect 1710 2948 1714 2952
rect 1726 2948 1730 2952
rect 1838 2948 1842 2952
rect 1902 2948 1906 2952
rect 1926 2948 1930 2952
rect 1950 2948 1954 2952
rect 1974 2948 1978 2952
rect 2006 2948 2010 2952
rect 2022 2948 2026 2952
rect 2038 2948 2042 2952
rect 2070 2948 2074 2952
rect 2078 2948 2082 2952
rect 2158 2948 2162 2952
rect 2214 2948 2218 2952
rect 2302 2958 2306 2962
rect 2510 2958 2514 2962
rect 2590 2958 2594 2962
rect 2694 2958 2698 2962
rect 2742 2958 2746 2962
rect 3086 2958 3090 2962
rect 3126 2958 3130 2962
rect 3166 2958 3170 2962
rect 3222 2958 3226 2962
rect 3278 2958 3282 2962
rect 3302 2958 3306 2962
rect 3326 2958 3330 2962
rect 3342 2958 3346 2962
rect 3374 2958 3378 2962
rect 3406 2958 3410 2962
rect 3430 2958 3434 2962
rect 3534 2958 3538 2962
rect 3582 2958 3586 2962
rect 3630 2958 3634 2962
rect 3686 2958 3690 2962
rect 3734 2958 3738 2962
rect 3798 2958 3802 2962
rect 3910 2958 3914 2962
rect 4438 2958 4442 2962
rect 4494 2958 4498 2962
rect 4542 2958 4546 2962
rect 4902 2958 4906 2962
rect 5166 2958 5170 2962
rect 2318 2948 2322 2952
rect 150 2938 154 2942
rect 198 2938 202 2942
rect 278 2938 282 2942
rect 398 2938 402 2942
rect 430 2938 434 2942
rect 494 2938 498 2942
rect 542 2938 546 2942
rect 566 2938 570 2942
rect 630 2938 634 2942
rect 694 2938 698 2942
rect 710 2938 714 2942
rect 758 2938 762 2942
rect 822 2938 826 2942
rect 870 2938 874 2942
rect 982 2938 986 2942
rect 1110 2938 1114 2942
rect 1158 2938 1162 2942
rect 1222 2938 1226 2942
rect 1286 2938 1290 2942
rect 1390 2938 1394 2942
rect 1550 2938 1554 2942
rect 1822 2938 1826 2942
rect 1838 2938 1842 2942
rect 1862 2938 1866 2942
rect 1894 2938 1898 2942
rect 1910 2938 1914 2942
rect 1918 2938 1922 2942
rect 1982 2938 1986 2942
rect 2038 2938 2042 2942
rect 2062 2938 2066 2942
rect 2070 2938 2074 2942
rect 2182 2938 2186 2942
rect 2238 2938 2242 2942
rect 2286 2938 2290 2942
rect 2310 2938 2314 2942
rect 2478 2947 2482 2951
rect 2526 2948 2530 2952
rect 2614 2948 2618 2952
rect 2622 2948 2626 2952
rect 2630 2948 2634 2952
rect 2710 2948 2714 2952
rect 2734 2948 2738 2952
rect 2750 2948 2754 2952
rect 2798 2948 2802 2952
rect 2854 2948 2858 2952
rect 2862 2948 2866 2952
rect 2878 2948 2882 2952
rect 2934 2948 2938 2952
rect 3070 2948 3074 2952
rect 3102 2948 3106 2952
rect 3150 2948 3154 2952
rect 3190 2948 3194 2952
rect 2390 2938 2394 2942
rect 2494 2938 2498 2942
rect 2526 2938 2530 2942
rect 2582 2938 2586 2942
rect 2606 2938 2610 2942
rect 2654 2938 2658 2942
rect 2670 2938 2674 2942
rect 2718 2938 2722 2942
rect 2774 2938 2778 2942
rect 2790 2938 2794 2942
rect 2846 2938 2850 2942
rect 2942 2938 2946 2942
rect 3006 2938 3010 2942
rect 3038 2938 3042 2942
rect 3062 2938 3066 2942
rect 3134 2938 3138 2942
rect 3142 2938 3146 2942
rect 3238 2948 3242 2952
rect 3262 2948 3266 2952
rect 3366 2948 3370 2952
rect 3390 2948 3394 2952
rect 3422 2948 3426 2952
rect 3454 2948 3458 2952
rect 3526 2948 3530 2952
rect 3542 2948 3546 2952
rect 3574 2948 3578 2952
rect 3598 2948 3602 2952
rect 3606 2948 3610 2952
rect 3638 2948 3642 2952
rect 3678 2948 3682 2952
rect 3694 2948 3698 2952
rect 3742 2948 3746 2952
rect 3774 2948 3778 2952
rect 3806 2948 3810 2952
rect 3830 2948 3834 2952
rect 3958 2948 3962 2952
rect 4006 2948 4010 2952
rect 4086 2948 4090 2952
rect 4166 2948 4170 2952
rect 4222 2948 4226 2952
rect 4302 2948 4306 2952
rect 4326 2948 4330 2952
rect 4470 2948 4474 2952
rect 4526 2948 4530 2952
rect 4574 2948 4578 2952
rect 4614 2948 4618 2952
rect 4710 2948 4714 2952
rect 4734 2948 4738 2952
rect 4750 2948 4754 2952
rect 3254 2938 3258 2942
rect 3286 2938 3290 2942
rect 3302 2938 3306 2942
rect 3342 2938 3346 2942
rect 3358 2938 3362 2942
rect 3382 2938 3386 2942
rect 3446 2938 3450 2942
rect 3470 2938 3474 2942
rect 3494 2938 3498 2942
rect 3542 2938 3546 2942
rect 3566 2938 3570 2942
rect 3590 2938 3594 2942
rect 3606 2938 3610 2942
rect 4782 2947 4786 2951
rect 4886 2948 4890 2952
rect 4942 2948 4946 2952
rect 4950 2948 4954 2952
rect 4990 2948 4994 2952
rect 4998 2948 5002 2952
rect 5038 2948 5042 2952
rect 5062 2948 5066 2952
rect 5070 2948 5074 2952
rect 5126 2948 5130 2952
rect 5134 2948 5138 2952
rect 5198 2947 5202 2951
rect 5294 2948 5298 2952
rect 3630 2938 3634 2942
rect 3654 2938 3658 2942
rect 3670 2938 3674 2942
rect 3718 2938 3722 2942
rect 3750 2938 3754 2942
rect 3822 2938 3826 2942
rect 3854 2938 3858 2942
rect 3902 2938 3906 2942
rect 3966 2938 3970 2942
rect 3982 2938 3986 2942
rect 4038 2938 4042 2942
rect 4086 2938 4090 2942
rect 4134 2938 4138 2942
rect 4158 2938 4162 2942
rect 4214 2938 4218 2942
rect 4246 2938 4250 2942
rect 4294 2938 4298 2942
rect 4350 2938 4354 2942
rect 4406 2938 4410 2942
rect 4414 2940 4418 2944
rect 4454 2938 4458 2942
rect 4478 2938 4482 2942
rect 4518 2938 4522 2942
rect 4566 2938 4570 2942
rect 4638 2938 4642 2942
rect 4702 2938 4706 2942
rect 4766 2938 4770 2942
rect 4870 2940 4874 2944
rect 4886 2938 4890 2942
rect 4950 2938 4954 2942
rect 5182 2938 5186 2942
rect 5206 2938 5210 2942
rect 5286 2938 5290 2942
rect 14 2927 18 2931
rect 70 2928 74 2932
rect 118 2928 122 2932
rect 166 2928 170 2932
rect 310 2928 314 2932
rect 374 2928 378 2932
rect 486 2928 490 2932
rect 558 2928 562 2932
rect 718 2928 722 2932
rect 750 2928 754 2932
rect 934 2928 938 2932
rect 998 2928 1002 2932
rect 1078 2928 1082 2932
rect 1158 2928 1162 2932
rect 1166 2928 1170 2932
rect 1438 2928 1442 2932
rect 1446 2928 1450 2932
rect 1454 2928 1458 2932
rect 1574 2928 1578 2932
rect 1774 2928 1778 2932
rect 1990 2928 1994 2932
rect 1998 2928 2002 2932
rect 2046 2928 2050 2932
rect 2110 2928 2114 2932
rect 2134 2928 2138 2932
rect 2198 2928 2202 2932
rect 2238 2928 2242 2932
rect 2598 2928 2602 2932
rect 2646 2928 2650 2932
rect 2686 2928 2690 2932
rect 2726 2928 2730 2932
rect 2774 2928 2778 2932
rect 2806 2928 2810 2932
rect 2854 2928 2858 2932
rect 3046 2928 3050 2932
rect 3214 2928 3218 2932
rect 3318 2928 3322 2932
rect 3486 2928 3490 2932
rect 3638 2928 3642 2932
rect 3654 2928 3658 2932
rect 3766 2928 3770 2932
rect 3782 2927 3786 2931
rect 3846 2928 3850 2932
rect 3974 2928 3978 2932
rect 4046 2928 4050 2932
rect 4078 2928 4082 2932
rect 4142 2928 4146 2932
rect 4454 2928 4458 2932
rect 4502 2928 4506 2932
rect 4550 2928 4554 2932
rect 4726 2928 4730 2932
rect 4974 2928 4978 2932
rect 5006 2928 5010 2932
rect 5118 2928 5122 2932
rect 5270 2928 5274 2932
rect 574 2918 578 2922
rect 1798 2918 1802 2922
rect 1830 2918 1834 2922
rect 1846 2918 1850 2922
rect 1950 2918 1954 2922
rect 2158 2918 2162 2922
rect 2302 2918 2306 2922
rect 2358 2918 2362 2922
rect 3038 2918 3042 2922
rect 3246 2918 3250 2922
rect 3278 2918 3282 2922
rect 3438 2918 3442 2922
rect 3462 2918 3466 2922
rect 3566 2918 3570 2922
rect 3710 2918 3714 2922
rect 4158 2918 4162 2922
rect 4478 2918 4482 2922
rect 4494 2918 4498 2922
rect 4542 2918 4546 2922
rect 4590 2918 4594 2922
rect 4710 2918 4714 2922
rect 4854 2918 4858 2922
rect 4886 2918 4890 2922
rect 4910 2918 4914 2922
rect 4950 2918 4954 2922
rect 5262 2918 5266 2922
rect 5278 2918 5282 2922
rect 502 2908 506 2912
rect 1158 2908 1162 2912
rect 4726 2908 4730 2912
rect 858 2903 862 2907
rect 865 2903 869 2907
rect 1874 2903 1878 2907
rect 1881 2903 1885 2907
rect 2906 2903 2910 2907
rect 2913 2903 2917 2907
rect 3930 2903 3934 2907
rect 3937 2903 3941 2907
rect 4954 2903 4958 2907
rect 4961 2903 4965 2907
rect 1110 2898 1114 2902
rect 1526 2898 1530 2902
rect 1910 2898 1914 2902
rect 4414 2898 4418 2902
rect 4550 2898 4554 2902
rect 4878 2898 4882 2902
rect 5070 2898 5074 2902
rect 14 2888 18 2892
rect 22 2888 26 2892
rect 150 2888 154 2892
rect 198 2888 202 2892
rect 310 2888 314 2892
rect 390 2888 394 2892
rect 406 2888 410 2892
rect 478 2888 482 2892
rect 510 2888 514 2892
rect 702 2888 706 2892
rect 758 2888 762 2892
rect 838 2888 842 2892
rect 934 2888 938 2892
rect 1038 2888 1042 2892
rect 1102 2888 1106 2892
rect 1198 2888 1202 2892
rect 1222 2888 1226 2892
rect 1406 2888 1410 2892
rect 1510 2888 1514 2892
rect 1542 2888 1546 2892
rect 1606 2888 1610 2892
rect 1862 2888 1866 2892
rect 2006 2888 2010 2892
rect 2142 2888 2146 2892
rect 2254 2888 2258 2892
rect 2422 2888 2426 2892
rect 2462 2888 2466 2892
rect 2558 2888 2562 2892
rect 2702 2888 2706 2892
rect 2854 2888 2858 2892
rect 3054 2888 3058 2892
rect 3086 2888 3090 2892
rect 3126 2888 3130 2892
rect 3262 2888 3266 2892
rect 3278 2888 3282 2892
rect 3326 2888 3330 2892
rect 3406 2888 3410 2892
rect 3462 2888 3466 2892
rect 3494 2888 3498 2892
rect 3574 2888 3578 2892
rect 3654 2888 3658 2892
rect 3742 2888 3746 2892
rect 3982 2888 3986 2892
rect 4054 2888 4058 2892
rect 4222 2888 4226 2892
rect 4326 2888 4330 2892
rect 4438 2888 4442 2892
rect 4454 2888 4458 2892
rect 4470 2888 4474 2892
rect 4614 2888 4618 2892
rect 5078 2888 5082 2892
rect 5174 2888 5178 2892
rect 142 2878 146 2882
rect 398 2878 402 2882
rect 678 2878 682 2882
rect 1254 2878 1258 2882
rect 1286 2878 1290 2882
rect 1526 2878 1530 2882
rect 1662 2878 1666 2882
rect 1742 2878 1746 2882
rect 1790 2878 1794 2882
rect 2070 2878 2074 2882
rect 6 2868 10 2872
rect 54 2868 58 2872
rect 86 2868 90 2872
rect 142 2868 146 2872
rect 158 2868 162 2872
rect 190 2868 194 2872
rect 278 2868 282 2872
rect 294 2868 298 2872
rect 342 2868 346 2872
rect 366 2868 370 2872
rect 422 2868 426 2872
rect 438 2868 442 2872
rect 454 2868 458 2872
rect 502 2868 506 2872
rect 590 2868 594 2872
rect 606 2868 610 2872
rect 654 2868 658 2872
rect 734 2868 738 2872
rect 742 2868 746 2872
rect 790 2868 794 2872
rect 798 2868 802 2872
rect 822 2868 826 2872
rect 918 2868 922 2872
rect 1014 2868 1018 2872
rect 1094 2868 1098 2872
rect 1182 2868 1186 2872
rect 1214 2868 1218 2872
rect 1302 2868 1306 2872
rect 1318 2868 1322 2872
rect 1382 2868 1386 2872
rect 1502 2868 1506 2872
rect 1526 2868 1530 2872
rect 1542 2868 1546 2872
rect 1582 2868 1586 2872
rect 1598 2868 1602 2872
rect 1678 2868 1682 2872
rect 1718 2868 1722 2872
rect 1734 2868 1738 2872
rect 78 2858 82 2862
rect 158 2858 162 2862
rect 182 2858 186 2862
rect 262 2859 266 2863
rect 374 2858 378 2862
rect 430 2858 434 2862
rect 574 2859 578 2863
rect 622 2858 626 2862
rect 662 2858 666 2862
rect 902 2859 906 2863
rect 998 2859 1002 2863
rect 1166 2859 1170 2863
rect 1278 2858 1282 2862
rect 1438 2858 1442 2862
rect 1470 2859 1474 2863
rect 1558 2858 1562 2862
rect 1606 2858 1610 2862
rect 1646 2858 1650 2862
rect 1670 2858 1674 2862
rect 1694 2858 1698 2862
rect 1726 2858 1730 2862
rect 1854 2868 1858 2872
rect 1918 2868 1922 2872
rect 1966 2868 1970 2872
rect 1974 2868 1978 2872
rect 1990 2868 1994 2872
rect 2022 2868 2026 2872
rect 2126 2878 2130 2882
rect 2134 2878 2138 2882
rect 2342 2878 2346 2882
rect 2374 2878 2378 2882
rect 2430 2878 2434 2882
rect 2494 2878 2498 2882
rect 2654 2878 2658 2882
rect 2790 2878 2794 2882
rect 3118 2878 3122 2882
rect 3134 2878 3138 2882
rect 3206 2878 3210 2882
rect 3270 2878 3274 2882
rect 2086 2868 2090 2872
rect 2094 2868 2098 2872
rect 2126 2868 2130 2872
rect 2150 2868 2154 2872
rect 2198 2868 2202 2872
rect 2246 2868 2250 2872
rect 2286 2868 2290 2872
rect 2302 2868 2306 2872
rect 2374 2868 2378 2872
rect 2566 2868 2570 2872
rect 2614 2868 2618 2872
rect 2622 2868 2626 2872
rect 2678 2868 2682 2872
rect 2718 2868 2722 2872
rect 2734 2868 2738 2872
rect 2750 2868 2754 2872
rect 2814 2868 2818 2872
rect 2846 2868 2850 2872
rect 2862 2868 2866 2872
rect 2878 2868 2882 2872
rect 2910 2868 2914 2872
rect 2926 2868 2930 2872
rect 2966 2868 2970 2872
rect 2998 2868 3002 2872
rect 3006 2868 3010 2872
rect 3030 2868 3034 2872
rect 3078 2868 3082 2872
rect 3142 2868 3146 2872
rect 3230 2868 3234 2872
rect 3238 2868 3242 2872
rect 3302 2868 3306 2872
rect 3446 2878 3450 2882
rect 3622 2878 3626 2882
rect 3662 2878 3666 2882
rect 3798 2878 3802 2882
rect 3846 2878 3850 2882
rect 3918 2878 3922 2882
rect 4086 2878 4090 2882
rect 4094 2878 4098 2882
rect 4150 2878 4154 2882
rect 1766 2858 1770 2862
rect 1790 2858 1794 2862
rect 1806 2858 1810 2862
rect 1822 2858 1826 2862
rect 1846 2858 1850 2862
rect 1934 2858 1938 2862
rect 1982 2858 1986 2862
rect 2038 2858 2042 2862
rect 2102 2858 2106 2862
rect 2110 2858 2114 2862
rect 2158 2858 2162 2862
rect 2174 2858 2178 2862
rect 2294 2858 2298 2862
rect 2334 2858 2338 2862
rect 2358 2858 2362 2862
rect 2382 2858 2386 2862
rect 2502 2858 2506 2862
rect 2526 2858 2530 2862
rect 2630 2858 2634 2862
rect 2670 2858 2674 2862
rect 2742 2858 2746 2862
rect 2774 2858 2778 2862
rect 2822 2858 2826 2862
rect 2838 2858 2842 2862
rect 2870 2858 2874 2862
rect 2918 2858 2922 2862
rect 2974 2858 2978 2862
rect 2998 2858 3002 2862
rect 3046 2858 3050 2862
rect 3102 2858 3106 2862
rect 3134 2858 3138 2862
rect 3166 2858 3170 2862
rect 3190 2858 3194 2862
rect 3222 2858 3226 2862
rect 3254 2858 3258 2862
rect 3294 2858 3298 2862
rect 3374 2868 3378 2872
rect 3422 2868 3426 2872
rect 3494 2868 3498 2872
rect 3510 2868 3514 2872
rect 3542 2868 3546 2872
rect 3334 2858 3338 2862
rect 3446 2858 3450 2862
rect 3478 2858 3482 2862
rect 3534 2858 3538 2862
rect 3598 2868 3602 2872
rect 3638 2868 3642 2872
rect 3710 2868 3714 2872
rect 3638 2858 3642 2862
rect 3662 2858 3666 2862
rect 3686 2858 3690 2862
rect 3798 2868 3802 2872
rect 3862 2868 3866 2872
rect 3886 2868 3890 2872
rect 3902 2868 3906 2872
rect 3950 2868 3954 2872
rect 3966 2868 3970 2872
rect 3990 2868 3994 2872
rect 3998 2868 4002 2872
rect 4014 2868 4018 2872
rect 4038 2868 4042 2872
rect 4078 2868 4082 2872
rect 4134 2868 4138 2872
rect 4166 2868 4170 2872
rect 4198 2868 4202 2872
rect 4550 2878 4554 2882
rect 4638 2878 4642 2882
rect 4774 2878 4778 2882
rect 4790 2878 4794 2882
rect 4878 2878 4882 2882
rect 4918 2878 4922 2882
rect 5038 2878 5042 2882
rect 5070 2878 5074 2882
rect 5302 2879 5306 2883
rect 4222 2868 4226 2872
rect 4270 2868 4274 2872
rect 4342 2868 4346 2872
rect 4446 2868 4450 2872
rect 4494 2868 4498 2872
rect 4558 2868 4562 2872
rect 4622 2868 4626 2872
rect 4638 2868 4642 2872
rect 4702 2868 4706 2872
rect 4734 2868 4738 2872
rect 4814 2868 4818 2872
rect 4854 2868 4858 2872
rect 4886 2868 4890 2872
rect 5022 2868 5026 2872
rect 5062 2868 5066 2872
rect 3782 2858 3786 2862
rect 3814 2858 3818 2862
rect 3830 2858 3834 2862
rect 3870 2858 3874 2862
rect 3878 2858 3882 2862
rect 3966 2858 3970 2862
rect 4030 2858 4034 2862
rect 4086 2858 4090 2862
rect 4110 2858 4114 2862
rect 4150 2858 4154 2862
rect 4190 2858 4194 2862
rect 4278 2858 4282 2862
rect 4310 2858 4314 2862
rect 4358 2859 4362 2863
rect 4518 2858 4522 2862
rect 4542 2858 4546 2862
rect 4598 2858 4602 2862
rect 4614 2858 4618 2862
rect 4662 2858 4666 2862
rect 4694 2858 4698 2862
rect 4726 2858 4730 2862
rect 4750 2858 4754 2862
rect 4790 2858 4794 2862
rect 4854 2858 4858 2862
rect 4862 2858 4866 2862
rect 4942 2858 4946 2862
rect 4990 2858 4994 2862
rect 5014 2858 5018 2862
rect 5110 2858 5114 2862
rect 5118 2858 5122 2862
rect 5206 2858 5210 2862
rect 5222 2858 5226 2862
rect 5270 2858 5274 2862
rect 5310 2858 5314 2862
rect 166 2848 170 2852
rect 446 2848 450 2852
rect 798 2848 802 2852
rect 1198 2848 1202 2852
rect 1502 2848 1506 2852
rect 1622 2848 1626 2852
rect 1654 2848 1658 2852
rect 1782 2848 1786 2852
rect 1814 2848 1818 2852
rect 1894 2848 1898 2852
rect 2006 2848 2010 2852
rect 2030 2848 2034 2852
rect 2166 2848 2170 2852
rect 2310 2848 2314 2852
rect 2366 2848 2370 2852
rect 2430 2848 2434 2852
rect 2462 2848 2466 2852
rect 2646 2848 2650 2852
rect 2694 2848 2698 2852
rect 2726 2848 2730 2852
rect 2790 2848 2794 2852
rect 2830 2848 2834 2852
rect 2894 2848 2898 2852
rect 2950 2848 2954 2852
rect 2974 2848 2978 2852
rect 3022 2848 3026 2852
rect 3086 2848 3090 2852
rect 3198 2848 3202 2852
rect 3206 2848 3210 2852
rect 3254 2848 3258 2852
rect 3270 2848 3274 2852
rect 3494 2848 3498 2852
rect 3614 2848 3618 2852
rect 3654 2848 3658 2852
rect 3678 2848 3682 2852
rect 3942 2848 3946 2852
rect 3974 2848 3978 2852
rect 4014 2848 4018 2852
rect 4022 2848 4026 2852
rect 4174 2848 4178 2852
rect 4294 2848 4298 2852
rect 4606 2848 4610 2852
rect 4670 2848 4674 2852
rect 4678 2848 4682 2852
rect 4710 2848 4714 2852
rect 4742 2848 4746 2852
rect 4830 2848 4834 2852
rect 4982 2848 4986 2852
rect 5046 2848 5050 2852
rect 102 2838 106 2842
rect 1558 2838 1562 2842
rect 1582 2838 1586 2842
rect 1638 2838 1642 2842
rect 1830 2838 1834 2842
rect 2046 2838 2050 2842
rect 2070 2838 2074 2842
rect 2182 2838 2186 2842
rect 2254 2838 2258 2842
rect 2630 2838 2634 2842
rect 2678 2838 2682 2842
rect 2686 2838 2690 2842
rect 2766 2838 2770 2842
rect 2790 2838 2794 2842
rect 2814 2838 2818 2842
rect 2942 2838 2946 2842
rect 3182 2838 3186 2842
rect 3694 2838 3698 2842
rect 4038 2838 4042 2842
rect 4118 2838 4122 2842
rect 4142 2838 4146 2842
rect 4574 2838 4578 2842
rect 4590 2838 4594 2842
rect 4654 2838 4658 2842
rect 4662 2838 4666 2842
rect 4758 2838 4762 2842
rect 4862 2838 4866 2842
rect 4950 2838 4954 2842
rect 4998 2838 5002 2842
rect 5286 2838 5290 2842
rect 2038 2828 2042 2832
rect 2774 2828 2778 2832
rect 3686 2828 3690 2832
rect 4110 2828 4114 2832
rect 4598 2828 4602 2832
rect 4942 2828 4946 2832
rect 1542 2818 1546 2822
rect 1606 2818 1610 2822
rect 1646 2818 1650 2822
rect 1822 2818 1826 2822
rect 2174 2818 2178 2822
rect 2222 2818 2226 2822
rect 2350 2818 2354 2822
rect 4662 2818 4666 2822
rect 4694 2818 4698 2822
rect 4726 2818 4730 2822
rect 4750 2818 4754 2822
rect 4782 2818 4786 2822
rect 4798 2818 4802 2822
rect 4894 2818 4898 2822
rect 4990 2818 4994 2822
rect 5038 2818 5042 2822
rect 346 2803 350 2807
rect 353 2803 357 2807
rect 1370 2803 1374 2807
rect 1377 2803 1381 2807
rect 2394 2803 2398 2807
rect 2401 2803 2405 2807
rect 3418 2803 3422 2807
rect 3425 2803 3429 2807
rect 4442 2803 4446 2807
rect 4449 2803 4453 2807
rect 254 2788 258 2792
rect 278 2788 282 2792
rect 374 2788 378 2792
rect 470 2788 474 2792
rect 550 2788 554 2792
rect 646 2788 650 2792
rect 774 2788 778 2792
rect 822 2788 826 2792
rect 918 2788 922 2792
rect 1230 2788 1234 2792
rect 1326 2788 1330 2792
rect 1358 2788 1362 2792
rect 1654 2788 1658 2792
rect 1678 2788 1682 2792
rect 1774 2788 1778 2792
rect 1790 2788 1794 2792
rect 1830 2788 1834 2792
rect 1862 2788 1866 2792
rect 1998 2788 2002 2792
rect 2054 2788 2058 2792
rect 2126 2788 2130 2792
rect 2310 2788 2314 2792
rect 2342 2788 2346 2792
rect 2374 2788 2378 2792
rect 2518 2788 2522 2792
rect 2614 2788 2618 2792
rect 2702 2788 2706 2792
rect 2894 2788 2898 2792
rect 2990 2788 2994 2792
rect 3022 2788 3026 2792
rect 3150 2788 3154 2792
rect 3222 2788 3226 2792
rect 3270 2788 3274 2792
rect 3294 2788 3298 2792
rect 3470 2788 3474 2792
rect 3694 2788 3698 2792
rect 3734 2788 3738 2792
rect 3766 2788 3770 2792
rect 3886 2788 3890 2792
rect 4014 2788 4018 2792
rect 4038 2788 4042 2792
rect 4086 2788 4090 2792
rect 4166 2788 4170 2792
rect 4566 2788 4570 2792
rect 5150 2788 5154 2792
rect 1646 2778 1650 2782
rect 2622 2778 2626 2782
rect 78 2768 82 2772
rect 102 2768 106 2772
rect 262 2768 266 2772
rect 302 2768 306 2772
rect 478 2768 482 2772
rect 542 2768 546 2772
rect 782 2768 786 2772
rect 798 2768 802 2772
rect 1630 2768 1634 2772
rect 1822 2768 1826 2772
rect 1950 2768 1954 2772
rect 1990 2768 1994 2772
rect 2006 2768 2010 2772
rect 2334 2768 2338 2772
rect 2350 2768 2354 2772
rect 2382 2768 2386 2772
rect 2862 2768 2866 2772
rect 3190 2778 3194 2782
rect 4414 2778 4418 2782
rect 2894 2768 2898 2772
rect 2902 2768 2906 2772
rect 2918 2768 2922 2772
rect 2958 2768 2962 2772
rect 2998 2768 3002 2772
rect 3174 2768 3178 2772
rect 3262 2768 3266 2772
rect 3310 2768 3314 2772
rect 3686 2768 3690 2772
rect 3758 2768 3762 2772
rect 3774 2768 3778 2772
rect 3798 2768 3802 2772
rect 3966 2768 3970 2772
rect 4030 2768 4034 2772
rect 4342 2768 4346 2772
rect 4358 2768 4362 2772
rect 4390 2768 4394 2772
rect 4406 2768 4410 2772
rect 4614 2768 4618 2772
rect 54 2758 58 2762
rect 62 2758 66 2762
rect 110 2758 114 2762
rect 222 2758 226 2762
rect 238 2758 242 2762
rect 246 2758 250 2762
rect 22 2748 26 2752
rect 30 2748 34 2752
rect 70 2748 74 2752
rect 86 2748 90 2752
rect 134 2748 138 2752
rect 174 2748 178 2752
rect 182 2748 186 2752
rect 254 2748 258 2752
rect 278 2748 282 2752
rect 390 2758 394 2762
rect 462 2758 466 2762
rect 526 2758 530 2762
rect 806 2758 810 2762
rect 854 2758 858 2762
rect 1190 2758 1194 2762
rect 1246 2758 1250 2762
rect 1702 2758 1706 2762
rect 1758 2758 1762 2762
rect 1782 2758 1786 2762
rect 1814 2758 1818 2762
rect 1902 2758 1906 2762
rect 1934 2758 1938 2762
rect 2334 2758 2338 2762
rect 2366 2758 2370 2762
rect 2406 2758 2410 2762
rect 2790 2758 2794 2762
rect 2830 2758 2834 2762
rect 2838 2758 2842 2762
rect 2878 2758 2882 2762
rect 2886 2758 2890 2762
rect 2934 2758 2938 2762
rect 2982 2758 2986 2762
rect 3158 2758 3162 2762
rect 3286 2758 3290 2762
rect 3302 2758 3306 2762
rect 3598 2758 3602 2762
rect 3630 2758 3634 2762
rect 3670 2758 3674 2762
rect 3702 2758 3706 2762
rect 3742 2758 3746 2762
rect 3814 2758 3818 2762
rect 3846 2758 3850 2762
rect 3982 2758 3986 2762
rect 4046 2758 4050 2762
rect 4062 2758 4066 2762
rect 334 2748 338 2752
rect 350 2748 354 2752
rect 422 2748 426 2752
rect 470 2748 474 2752
rect 494 2748 498 2752
rect 590 2748 594 2752
rect 38 2738 42 2742
rect 118 2738 122 2742
rect 142 2738 146 2742
rect 614 2747 618 2751
rect 678 2748 682 2752
rect 710 2747 714 2751
rect 742 2748 746 2752
rect 774 2748 778 2752
rect 822 2748 826 2752
rect 894 2748 898 2752
rect 958 2748 962 2752
rect 974 2748 978 2752
rect 998 2748 1002 2752
rect 1078 2748 1082 2752
rect 1110 2748 1114 2752
rect 1118 2748 1122 2752
rect 1158 2748 1162 2752
rect 1182 2748 1186 2752
rect 1198 2748 1202 2752
rect 1230 2748 1234 2752
rect 206 2738 210 2742
rect 310 2738 314 2742
rect 342 2738 346 2742
rect 366 2738 370 2742
rect 414 2738 418 2742
rect 510 2740 514 2744
rect 526 2738 530 2742
rect 542 2738 546 2742
rect 830 2738 834 2742
rect 838 2738 842 2742
rect 902 2738 906 2742
rect 950 2738 954 2742
rect 1022 2738 1026 2742
rect 1086 2738 1090 2742
rect 1118 2738 1122 2742
rect 1422 2747 1426 2751
rect 1550 2748 1554 2752
rect 1582 2747 1586 2751
rect 1734 2748 1738 2752
rect 1814 2748 1818 2752
rect 1838 2748 1842 2752
rect 1918 2748 1922 2752
rect 1934 2748 1938 2752
rect 1998 2748 2002 2752
rect 2022 2748 2026 2752
rect 2182 2748 2186 2752
rect 2246 2747 2250 2751
rect 2342 2748 2346 2752
rect 2374 2748 2378 2752
rect 2454 2747 2458 2751
rect 2550 2747 2554 2751
rect 2582 2748 2586 2752
rect 2726 2748 2730 2752
rect 2814 2748 2818 2752
rect 2830 2748 2834 2752
rect 2870 2748 2874 2752
rect 2894 2748 2898 2752
rect 2942 2748 2946 2752
rect 2974 2748 2978 2752
rect 2990 2748 2994 2752
rect 3014 2748 3018 2752
rect 3038 2748 3042 2752
rect 3126 2748 3130 2752
rect 3166 2748 3170 2752
rect 3246 2748 3250 2752
rect 3270 2748 3274 2752
rect 3326 2748 3330 2752
rect 3414 2748 3418 2752
rect 3454 2748 3458 2752
rect 3462 2748 3466 2752
rect 3598 2748 3602 2752
rect 3630 2748 3634 2752
rect 3654 2748 3658 2752
rect 3670 2748 3674 2752
rect 3694 2748 3698 2752
rect 3710 2748 3714 2752
rect 3750 2748 3754 2752
rect 3798 2748 3802 2752
rect 3822 2748 3826 2752
rect 3838 2748 3842 2752
rect 3862 2748 3866 2752
rect 3942 2748 3946 2752
rect 3998 2748 4002 2752
rect 4038 2748 4042 2752
rect 4054 2748 4058 2752
rect 4102 2758 4106 2762
rect 4142 2758 4146 2762
rect 4446 2758 4450 2762
rect 4510 2758 4514 2762
rect 4598 2758 4602 2762
rect 4630 2758 4634 2762
rect 4710 2758 4714 2762
rect 4718 2758 4722 2762
rect 4926 2758 4930 2762
rect 5278 2758 5282 2762
rect 4150 2748 4154 2752
rect 4206 2748 4210 2752
rect 1190 2738 1194 2742
rect 1214 2738 1218 2742
rect 1222 2738 1226 2742
rect 1254 2738 1258 2742
rect 1270 2738 1274 2742
rect 1438 2738 1442 2742
rect 1454 2738 1458 2742
rect 1518 2738 1522 2742
rect 1566 2738 1570 2742
rect 1702 2738 1706 2742
rect 1726 2738 1730 2742
rect 1742 2738 1746 2742
rect 1766 2738 1770 2742
rect 1838 2738 1842 2742
rect 1910 2738 1914 2742
rect 1926 2738 1930 2742
rect 1950 2738 1954 2742
rect 1966 2738 1970 2742
rect 2070 2738 2074 2742
rect 2118 2738 2122 2742
rect 2438 2738 2442 2742
rect 2534 2738 2538 2742
rect 2638 2738 2642 2742
rect 2686 2738 2690 2742
rect 2734 2738 2738 2742
rect 2782 2738 2786 2742
rect 2790 2738 2794 2742
rect 2806 2738 2810 2742
rect 4294 2747 4298 2751
rect 4414 2748 4418 2752
rect 4430 2748 4434 2752
rect 4462 2748 4466 2752
rect 4494 2748 4498 2752
rect 4502 2748 4506 2752
rect 4542 2748 4546 2752
rect 4622 2748 4626 2752
rect 4742 2748 4746 2752
rect 4758 2748 4762 2752
rect 4886 2748 4890 2752
rect 4966 2748 4970 2752
rect 5014 2748 5018 2752
rect 5030 2748 5034 2752
rect 5102 2748 5106 2752
rect 5214 2747 5218 2751
rect 5262 2748 5266 2752
rect 5302 2748 5306 2752
rect 3030 2738 3034 2742
rect 3070 2738 3074 2742
rect 3118 2738 3122 2742
rect 3134 2738 3138 2742
rect 3182 2738 3186 2742
rect 3238 2738 3242 2742
rect 3286 2738 3290 2742
rect 3334 2738 3338 2742
rect 3342 2738 3346 2742
rect 3390 2738 3394 2742
rect 3486 2738 3490 2742
rect 3534 2738 3538 2742
rect 3542 2738 3546 2742
rect 3590 2738 3594 2742
rect 3622 2738 3626 2742
rect 3646 2738 3650 2742
rect 3718 2738 3722 2742
rect 3790 2738 3794 2742
rect 3870 2738 3874 2742
rect 3894 2738 3898 2742
rect 3958 2738 3962 2742
rect 3966 2738 3970 2742
rect 3982 2738 3986 2742
rect 4078 2738 4082 2742
rect 4094 2738 4098 2742
rect 4142 2738 4146 2742
rect 4182 2738 4186 2742
rect 54 2728 58 2732
rect 102 2728 106 2732
rect 190 2728 194 2732
rect 294 2728 298 2732
rect 318 2728 322 2732
rect 414 2728 418 2732
rect 742 2728 746 2732
rect 798 2728 802 2732
rect 958 2728 962 2732
rect 982 2728 986 2732
rect 1134 2728 1138 2732
rect 1158 2728 1162 2732
rect 1262 2728 1266 2732
rect 1662 2728 1666 2732
rect 1670 2728 1674 2732
rect 1758 2728 1762 2732
rect 1798 2728 1802 2732
rect 1878 2728 1882 2732
rect 1974 2728 1978 2732
rect 2038 2728 2042 2732
rect 2062 2728 2066 2732
rect 2246 2728 2250 2732
rect 4278 2738 4282 2742
rect 4374 2738 4378 2742
rect 4486 2738 4490 2742
rect 4534 2738 4538 2742
rect 4582 2738 4586 2742
rect 4638 2738 4642 2742
rect 4686 2738 4690 2742
rect 4694 2738 4698 2742
rect 4742 2738 4746 2742
rect 4774 2738 4778 2742
rect 4814 2738 4818 2742
rect 4830 2738 4834 2742
rect 4846 2738 4850 2742
rect 4878 2738 4882 2742
rect 4902 2738 4906 2742
rect 4942 2738 4946 2742
rect 4974 2738 4978 2742
rect 5022 2738 5026 2742
rect 5110 2738 5114 2742
rect 5206 2738 5210 2742
rect 2422 2728 2426 2732
rect 2630 2728 2634 2732
rect 2694 2728 2698 2732
rect 2718 2727 2722 2731
rect 2790 2728 2794 2732
rect 2838 2728 2842 2732
rect 2974 2728 2978 2732
rect 3030 2728 3034 2732
rect 3054 2728 3058 2732
rect 3062 2728 3066 2732
rect 3150 2728 3154 2732
rect 3198 2728 3202 2732
rect 3206 2728 3210 2732
rect 3478 2728 3482 2732
rect 3630 2728 3634 2732
rect 3734 2728 3738 2732
rect 3782 2728 3786 2732
rect 3838 2728 3842 2732
rect 3846 2728 3850 2732
rect 3886 2728 3890 2732
rect 4070 2728 4074 2732
rect 4126 2728 4130 2732
rect 4230 2728 4234 2732
rect 4366 2728 4370 2732
rect 4430 2728 4434 2732
rect 4478 2728 4482 2732
rect 4526 2728 4530 2732
rect 4758 2728 4762 2732
rect 4790 2728 4794 2732
rect 4798 2728 4802 2732
rect 4814 2728 4818 2732
rect 4862 2728 4866 2732
rect 4870 2728 4874 2732
rect 4894 2728 4898 2732
rect 4990 2728 4994 2732
rect 4998 2728 5002 2732
rect 5278 2728 5282 2732
rect 166 2718 170 2722
rect 414 2718 418 2722
rect 862 2718 866 2722
rect 990 2718 994 2722
rect 1118 2718 1122 2722
rect 1166 2718 1170 2722
rect 1230 2718 1234 2722
rect 1718 2718 1722 2722
rect 1958 2718 1962 2722
rect 2102 2718 2106 2722
rect 2654 2718 2658 2722
rect 3078 2718 3082 2722
rect 3102 2718 3106 2722
rect 3310 2718 3314 2722
rect 3374 2718 3378 2722
rect 3382 2718 3386 2722
rect 3518 2718 3522 2722
rect 3526 2718 3530 2722
rect 3574 2718 3578 2722
rect 3582 2718 3586 2722
rect 3614 2718 3618 2722
rect 3798 2718 3802 2722
rect 3958 2718 3962 2722
rect 4262 2718 4266 2722
rect 4454 2718 4458 2722
rect 4574 2718 4578 2722
rect 4598 2718 4602 2722
rect 4622 2718 4626 2722
rect 4670 2718 4674 2722
rect 4710 2718 4714 2722
rect 4726 2718 4730 2722
rect 4750 2718 4754 2722
rect 4782 2718 4786 2722
rect 4822 2718 4826 2722
rect 4854 2718 4858 2722
rect 4918 2718 4922 2722
rect 4982 2718 4986 2722
rect 5006 2718 5010 2722
rect 5046 2718 5050 2722
rect 5054 2718 5058 2722
rect 462 2708 466 2712
rect 1158 2708 1162 2712
rect 3198 2708 3202 2712
rect 3478 2708 3482 2712
rect 3838 2708 3842 2712
rect 4054 2708 4058 2712
rect 4070 2708 4074 2712
rect 4366 2708 4370 2712
rect 4478 2708 4482 2712
rect 5278 2708 5282 2712
rect 858 2703 862 2707
rect 865 2703 869 2707
rect 1874 2703 1878 2707
rect 1881 2703 1885 2707
rect 2906 2703 2910 2707
rect 2913 2703 2917 2707
rect 3930 2703 3934 2707
rect 3937 2703 3941 2707
rect 4954 2703 4958 2707
rect 4961 2703 4965 2707
rect 30 2698 34 2702
rect 614 2698 618 2702
rect 998 2698 1002 2702
rect 1966 2698 1970 2702
rect 2310 2698 2314 2702
rect 3166 2698 3170 2702
rect 3334 2698 3338 2702
rect 3350 2698 3354 2702
rect 3622 2698 3626 2702
rect 3646 2698 3650 2702
rect 3910 2698 3914 2702
rect 4278 2698 4282 2702
rect 62 2688 66 2692
rect 86 2688 90 2692
rect 182 2688 186 2692
rect 230 2688 234 2692
rect 390 2688 394 2692
rect 486 2688 490 2692
rect 502 2688 506 2692
rect 518 2688 522 2692
rect 558 2688 562 2692
rect 574 2688 578 2692
rect 606 2688 610 2692
rect 654 2688 658 2692
rect 686 2688 690 2692
rect 766 2688 770 2692
rect 814 2688 818 2692
rect 838 2688 842 2692
rect 854 2688 858 2692
rect 934 2688 938 2692
rect 1006 2688 1010 2692
rect 1038 2688 1042 2692
rect 1086 2688 1090 2692
rect 1094 2688 1098 2692
rect 1182 2688 1186 2692
rect 1286 2688 1290 2692
rect 1326 2688 1330 2692
rect 1398 2688 1402 2692
rect 1494 2688 1498 2692
rect 1590 2688 1594 2692
rect 1798 2688 1802 2692
rect 1894 2688 1898 2692
rect 1934 2688 1938 2692
rect 2046 2688 2050 2692
rect 2078 2688 2082 2692
rect 2142 2688 2146 2692
rect 2230 2688 2234 2692
rect 2342 2688 2346 2692
rect 2398 2688 2402 2692
rect 2414 2688 2418 2692
rect 2518 2688 2522 2692
rect 2566 2688 2570 2692
rect 2598 2688 2602 2692
rect 2662 2688 2666 2692
rect 2758 2688 2762 2692
rect 2926 2688 2930 2692
rect 3038 2688 3042 2692
rect 3054 2688 3058 2692
rect 3134 2688 3138 2692
rect 3174 2688 3178 2692
rect 3238 2688 3242 2692
rect 3294 2688 3298 2692
rect 3446 2688 3450 2692
rect 3470 2688 3474 2692
rect 3574 2688 3578 2692
rect 3582 2688 3586 2692
rect 3662 2688 3666 2692
rect 3686 2688 3690 2692
rect 3782 2688 3786 2692
rect 3798 2688 3802 2692
rect 3814 2688 3818 2692
rect 3854 2688 3858 2692
rect 3862 2688 3866 2692
rect 3894 2688 3898 2692
rect 3950 2688 3954 2692
rect 4078 2688 4082 2692
rect 4302 2688 4306 2692
rect 4350 2688 4354 2692
rect 4414 2688 4418 2692
rect 4430 2688 4434 2692
rect 4478 2688 4482 2692
rect 4494 2688 4498 2692
rect 4614 2688 4618 2692
rect 4934 2688 4938 2692
rect 30 2678 34 2682
rect 118 2678 122 2682
rect 262 2678 266 2682
rect 358 2678 362 2682
rect 478 2678 482 2682
rect 614 2678 618 2682
rect 662 2678 666 2682
rect 742 2678 746 2682
rect 822 2678 826 2682
rect 926 2678 930 2682
rect 998 2678 1002 2682
rect 1062 2678 1066 2682
rect 1158 2678 1162 2682
rect 1694 2679 1698 2683
rect 1918 2678 1922 2682
rect 1966 2678 1970 2682
rect 2134 2678 2138 2682
rect 2286 2678 2290 2682
rect 2302 2678 2306 2682
rect 2310 2678 2314 2682
rect 2638 2678 2642 2682
rect 2902 2678 2906 2682
rect 2942 2678 2946 2682
rect 3166 2678 3170 2682
rect 3230 2678 3234 2682
rect 3262 2678 3266 2682
rect 3350 2678 3354 2682
rect 3622 2678 3626 2682
rect 3822 2678 3826 2682
rect 3910 2678 3914 2682
rect 54 2668 58 2672
rect 70 2668 74 2672
rect 78 2668 82 2672
rect 110 2668 114 2672
rect 142 2668 146 2672
rect 158 2668 162 2672
rect 198 2668 202 2672
rect 206 2668 210 2672
rect 254 2668 258 2672
rect 294 2668 298 2672
rect 350 2668 354 2672
rect 374 2668 378 2672
rect 406 2668 410 2672
rect 414 2668 418 2672
rect 430 2668 434 2672
rect 438 2668 442 2672
rect 462 2668 466 2672
rect 510 2668 514 2672
rect 542 2668 546 2672
rect 550 2668 554 2672
rect 590 2668 594 2672
rect 614 2668 618 2672
rect 638 2668 642 2672
rect 670 2668 674 2672
rect 718 2668 722 2672
rect 742 2668 746 2672
rect 798 2668 802 2672
rect 846 2668 850 2672
rect 894 2668 898 2672
rect 942 2668 946 2672
rect 1030 2668 1034 2672
rect 1062 2668 1066 2672
rect 1078 2668 1082 2672
rect 1118 2668 1122 2672
rect 1222 2668 1226 2672
rect 1238 2668 1242 2672
rect 1254 2668 1258 2672
rect 1262 2668 1266 2672
rect 1358 2668 1362 2672
rect 1374 2668 1378 2672
rect 1550 2668 1554 2672
rect 1718 2668 1722 2672
rect 1814 2668 1818 2672
rect 1926 2668 1930 2672
rect 1966 2668 1970 2672
rect 1990 2668 1994 2672
rect 2006 2668 2010 2672
rect 4142 2678 4146 2682
rect 4198 2678 4202 2682
rect 4262 2678 4266 2682
rect 4278 2678 4282 2682
rect 4366 2678 4370 2682
rect 4398 2679 4402 2683
rect 4646 2678 4650 2682
rect 5182 2678 5186 2682
rect 2022 2666 2026 2670
rect 2126 2668 2130 2672
rect 2174 2668 2178 2672
rect 2214 2666 2218 2670
rect 2254 2666 2258 2670
rect 2262 2668 2266 2672
rect 2270 2668 2274 2672
rect 2310 2668 2314 2672
rect 2398 2668 2402 2672
rect 2406 2668 2410 2672
rect 2438 2668 2442 2672
rect 2526 2668 2530 2672
rect 2574 2668 2578 2672
rect 2582 2668 2586 2672
rect 2742 2668 2746 2672
rect 2838 2668 2842 2672
rect 2854 2668 2858 2672
rect 2886 2668 2890 2672
rect 2894 2668 2898 2672
rect 2958 2668 2962 2672
rect 3046 2668 3050 2672
rect 3094 2668 3098 2672
rect 3126 2668 3130 2672
rect 3142 2668 3146 2672
rect 3198 2668 3202 2672
rect 3206 2668 3210 2672
rect 3222 2668 3226 2672
rect 3246 2668 3250 2672
rect 3334 2668 3338 2672
rect 3550 2668 3554 2672
rect 3566 2668 3570 2672
rect 3614 2668 3618 2672
rect 3646 2668 3650 2672
rect 3670 2668 3674 2672
rect 3726 2668 3730 2672
rect 3790 2668 3794 2672
rect 3838 2668 3842 2672
rect 3894 2668 3898 2672
rect 3918 2668 3922 2672
rect 4054 2668 4058 2672
rect 4086 2668 4090 2672
rect 4094 2668 4098 2672
rect 4126 2668 4130 2672
rect 4150 2668 4154 2672
rect 4214 2668 4218 2672
rect 4286 2668 4290 2672
rect 4302 2668 4306 2672
rect 4334 2668 4338 2672
rect 4358 2668 4362 2672
rect 4374 2668 4378 2672
rect 4382 2668 4386 2672
rect 4430 2668 4434 2672
rect 4454 2668 4458 2672
rect 4486 2668 4490 2672
rect 4534 2668 4538 2672
rect 4542 2668 4546 2672
rect 4598 2668 4602 2672
rect 4614 2668 4618 2672
rect 4654 2668 4658 2672
rect 4702 2668 4706 2672
rect 4742 2668 4746 2672
rect 4790 2668 4794 2672
rect 4822 2668 4826 2672
rect 4878 2668 4882 2672
rect 4918 2668 4922 2672
rect 5142 2668 5146 2672
rect 5294 2668 5298 2672
rect 6 2658 10 2662
rect 46 2658 50 2662
rect 86 2658 90 2662
rect 102 2658 106 2662
rect 166 2658 170 2662
rect 302 2658 306 2662
rect 318 2658 322 2662
rect 382 2658 386 2662
rect 454 2658 458 2662
rect 462 2658 466 2662
rect 502 2658 506 2662
rect 534 2658 538 2662
rect 598 2658 602 2662
rect 614 2658 618 2662
rect 806 2658 810 2662
rect 886 2658 890 2662
rect 918 2658 922 2662
rect 950 2658 954 2662
rect 974 2658 978 2662
rect 982 2658 986 2662
rect 1022 2658 1026 2662
rect 1054 2658 1058 2662
rect 1086 2658 1090 2662
rect 1110 2658 1114 2662
rect 1142 2658 1146 2662
rect 1222 2658 1226 2662
rect 1246 2658 1250 2662
rect 1270 2658 1274 2662
rect 1302 2658 1306 2662
rect 1342 2658 1346 2662
rect 1438 2658 1442 2662
rect 1462 2659 1466 2663
rect 1558 2659 1562 2663
rect 1630 2658 1634 2662
rect 1646 2658 1650 2662
rect 1702 2658 1706 2662
rect 1734 2659 1738 2663
rect 1830 2659 1834 2663
rect 1950 2658 1954 2662
rect 1982 2658 1986 2662
rect 2038 2658 2042 2662
rect 2062 2658 2066 2662
rect 2094 2658 2098 2662
rect 2182 2658 2186 2662
rect 2286 2658 2290 2662
rect 2326 2658 2330 2662
rect 2374 2658 2378 2662
rect 2454 2659 2458 2663
rect 2558 2658 2562 2662
rect 2654 2658 2658 2662
rect 2702 2658 2706 2662
rect 2806 2658 2810 2662
rect 2862 2658 2866 2662
rect 2974 2659 2978 2663
rect 3118 2658 3122 2662
rect 3150 2658 3154 2662
rect 3166 2658 3170 2662
rect 3190 2658 3194 2662
rect 3254 2658 3258 2662
rect 3278 2658 3282 2662
rect 3294 2658 3298 2662
rect 3318 2658 3322 2662
rect 3382 2659 3386 2663
rect 3414 2658 3418 2662
rect 3510 2658 3514 2662
rect 3526 2658 3530 2662
rect 3638 2658 3642 2662
rect 3718 2659 3722 2663
rect 3798 2658 3802 2662
rect 3838 2658 3842 2662
rect 3878 2658 3882 2662
rect 3982 2659 3986 2663
rect 4014 2658 4018 2662
rect 4062 2658 4066 2662
rect 4102 2658 4106 2662
rect 4158 2658 4162 2662
rect 4222 2658 4226 2662
rect 4238 2658 4242 2662
rect 4262 2658 4266 2662
rect 4326 2658 4330 2662
rect 4390 2658 4394 2662
rect 4462 2658 4466 2662
rect 4502 2658 4506 2662
rect 4622 2658 4626 2662
rect 4718 2658 4722 2662
rect 4814 2658 4818 2662
rect 4894 2658 4898 2662
rect 4998 2658 5002 2662
rect 5038 2658 5042 2662
rect 5070 2658 5074 2662
rect 5094 2658 5098 2662
rect 5134 2658 5138 2662
rect 5198 2658 5202 2662
rect 5238 2658 5242 2662
rect 5270 2658 5274 2662
rect 5286 2658 5290 2662
rect 54 2648 58 2652
rect 126 2648 130 2652
rect 142 2648 146 2652
rect 174 2648 178 2652
rect 182 2648 186 2652
rect 310 2648 314 2652
rect 390 2648 394 2652
rect 414 2648 418 2652
rect 438 2648 442 2652
rect 478 2648 482 2652
rect 566 2648 570 2652
rect 646 2648 650 2652
rect 742 2648 746 2652
rect 830 2648 834 2652
rect 998 2648 1002 2652
rect 1038 2648 1042 2652
rect 1094 2648 1098 2652
rect 1198 2648 1202 2652
rect 1230 2648 1234 2652
rect 1294 2648 1298 2652
rect 1358 2648 1362 2652
rect 1374 2648 1378 2652
rect 1934 2648 1938 2652
rect 2006 2648 2010 2652
rect 2070 2648 2074 2652
rect 2198 2648 2202 2652
rect 2238 2648 2242 2652
rect 2286 2648 2290 2652
rect 2334 2648 2338 2652
rect 2358 2648 2362 2652
rect 2422 2648 2426 2652
rect 2878 2648 2882 2652
rect 3142 2648 3146 2652
rect 3174 2648 3178 2652
rect 3222 2648 3226 2652
rect 3294 2648 3298 2652
rect 3302 2648 3306 2652
rect 3662 2648 3666 2652
rect 3686 2648 3690 2652
rect 3822 2648 3826 2652
rect 3854 2648 3858 2652
rect 3862 2648 3866 2652
rect 3902 2648 3906 2652
rect 3934 2648 3938 2652
rect 4078 2648 4082 2652
rect 4190 2648 4194 2652
rect 4230 2648 4234 2652
rect 4286 2648 4290 2652
rect 4302 2648 4306 2652
rect 4414 2648 4418 2652
rect 4614 2648 4618 2652
rect 4710 2648 4714 2652
rect 4798 2648 4802 2652
rect 4854 2648 4858 2652
rect 4878 2648 4882 2652
rect 4990 2648 4994 2652
rect 5022 2648 5026 2652
rect 5046 2648 5050 2652
rect 5078 2648 5082 2652
rect 5086 2648 5090 2652
rect 5118 2648 5122 2652
rect 5182 2648 5186 2652
rect 5190 2648 5194 2652
rect 5270 2648 5274 2652
rect 158 2638 162 2642
rect 326 2638 330 2642
rect 966 2638 970 2642
rect 1134 2638 1138 2642
rect 1302 2638 1306 2642
rect 1310 2638 1314 2642
rect 1510 2638 1514 2642
rect 1606 2638 1610 2642
rect 1990 2638 1994 2642
rect 2054 2638 2058 2642
rect 3334 2638 3338 2642
rect 3646 2638 3650 2642
rect 4246 2638 4250 2642
rect 4334 2638 4338 2642
rect 4574 2638 4578 2642
rect 4646 2638 4650 2642
rect 4686 2638 4690 2642
rect 4726 2638 4730 2642
rect 4862 2638 4866 2642
rect 4902 2638 4906 2642
rect 5006 2638 5010 2642
rect 5030 2638 5034 2642
rect 5062 2638 5066 2642
rect 5094 2638 5098 2642
rect 5102 2638 5106 2642
rect 5158 2638 5162 2642
rect 958 2628 962 2632
rect 1998 2628 2002 2632
rect 5134 2628 5138 2632
rect 278 2618 282 2622
rect 318 2618 322 2622
rect 1126 2618 1130 2622
rect 3062 2618 3066 2622
rect 4046 2618 4050 2622
rect 4182 2618 4186 2622
rect 4238 2618 4242 2622
rect 4718 2618 4722 2622
rect 4758 2618 4762 2622
rect 4814 2618 4818 2622
rect 4870 2618 4874 2622
rect 4894 2618 4898 2622
rect 4998 2618 5002 2622
rect 5094 2618 5098 2622
rect 5286 2618 5290 2622
rect 346 2603 350 2607
rect 353 2603 357 2607
rect 1370 2603 1374 2607
rect 1377 2603 1381 2607
rect 2394 2603 2398 2607
rect 2401 2603 2405 2607
rect 3418 2603 3422 2607
rect 3425 2603 3429 2607
rect 4442 2603 4446 2607
rect 4449 2603 4453 2607
rect 94 2588 98 2592
rect 350 2588 354 2592
rect 446 2588 450 2592
rect 542 2588 546 2592
rect 550 2588 554 2592
rect 574 2588 578 2592
rect 662 2588 666 2592
rect 694 2588 698 2592
rect 718 2588 722 2592
rect 790 2588 794 2592
rect 822 2588 826 2592
rect 846 2588 850 2592
rect 894 2588 898 2592
rect 1006 2588 1010 2592
rect 1078 2588 1082 2592
rect 1102 2588 1106 2592
rect 1182 2588 1186 2592
rect 1214 2588 1218 2592
rect 1310 2588 1314 2592
rect 1342 2588 1346 2592
rect 1350 2588 1354 2592
rect 1454 2588 1458 2592
rect 1558 2588 1562 2592
rect 1654 2588 1658 2592
rect 1702 2588 1706 2592
rect 1726 2588 1730 2592
rect 1734 2588 1738 2592
rect 1750 2588 1754 2592
rect 1950 2588 1954 2592
rect 2142 2588 2146 2592
rect 2206 2588 2210 2592
rect 2366 2588 2370 2592
rect 2422 2588 2426 2592
rect 2510 2588 2514 2592
rect 2518 2588 2522 2592
rect 2654 2588 2658 2592
rect 2662 2588 2666 2592
rect 2910 2588 2914 2592
rect 3030 2588 3034 2592
rect 3054 2588 3058 2592
rect 3158 2588 3162 2592
rect 3262 2588 3266 2592
rect 3606 2588 3610 2592
rect 3702 2588 3706 2592
rect 3718 2588 3722 2592
rect 4262 2588 4266 2592
rect 4334 2588 4338 2592
rect 4910 2588 4914 2592
rect 486 2578 490 2582
rect 734 2578 738 2582
rect 1198 2578 1202 2582
rect 1958 2578 1962 2582
rect 2270 2578 2274 2582
rect 4670 2578 4674 2582
rect 742 2568 746 2572
rect 758 2568 762 2572
rect 1110 2568 1114 2572
rect 2622 2568 2626 2572
rect 3118 2568 3122 2572
rect 3150 2568 3154 2572
rect 3982 2568 3986 2572
rect 3990 2568 3994 2572
rect 4014 2568 4018 2572
rect 4174 2568 4178 2572
rect 4430 2568 4434 2572
rect 4470 2568 4474 2572
rect 4478 2568 4482 2572
rect 4494 2568 4498 2572
rect 4662 2568 4666 2572
rect 4846 2568 4850 2572
rect 5142 2568 5146 2572
rect 30 2558 34 2562
rect 142 2558 146 2562
rect 198 2558 202 2562
rect 278 2558 282 2562
rect 590 2558 594 2562
rect 614 2558 618 2562
rect 670 2558 674 2562
rect 678 2558 682 2562
rect 774 2558 778 2562
rect 862 2558 866 2562
rect 998 2558 1002 2562
rect 1086 2558 1090 2562
rect 1094 2558 1098 2562
rect 1662 2558 1666 2562
rect 2406 2558 2410 2562
rect 3038 2558 3042 2562
rect 3070 2558 3074 2562
rect 3110 2558 3114 2562
rect 3134 2558 3138 2562
rect 3166 2558 3170 2562
rect 3398 2558 3402 2562
rect 3854 2558 3858 2562
rect 4030 2558 4034 2562
rect 4390 2558 4394 2562
rect 4406 2558 4410 2562
rect 4414 2558 4418 2562
rect 4566 2558 4570 2562
rect 4582 2558 4586 2562
rect 4622 2558 4626 2562
rect 4678 2558 4682 2562
rect 4702 2558 4706 2562
rect 4830 2558 4834 2562
rect 4982 2558 4986 2562
rect 5014 2558 5018 2562
rect 14 2548 18 2552
rect 38 2548 42 2552
rect 54 2548 58 2552
rect 126 2548 130 2552
rect 150 2548 154 2552
rect 166 2548 170 2552
rect 262 2548 266 2552
rect 310 2548 314 2552
rect 390 2548 394 2552
rect 414 2548 418 2552
rect 454 2548 458 2552
rect 478 2548 482 2552
rect 502 2548 506 2552
rect 542 2548 546 2552
rect 574 2548 578 2552
rect 630 2548 634 2552
rect 702 2548 706 2552
rect 766 2548 770 2552
rect 782 2548 786 2552
rect 814 2548 818 2552
rect 854 2548 858 2552
rect 894 2548 898 2552
rect 982 2548 986 2552
rect 1046 2548 1050 2552
rect 1062 2548 1066 2552
rect 1102 2548 1106 2552
rect 6 2538 10 2542
rect 62 2538 66 2542
rect 118 2538 122 2542
rect 134 2538 138 2542
rect 174 2538 178 2542
rect 206 2538 210 2542
rect 254 2538 258 2542
rect 302 2538 306 2542
rect 318 2538 322 2542
rect 1278 2547 1282 2551
rect 1390 2548 1394 2552
rect 1422 2547 1426 2551
rect 1518 2547 1522 2551
rect 1614 2548 1618 2552
rect 1710 2548 1714 2552
rect 1814 2547 1818 2551
rect 1886 2547 1890 2551
rect 2022 2547 2026 2551
rect 2078 2547 2082 2551
rect 2110 2548 2114 2552
rect 2166 2548 2170 2552
rect 2238 2548 2242 2552
rect 2302 2547 2306 2551
rect 2334 2548 2338 2552
rect 2558 2548 2562 2552
rect 2726 2547 2730 2551
rect 2758 2548 2762 2552
rect 2854 2548 2858 2552
rect 2966 2547 2970 2551
rect 3062 2548 3066 2552
rect 3094 2548 3098 2552
rect 3110 2548 3114 2552
rect 3158 2548 3162 2552
rect 3198 2547 3202 2551
rect 3294 2547 3298 2551
rect 3326 2548 3330 2552
rect 3446 2548 3450 2552
rect 3478 2548 3482 2552
rect 3542 2547 3546 2551
rect 3574 2548 3578 2552
rect 3638 2547 3642 2551
rect 3670 2548 3674 2552
rect 3774 2548 3778 2552
rect 3814 2548 3818 2552
rect 3894 2548 3898 2552
rect 3902 2548 3906 2552
rect 3918 2548 3922 2552
rect 3990 2548 3994 2552
rect 4022 2548 4026 2552
rect 4062 2548 4066 2552
rect 4126 2547 4130 2551
rect 4158 2548 4162 2552
rect 4198 2548 4202 2552
rect 4422 2548 4426 2552
rect 4478 2548 4482 2552
rect 4510 2548 4514 2552
rect 4526 2548 4530 2552
rect 4542 2548 4546 2552
rect 4558 2548 4562 2552
rect 4582 2548 4586 2552
rect 4622 2548 4626 2552
rect 4630 2548 4634 2552
rect 4670 2548 4674 2552
rect 4710 2548 4714 2552
rect 4790 2548 4794 2552
rect 4798 2548 4802 2552
rect 4838 2548 4842 2552
rect 4862 2548 4866 2552
rect 4886 2548 4890 2552
rect 4934 2548 4938 2552
rect 5014 2548 5018 2552
rect 5286 2548 5290 2552
rect 566 2538 570 2542
rect 598 2538 602 2542
rect 638 2538 642 2542
rect 654 2538 658 2542
rect 710 2538 714 2542
rect 782 2538 786 2542
rect 806 2538 810 2542
rect 902 2538 906 2542
rect 950 2538 954 2542
rect 974 2538 978 2542
rect 990 2538 994 2542
rect 1054 2538 1058 2542
rect 1070 2538 1074 2542
rect 1126 2538 1130 2542
rect 1174 2538 1178 2542
rect 1206 2538 1210 2542
rect 1294 2538 1298 2542
rect 1438 2538 1442 2542
rect 1510 2538 1514 2542
rect 1606 2538 1610 2542
rect 1678 2538 1682 2542
rect 1806 2538 1810 2542
rect 2222 2538 2226 2542
rect 2254 2538 2258 2542
rect 2374 2538 2378 2542
rect 2398 2538 2402 2542
rect 2478 2538 2482 2542
rect 2494 2538 2498 2542
rect 2598 2538 2602 2542
rect 2638 2538 2642 2542
rect 2710 2538 2714 2542
rect 2774 2538 2778 2542
rect 2798 2538 2802 2542
rect 2830 2538 2834 2542
rect 2854 2538 2858 2542
rect 2950 2538 2954 2542
rect 3062 2538 3066 2542
rect 3086 2538 3090 2542
rect 3118 2538 3122 2542
rect 3406 2538 3410 2542
rect 3550 2538 3554 2542
rect 3742 2538 3746 2542
rect 3838 2538 3842 2542
rect 3878 2538 3882 2542
rect 3910 2538 3914 2542
rect 4054 2538 4058 2542
rect 4086 2538 4090 2542
rect 4246 2538 4250 2542
rect 4302 2538 4306 2542
rect 4350 2538 4354 2542
rect 4366 2538 4370 2542
rect 4390 2538 4394 2542
rect 4406 2538 4410 2542
rect 4534 2538 4538 2542
rect 4590 2538 4594 2542
rect 4686 2538 4690 2542
rect 4718 2538 4722 2542
rect 4734 2538 4738 2542
rect 4806 2538 4810 2542
rect 4894 2538 4898 2542
rect 4942 2538 4946 2542
rect 4966 2538 4970 2542
rect 4990 2538 4994 2542
rect 5022 2538 5026 2542
rect 5070 2538 5074 2542
rect 5094 2538 5098 2542
rect 5110 2538 5114 2542
rect 5158 2538 5162 2542
rect 5182 2538 5186 2542
rect 5198 2538 5202 2542
rect 5246 2538 5250 2542
rect 5254 2538 5258 2542
rect 38 2528 42 2532
rect 150 2528 154 2532
rect 438 2528 442 2532
rect 494 2528 498 2532
rect 518 2528 522 2532
rect 526 2528 530 2532
rect 558 2528 562 2532
rect 726 2528 730 2532
rect 742 2528 746 2532
rect 830 2528 834 2532
rect 838 2528 842 2532
rect 966 2528 970 2532
rect 1014 2528 1018 2532
rect 1022 2528 1026 2532
rect 1190 2528 1194 2532
rect 1318 2528 1322 2532
rect 1326 2528 1330 2532
rect 1550 2528 1554 2532
rect 1686 2528 1690 2532
rect 1694 2528 1698 2532
rect 1718 2528 1722 2532
rect 1742 2528 1746 2532
rect 2158 2527 2162 2531
rect 2198 2528 2202 2532
rect 2214 2528 2218 2532
rect 2246 2528 2250 2532
rect 2486 2528 2490 2532
rect 2622 2528 2626 2532
rect 2630 2528 2634 2532
rect 2782 2528 2786 2532
rect 2790 2528 2794 2532
rect 3070 2528 3074 2532
rect 3198 2528 3202 2532
rect 3374 2528 3378 2532
rect 3430 2528 3434 2532
rect 3462 2528 3466 2532
rect 3806 2527 3810 2531
rect 3822 2528 3826 2532
rect 3886 2528 3890 2532
rect 3942 2528 3946 2532
rect 4038 2528 4042 2532
rect 4094 2528 4098 2532
rect 4494 2528 4498 2532
rect 4558 2528 4562 2532
rect 4734 2528 4738 2532
rect 4822 2528 4826 2532
rect 4910 2528 4914 2532
rect 5102 2528 5106 2532
rect 5190 2528 5194 2532
rect 5270 2528 5274 2532
rect 14 2518 18 2522
rect 30 2518 34 2522
rect 102 2518 106 2522
rect 198 2518 202 2522
rect 294 2518 298 2522
rect 510 2518 514 2522
rect 574 2518 578 2522
rect 1158 2518 1162 2522
rect 1166 2518 1170 2522
rect 2814 2518 2818 2522
rect 3054 2518 3058 2522
rect 3094 2518 3098 2522
rect 3358 2518 3362 2522
rect 3470 2518 3474 2522
rect 3830 2518 3834 2522
rect 3950 2518 3954 2522
rect 4022 2518 4026 2522
rect 4046 2518 4050 2522
rect 4190 2518 4194 2522
rect 4310 2518 4314 2522
rect 4430 2518 4434 2522
rect 4702 2518 4706 2522
rect 4726 2518 4730 2522
rect 4774 2518 4778 2522
rect 4814 2518 4818 2522
rect 4870 2518 4874 2522
rect 4918 2518 4922 2522
rect 4974 2518 4978 2522
rect 5038 2518 5042 2522
rect 5078 2518 5082 2522
rect 5166 2518 5170 2522
rect 5214 2518 5218 2522
rect 5262 2518 5266 2522
rect 5302 2518 5306 2522
rect 438 2508 442 2512
rect 526 2508 530 2512
rect 542 2508 546 2512
rect 622 2508 626 2512
rect 3430 2508 3434 2512
rect 3574 2508 3578 2512
rect 3886 2508 3890 2512
rect 4094 2508 4098 2512
rect 5190 2508 5194 2512
rect 5238 2508 5242 2512
rect 858 2503 862 2507
rect 865 2503 869 2507
rect 1874 2503 1878 2507
rect 1881 2503 1885 2507
rect 2906 2503 2910 2507
rect 2913 2503 2917 2507
rect 3930 2503 3934 2507
rect 3937 2503 3941 2507
rect 4954 2503 4958 2507
rect 4961 2503 4965 2507
rect 478 2498 482 2502
rect 1150 2498 1154 2502
rect 1350 2498 1354 2502
rect 3414 2498 3418 2502
rect 3470 2498 3474 2502
rect 3654 2498 3658 2502
rect 3774 2498 3778 2502
rect 4014 2498 4018 2502
rect 4942 2498 4946 2502
rect 5070 2498 5074 2502
rect 5294 2498 5298 2502
rect 38 2488 42 2492
rect 118 2488 122 2492
rect 142 2488 146 2492
rect 206 2488 210 2492
rect 246 2488 250 2492
rect 454 2488 458 2492
rect 518 2488 522 2492
rect 606 2488 610 2492
rect 646 2488 650 2492
rect 686 2488 690 2492
rect 734 2488 738 2492
rect 766 2488 770 2492
rect 790 2488 794 2492
rect 854 2488 858 2492
rect 910 2488 914 2492
rect 966 2488 970 2492
rect 1102 2488 1106 2492
rect 1174 2488 1178 2492
rect 1222 2488 1226 2492
rect 1254 2488 1258 2492
rect 1302 2488 1306 2492
rect 1334 2488 1338 2492
rect 1382 2488 1386 2492
rect 1542 2488 1546 2492
rect 1566 2488 1570 2492
rect 1598 2488 1602 2492
rect 1798 2488 1802 2492
rect 1822 2488 1826 2492
rect 1966 2488 1970 2492
rect 1974 2488 1978 2492
rect 2014 2488 2018 2492
rect 2038 2488 2042 2492
rect 2134 2488 2138 2492
rect 2158 2488 2162 2492
rect 2254 2488 2258 2492
rect 2382 2488 2386 2492
rect 2494 2488 2498 2492
rect 2550 2488 2554 2492
rect 2558 2488 2562 2492
rect 2742 2488 2746 2492
rect 2774 2488 2778 2492
rect 2886 2488 2890 2492
rect 2950 2488 2954 2492
rect 3054 2488 3058 2492
rect 3150 2488 3154 2492
rect 3246 2488 3250 2492
rect 3334 2488 3338 2492
rect 3462 2488 3466 2492
rect 3550 2488 3554 2492
rect 3598 2488 3602 2492
rect 3982 2488 3986 2492
rect 4086 2488 4090 2492
rect 4094 2488 4098 2492
rect 4110 2488 4114 2492
rect 4638 2488 4642 2492
rect 4854 2488 4858 2492
rect 4878 2488 4882 2492
rect 4910 2488 4914 2492
rect 5270 2488 5274 2492
rect 14 2479 18 2483
rect 30 2478 34 2482
rect 78 2478 82 2482
rect 94 2478 98 2482
rect 294 2478 298 2482
rect 318 2478 322 2482
rect 366 2478 370 2482
rect 742 2478 746 2482
rect 774 2478 778 2482
rect 814 2478 818 2482
rect 838 2478 842 2482
rect 958 2478 962 2482
rect 1150 2478 1154 2482
rect 1206 2478 1210 2482
rect 1246 2478 1250 2482
rect 1350 2478 1354 2482
rect 1518 2478 1522 2482
rect 1774 2478 1778 2482
rect 1934 2478 1938 2482
rect 2262 2478 2266 2482
rect 2750 2478 2754 2482
rect 3022 2478 3026 2482
rect 3262 2479 3266 2483
rect 3414 2478 3418 2482
rect 3470 2478 3474 2482
rect 3558 2478 3562 2482
rect 3654 2478 3658 2482
rect 3670 2478 3674 2482
rect 3942 2478 3946 2482
rect 3974 2478 3978 2482
rect 4014 2478 4018 2482
rect 4238 2478 4242 2482
rect 4422 2478 4426 2482
rect 4494 2478 4498 2482
rect 4510 2478 4514 2482
rect 4590 2478 4594 2482
rect 4606 2478 4610 2482
rect 4670 2478 4674 2482
rect 4694 2478 4698 2482
rect 4766 2478 4770 2482
rect 4782 2478 4786 2482
rect 4790 2478 4794 2482
rect 4814 2478 4818 2482
rect 4942 2478 4946 2482
rect 5142 2478 5146 2482
rect 5254 2479 5258 2483
rect 5294 2478 5298 2482
rect 46 2468 50 2472
rect 110 2468 114 2472
rect 126 2468 130 2472
rect 174 2468 178 2472
rect 214 2468 218 2472
rect 294 2468 298 2472
rect 326 2468 330 2472
rect 374 2468 378 2472
rect 6 2458 10 2462
rect 54 2458 58 2462
rect 78 2458 82 2462
rect 134 2458 138 2462
rect 158 2458 162 2462
rect 222 2458 226 2462
rect 246 2458 250 2462
rect 270 2458 274 2462
rect 302 2458 306 2462
rect 334 2458 338 2462
rect 366 2458 370 2462
rect 414 2458 418 2462
rect 486 2468 490 2472
rect 494 2468 498 2472
rect 542 2468 546 2472
rect 574 2468 578 2472
rect 622 2468 626 2472
rect 630 2468 634 2472
rect 726 2468 730 2472
rect 758 2468 762 2472
rect 902 2468 906 2472
rect 934 2468 938 2472
rect 1046 2468 1050 2472
rect 1062 2468 1066 2472
rect 1110 2468 1114 2472
rect 1134 2468 1138 2472
rect 1174 2468 1178 2472
rect 1214 2468 1218 2472
rect 1246 2468 1250 2472
rect 1294 2468 1298 2472
rect 1334 2468 1338 2472
rect 1358 2468 1362 2472
rect 1446 2468 1450 2472
rect 1526 2468 1530 2472
rect 526 2458 530 2462
rect 678 2458 682 2462
rect 702 2458 706 2462
rect 718 2458 722 2462
rect 750 2458 754 2462
rect 790 2458 794 2462
rect 862 2458 866 2462
rect 926 2458 930 2462
rect 1030 2459 1034 2463
rect 1126 2458 1130 2462
rect 1166 2458 1170 2462
rect 1214 2458 1218 2462
rect 1270 2458 1274 2462
rect 1318 2458 1322 2462
rect 1566 2458 1570 2462
rect 1606 2468 1610 2472
rect 1670 2468 1674 2472
rect 1726 2468 1730 2472
rect 1814 2468 1818 2472
rect 1990 2468 1994 2472
rect 1998 2468 2002 2472
rect 2022 2468 2026 2472
rect 2142 2468 2146 2472
rect 2158 2468 2162 2472
rect 2262 2468 2266 2472
rect 2286 2468 2290 2472
rect 2302 2468 2306 2472
rect 2414 2468 2418 2472
rect 2518 2468 2522 2472
rect 1742 2459 1746 2463
rect 1790 2458 1794 2462
rect 1854 2458 1858 2462
rect 1886 2459 1890 2463
rect 2070 2459 2074 2463
rect 2102 2458 2106 2462
rect 2198 2458 2202 2462
rect 2222 2458 2226 2462
rect 2318 2459 2322 2463
rect 2350 2458 2354 2462
rect 2430 2459 2434 2463
rect 2758 2468 2762 2472
rect 2782 2468 2786 2472
rect 2846 2468 2850 2472
rect 2854 2468 2858 2472
rect 2894 2468 2898 2472
rect 2974 2468 2978 2472
rect 3070 2468 3074 2472
rect 3166 2468 3170 2472
rect 3198 2468 3202 2472
rect 3278 2468 3282 2472
rect 3326 2468 3330 2472
rect 3334 2468 3338 2472
rect 3406 2468 3410 2472
rect 3438 2468 3442 2472
rect 3478 2468 3482 2472
rect 3534 2468 3538 2472
rect 3550 2468 3554 2472
rect 3574 2468 3578 2472
rect 3630 2468 3634 2472
rect 3782 2468 3786 2472
rect 3822 2468 3826 2472
rect 3918 2468 3922 2472
rect 3934 2468 3938 2472
rect 4006 2468 4010 2472
rect 4030 2468 4034 2472
rect 4094 2468 4098 2472
rect 4102 2468 4106 2472
rect 4150 2468 4154 2472
rect 4182 2468 4186 2472
rect 4214 2468 4218 2472
rect 4270 2468 4274 2472
rect 4310 2468 4314 2472
rect 4398 2468 4402 2472
rect 4430 2468 4434 2472
rect 4470 2468 4474 2472
rect 4486 2468 4490 2472
rect 4582 2468 4586 2472
rect 4606 2468 4610 2472
rect 4630 2468 4634 2472
rect 4662 2468 4666 2472
rect 4742 2468 4746 2472
rect 4766 2468 4770 2472
rect 4798 2468 4802 2472
rect 4870 2468 4874 2472
rect 4910 2468 4914 2472
rect 4934 2468 4938 2472
rect 4966 2468 4970 2472
rect 5022 2468 5026 2472
rect 5158 2468 5162 2472
rect 5182 2468 5186 2472
rect 5214 2468 5218 2472
rect 5286 2468 5290 2472
rect 86 2448 90 2452
rect 166 2448 170 2452
rect 190 2448 194 2452
rect 278 2448 282 2452
rect 398 2448 402 2452
rect 710 2448 714 2452
rect 782 2448 786 2452
rect 886 2448 890 2452
rect 902 2448 906 2452
rect 1142 2448 1146 2452
rect 1174 2448 1178 2452
rect 1238 2448 1242 2452
rect 1278 2448 1282 2452
rect 1574 2448 1578 2452
rect 1598 2448 1602 2452
rect 1798 2448 1802 2452
rect 1966 2448 1970 2452
rect 1974 2448 1978 2452
rect 2014 2448 2018 2452
rect 2038 2448 2042 2452
rect 2158 2448 2162 2452
rect 70 2438 74 2442
rect 150 2438 154 2442
rect 694 2438 698 2442
rect 798 2438 802 2442
rect 822 2438 826 2442
rect 942 2438 946 2442
rect 1206 2438 1210 2442
rect 1294 2438 1298 2442
rect 1558 2438 1562 2442
rect 1678 2438 1682 2442
rect 1790 2438 1794 2442
rect 2510 2438 2514 2442
rect 2622 2459 2626 2463
rect 2678 2459 2682 2463
rect 2710 2458 2714 2462
rect 2990 2459 2994 2463
rect 3086 2459 3090 2463
rect 3182 2459 3186 2463
rect 3270 2458 3274 2462
rect 3310 2458 3314 2462
rect 3334 2458 3338 2462
rect 3358 2458 3362 2462
rect 3366 2458 3370 2462
rect 3446 2458 3450 2462
rect 3518 2458 3522 2462
rect 3566 2458 3570 2462
rect 3582 2458 3586 2462
rect 3622 2458 3626 2462
rect 3638 2458 3642 2462
rect 3654 2458 3658 2462
rect 3686 2458 3690 2462
rect 3718 2458 3722 2462
rect 3734 2458 3738 2462
rect 3766 2458 3770 2462
rect 3798 2458 3802 2462
rect 3862 2458 3866 2462
rect 3886 2458 3890 2462
rect 3910 2458 3914 2462
rect 3958 2458 3962 2462
rect 3998 2458 4002 2462
rect 4038 2458 4042 2462
rect 4054 2458 4058 2462
rect 4118 2458 4122 2462
rect 4174 2458 4178 2462
rect 4206 2458 4210 2462
rect 4222 2458 4226 2462
rect 4238 2458 4242 2462
rect 4262 2458 4266 2462
rect 4278 2458 4282 2462
rect 4326 2459 4330 2463
rect 4534 2458 4538 2462
rect 4574 2458 4578 2462
rect 4590 2458 4594 2462
rect 4630 2458 4634 2462
rect 4670 2458 4674 2462
rect 4734 2458 4738 2462
rect 4750 2458 4754 2462
rect 4822 2458 4826 2462
rect 4838 2458 4842 2462
rect 5022 2458 5026 2462
rect 5062 2458 5066 2462
rect 5094 2458 5098 2462
rect 5126 2458 5130 2462
rect 5158 2458 5162 2462
rect 5174 2458 5178 2462
rect 5206 2458 5210 2462
rect 5238 2458 5242 2462
rect 5246 2458 5250 2462
rect 2526 2448 2530 2452
rect 2550 2448 2554 2452
rect 2870 2448 2874 2452
rect 3350 2448 3354 2452
rect 3526 2448 3530 2452
rect 3534 2448 3538 2452
rect 3606 2448 3610 2452
rect 3726 2448 3730 2452
rect 3758 2448 3762 2452
rect 3814 2448 3818 2452
rect 3870 2448 3874 2452
rect 3878 2448 3882 2452
rect 4006 2448 4010 2452
rect 4046 2448 4050 2452
rect 4078 2448 4082 2452
rect 4158 2448 4162 2452
rect 4190 2448 4194 2452
rect 4398 2448 4402 2452
rect 4454 2448 4458 2452
rect 4486 2448 4490 2452
rect 4510 2448 4514 2452
rect 4526 2448 4530 2452
rect 4558 2448 4562 2452
rect 4638 2448 4642 2452
rect 4718 2448 4722 2452
rect 4886 2448 4890 2452
rect 4894 2448 4898 2452
rect 5038 2448 5042 2452
rect 5070 2448 5074 2452
rect 5102 2448 5106 2452
rect 5134 2448 5138 2452
rect 5158 2448 5162 2452
rect 5190 2448 5194 2452
rect 2526 2438 2530 2442
rect 2574 2438 2578 2442
rect 3374 2438 3378 2442
rect 3390 2438 3394 2442
rect 3494 2438 3498 2442
rect 3510 2438 3514 2442
rect 3742 2438 3746 2442
rect 3886 2438 3890 2442
rect 4062 2438 4066 2442
rect 4206 2438 4210 2442
rect 4222 2438 4226 2442
rect 4526 2438 4530 2442
rect 4542 2438 4546 2442
rect 4750 2438 4754 2442
rect 4910 2438 4914 2442
rect 5054 2438 5058 2442
rect 5086 2438 5090 2442
rect 5118 2438 5122 2442
rect 1382 2428 1386 2432
rect 5094 2428 5098 2432
rect 350 2418 354 2422
rect 382 2418 386 2422
rect 830 2418 834 2422
rect 1126 2418 1130 2422
rect 1502 2418 1506 2422
rect 1662 2418 1666 2422
rect 1942 2418 1946 2422
rect 2950 2418 2954 2422
rect 3382 2418 3386 2422
rect 3518 2418 3522 2422
rect 3622 2418 3626 2422
rect 3750 2418 3754 2422
rect 3886 2418 3890 2422
rect 3934 2418 3938 2422
rect 4054 2418 4058 2422
rect 4174 2418 4178 2422
rect 4390 2418 4394 2422
rect 4550 2418 4554 2422
rect 4574 2418 4578 2422
rect 4686 2418 4690 2422
rect 4918 2418 4922 2422
rect 4990 2418 4994 2422
rect 5062 2418 5066 2422
rect 5110 2418 5114 2422
rect 5206 2418 5210 2422
rect 346 2403 350 2407
rect 353 2403 357 2407
rect 1370 2403 1374 2407
rect 1377 2403 1381 2407
rect 2394 2403 2398 2407
rect 2401 2403 2405 2407
rect 3418 2403 3422 2407
rect 3425 2403 3429 2407
rect 4442 2403 4446 2407
rect 4449 2403 4453 2407
rect 38 2388 42 2392
rect 86 2388 90 2392
rect 118 2388 122 2392
rect 198 2388 202 2392
rect 270 2388 274 2392
rect 310 2388 314 2392
rect 382 2388 386 2392
rect 494 2388 498 2392
rect 550 2388 554 2392
rect 638 2388 642 2392
rect 678 2388 682 2392
rect 774 2388 778 2392
rect 838 2388 842 2392
rect 998 2388 1002 2392
rect 1110 2388 1114 2392
rect 1286 2388 1290 2392
rect 1518 2388 1522 2392
rect 1558 2388 1562 2392
rect 1614 2388 1618 2392
rect 1710 2388 1714 2392
rect 1758 2388 1762 2392
rect 1782 2388 1786 2392
rect 1830 2388 1834 2392
rect 1926 2388 1930 2392
rect 1982 2388 1986 2392
rect 2006 2388 2010 2392
rect 2126 2388 2130 2392
rect 2166 2388 2170 2392
rect 2190 2388 2194 2392
rect 2246 2388 2250 2392
rect 2342 2388 2346 2392
rect 2606 2388 2610 2392
rect 2822 2388 2826 2392
rect 3454 2388 3458 2392
rect 3806 2388 3810 2392
rect 4046 2388 4050 2392
rect 4134 2388 4138 2392
rect 5182 2388 5186 2392
rect 1094 2378 1098 2382
rect 2990 2378 2994 2382
rect 4750 2378 4754 2382
rect 5214 2378 5218 2382
rect 30 2368 34 2372
rect 70 2368 74 2372
rect 110 2368 114 2372
rect 118 2368 122 2372
rect 190 2368 194 2372
rect 302 2368 306 2372
rect 414 2368 418 2372
rect 502 2368 506 2372
rect 590 2368 594 2372
rect 630 2368 634 2372
rect 662 2368 666 2372
rect 670 2368 674 2372
rect 710 2368 714 2372
rect 782 2368 786 2372
rect 1006 2368 1010 2372
rect 1030 2368 1034 2372
rect 1118 2368 1122 2372
rect 1190 2368 1194 2372
rect 1398 2368 1402 2372
rect 1702 2368 1706 2372
rect 1766 2368 1770 2372
rect 1798 2368 1802 2372
rect 1822 2368 1826 2372
rect 1966 2368 1970 2372
rect 1998 2368 2002 2372
rect 2006 2368 2010 2372
rect 2798 2368 2802 2372
rect 2814 2368 2818 2372
rect 2902 2368 2906 2372
rect 2966 2368 2970 2372
rect 3214 2368 3218 2372
rect 3238 2368 3242 2372
rect 3246 2368 3250 2372
rect 3366 2368 3370 2372
rect 3510 2368 3514 2372
rect 3958 2368 3962 2372
rect 3998 2368 4002 2372
rect 4054 2368 4058 2372
rect 4102 2368 4106 2372
rect 4246 2368 4250 2372
rect 4526 2368 4530 2372
rect 4542 2368 4546 2372
rect 4726 2368 4730 2372
rect 4758 2368 4762 2372
rect 4950 2368 4954 2372
rect 5014 2368 5018 2372
rect 5030 2368 5034 2372
rect 5070 2368 5074 2372
rect 5102 2368 5106 2372
rect 5126 2368 5130 2372
rect 14 2358 18 2362
rect 54 2358 58 2362
rect 174 2358 178 2362
rect 198 2358 202 2362
rect 286 2358 290 2362
rect 318 2358 322 2362
rect 454 2358 458 2362
rect 478 2358 482 2362
rect 486 2358 490 2362
rect 518 2358 522 2362
rect 614 2358 618 2362
rect 646 2358 650 2362
rect 654 2358 658 2362
rect 758 2358 762 2362
rect 766 2358 770 2362
rect 830 2358 834 2362
rect 998 2358 1002 2362
rect 1062 2358 1066 2362
rect 1086 2358 1090 2362
rect 1126 2358 1130 2362
rect 1670 2358 1674 2362
rect 1718 2358 1722 2362
rect 1742 2358 1746 2362
rect 1750 2358 1754 2362
rect 1838 2358 1842 2362
rect 1918 2358 1922 2362
rect 1958 2358 1962 2362
rect 2014 2358 2018 2362
rect 2366 2358 2370 2362
rect 2830 2358 2834 2362
rect 2870 2358 2874 2362
rect 2886 2358 2890 2362
rect 3046 2358 3050 2362
rect 3134 2358 3138 2362
rect 3198 2358 3202 2362
rect 3254 2358 3258 2362
rect 3262 2358 3266 2362
rect 3278 2358 3282 2362
rect 3310 2358 3314 2362
rect 3326 2358 3330 2362
rect 3342 2358 3346 2362
rect 3358 2358 3362 2362
rect 3382 2358 3386 2362
rect 3478 2358 3482 2362
rect 3518 2358 3522 2362
rect 3646 2358 3650 2362
rect 3694 2358 3698 2362
rect 3726 2358 3730 2362
rect 38 2348 42 2352
rect 86 2348 90 2352
rect 118 2348 122 2352
rect 158 2348 162 2352
rect 166 2348 170 2352
rect 198 2348 202 2352
rect 222 2348 226 2352
rect 238 2348 242 2352
rect 270 2348 274 2352
rect 310 2348 314 2352
rect 326 2348 330 2352
rect 438 2348 442 2352
rect 494 2348 498 2352
rect 638 2348 642 2352
rect 662 2348 666 2352
rect 694 2348 698 2352
rect 702 2348 706 2352
rect 742 2348 746 2352
rect 750 2348 754 2352
rect 774 2348 778 2352
rect 806 2348 810 2352
rect 822 2348 826 2352
rect 910 2347 914 2351
rect 950 2348 954 2352
rect 958 2348 962 2352
rect 974 2348 978 2352
rect 1006 2348 1010 2352
rect 1030 2348 1034 2352
rect 1126 2348 1130 2352
rect 1150 2348 1154 2352
rect 1166 2348 1170 2352
rect 1254 2347 1258 2351
rect 1342 2348 1346 2352
rect 1462 2347 1466 2351
rect 1494 2348 1498 2352
rect 1710 2348 1714 2352
rect 1766 2348 1770 2352
rect 1830 2348 1834 2352
rect 1846 2348 1850 2352
rect 1902 2348 1906 2352
rect 1918 2348 1922 2352
rect 1950 2348 1954 2352
rect 1966 2348 1970 2352
rect 2006 2348 2010 2352
rect 2030 2348 2034 2352
rect 94 2338 98 2342
rect 150 2338 154 2342
rect 214 2338 218 2342
rect 262 2338 266 2342
rect 334 2338 338 2342
rect 358 2338 362 2342
rect 390 2338 394 2342
rect 430 2338 434 2342
rect 534 2338 538 2342
rect 582 2338 586 2342
rect 686 2338 690 2342
rect 734 2338 738 2342
rect 798 2338 802 2342
rect 886 2338 890 2342
rect 926 2338 930 2342
rect 966 2338 970 2342
rect 1062 2338 1066 2342
rect 1078 2338 1082 2342
rect 1102 2338 1106 2342
rect 1158 2338 1162 2342
rect 1182 2338 1186 2342
rect 1270 2338 1274 2342
rect 1350 2338 1354 2342
rect 1478 2338 1482 2342
rect 1502 2338 1506 2342
rect 1574 2338 1578 2342
rect 1582 2338 1586 2342
rect 1630 2338 1634 2342
rect 1686 2338 1690 2342
rect 1726 2338 1730 2342
rect 1854 2338 1858 2342
rect 1886 2338 1890 2342
rect 1942 2338 1946 2342
rect 2062 2347 2066 2351
rect 2094 2348 2098 2352
rect 2214 2348 2218 2352
rect 2278 2347 2282 2351
rect 2302 2348 2306 2352
rect 2374 2348 2378 2352
rect 2414 2348 2418 2352
rect 2510 2348 2514 2352
rect 2542 2347 2546 2351
rect 2574 2348 2578 2352
rect 2638 2347 2642 2351
rect 2646 2348 2650 2352
rect 2670 2348 2674 2352
rect 2734 2347 2738 2351
rect 2766 2348 2770 2352
rect 2822 2348 2826 2352
rect 2878 2348 2882 2352
rect 2918 2348 2922 2352
rect 2998 2348 3002 2352
rect 3030 2348 3034 2352
rect 3054 2348 3058 2352
rect 3174 2348 3178 2352
rect 3190 2348 3194 2352
rect 3206 2348 3210 2352
rect 3246 2348 3250 2352
rect 3278 2348 3282 2352
rect 3326 2348 3330 2352
rect 3358 2348 3362 2352
rect 3518 2348 3522 2352
rect 3622 2348 3626 2352
rect 3662 2348 3666 2352
rect 3710 2348 3714 2352
rect 3910 2358 3914 2362
rect 3934 2358 3938 2362
rect 3974 2358 3978 2362
rect 4006 2358 4010 2362
rect 4070 2358 4074 2362
rect 4078 2358 4082 2362
rect 4094 2358 4098 2362
rect 4270 2358 4274 2362
rect 4310 2358 4314 2362
rect 4470 2358 4474 2362
rect 4510 2358 4514 2362
rect 4590 2358 4594 2362
rect 4742 2358 4746 2362
rect 4830 2358 4834 2362
rect 4862 2358 4866 2362
rect 4998 2358 5002 2362
rect 5046 2358 5050 2362
rect 5054 2358 5058 2362
rect 5086 2358 5090 2362
rect 5198 2358 5202 2362
rect 3782 2348 3786 2352
rect 3798 2348 3802 2352
rect 3822 2348 3826 2352
rect 3854 2348 3858 2352
rect 3966 2348 3970 2352
rect 3982 2348 3986 2352
rect 3998 2348 4002 2352
rect 4038 2348 4042 2352
rect 4062 2348 4066 2352
rect 4166 2348 4170 2352
rect 4206 2348 4210 2352
rect 4302 2348 4306 2352
rect 4326 2348 4330 2352
rect 4366 2348 4370 2352
rect 4398 2348 4402 2352
rect 4422 2348 4426 2352
rect 4502 2348 4506 2352
rect 4518 2348 4522 2352
rect 4590 2348 4594 2352
rect 4678 2348 4682 2352
rect 4710 2348 4714 2352
rect 4734 2348 4738 2352
rect 4766 2348 4770 2352
rect 4798 2348 4802 2352
rect 4814 2348 4818 2352
rect 4846 2348 4850 2352
rect 4878 2348 4882 2352
rect 4894 2348 4898 2352
rect 4910 2348 4914 2352
rect 4982 2348 4986 2352
rect 5038 2348 5042 2352
rect 5062 2348 5066 2352
rect 5094 2348 5098 2352
rect 5118 2348 5122 2352
rect 5134 2348 5138 2352
rect 5182 2348 5186 2352
rect 5214 2348 5218 2352
rect 5230 2348 5234 2352
rect 5254 2348 5258 2352
rect 5294 2348 5298 2352
rect 2182 2338 2186 2342
rect 2206 2338 2210 2342
rect 2230 2338 2234 2342
rect 2350 2338 2354 2342
rect 2478 2338 2482 2342
rect 2846 2338 2850 2342
rect 2926 2338 2930 2342
rect 2942 2338 2946 2342
rect 2966 2338 2970 2342
rect 2974 2340 2978 2344
rect 3014 2338 3018 2342
rect 3054 2338 3058 2342
rect 3070 2338 3074 2342
rect 3118 2338 3122 2342
rect 3158 2338 3162 2342
rect 3166 2338 3170 2342
rect 14 2328 18 2332
rect 54 2328 58 2332
rect 254 2328 258 2332
rect 374 2328 378 2332
rect 414 2328 418 2332
rect 518 2328 522 2332
rect 590 2328 594 2332
rect 614 2328 618 2332
rect 726 2328 730 2332
rect 950 2328 954 2332
rect 982 2328 986 2332
rect 1038 2328 1042 2332
rect 1054 2328 1058 2332
rect 1518 2328 1522 2332
rect 1734 2328 1738 2332
rect 1790 2328 1794 2332
rect 1798 2328 1802 2332
rect 1870 2328 1874 2332
rect 1926 2328 1930 2332
rect 2030 2328 2034 2332
rect 2190 2328 2194 2332
rect 2222 2328 2226 2332
rect 2358 2328 2362 2332
rect 2382 2327 2386 2331
rect 2950 2328 2954 2332
rect 3014 2328 3018 2332
rect 3062 2328 3066 2332
rect 3142 2328 3146 2332
rect 3246 2338 3250 2342
rect 3286 2338 3290 2342
rect 3294 2338 3298 2342
rect 3318 2338 3322 2342
rect 3398 2338 3402 2342
rect 3422 2338 3426 2342
rect 3470 2338 3474 2342
rect 3494 2338 3498 2342
rect 3534 2338 3538 2342
rect 3582 2338 3586 2342
rect 3590 2338 3594 2342
rect 3638 2338 3642 2342
rect 3678 2338 3682 2342
rect 3718 2338 3722 2342
rect 3750 2338 3754 2342
rect 3774 2338 3778 2342
rect 3782 2338 3786 2342
rect 3894 2340 3898 2344
rect 3910 2338 3914 2342
rect 3942 2338 3946 2342
rect 4030 2338 4034 2342
rect 4078 2338 4082 2342
rect 4118 2338 4122 2342
rect 4270 2338 4274 2342
rect 4334 2338 4338 2342
rect 4446 2338 4450 2342
rect 4494 2338 4498 2342
rect 4558 2338 4562 2342
rect 4574 2338 4578 2342
rect 4598 2338 4602 2342
rect 4654 2338 4658 2342
rect 4670 2338 4674 2342
rect 4822 2338 4826 2342
rect 4894 2338 4898 2342
rect 4910 2338 4914 2342
rect 4918 2338 4922 2342
rect 4998 2338 5002 2342
rect 5014 2338 5018 2342
rect 5070 2338 5074 2342
rect 5190 2338 5194 2342
rect 5222 2338 5226 2342
rect 5310 2338 5314 2342
rect 3190 2328 3194 2332
rect 3206 2328 3210 2332
rect 3390 2328 3394 2332
rect 3518 2328 3522 2332
rect 3758 2328 3762 2332
rect 3830 2328 3834 2332
rect 3870 2328 3874 2332
rect 4014 2328 4018 2332
rect 4126 2328 4130 2332
rect 4142 2328 4146 2332
rect 4198 2328 4202 2332
rect 4286 2328 4290 2332
rect 4302 2328 4306 2332
rect 4350 2328 4354 2332
rect 4478 2328 4482 2332
rect 4566 2328 4570 2332
rect 4654 2328 4658 2332
rect 4686 2328 4690 2332
rect 4790 2328 4794 2332
rect 4910 2328 4914 2332
rect 4942 2328 4946 2332
rect 5094 2328 5098 2332
rect 5150 2328 5154 2332
rect 246 2318 250 2322
rect 398 2318 402 2322
rect 478 2318 482 2322
rect 574 2318 578 2322
rect 1862 2318 1866 2322
rect 2494 2318 2498 2322
rect 2702 2318 2706 2322
rect 2878 2318 2882 2322
rect 3102 2318 3106 2322
rect 3134 2318 3138 2322
rect 3150 2318 3154 2322
rect 5238 2327 5242 2331
rect 5262 2327 5266 2331
rect 3302 2318 3306 2322
rect 3366 2318 3370 2322
rect 3478 2318 3482 2322
rect 3550 2318 3554 2322
rect 3606 2318 3610 2322
rect 3734 2318 3738 2322
rect 3766 2318 3770 2322
rect 3878 2318 3882 2322
rect 3910 2318 3914 2322
rect 4022 2318 4026 2322
rect 4310 2318 4314 2322
rect 4398 2318 4402 2322
rect 4446 2318 4450 2322
rect 4470 2318 4474 2322
rect 4486 2318 4490 2322
rect 4534 2318 4538 2322
rect 4590 2318 4594 2322
rect 4606 2318 4610 2322
rect 4662 2318 4666 2322
rect 4694 2318 4698 2322
rect 4830 2318 4834 2322
rect 4894 2318 4898 2322
rect 4950 2318 4954 2322
rect 5006 2318 5010 2322
rect 5278 2318 5282 2322
rect 766 2308 770 2312
rect 982 2308 986 2312
rect 1054 2308 1058 2312
rect 3014 2308 3018 2312
rect 4286 2308 4290 2312
rect 4566 2308 4570 2312
rect 4910 2308 4914 2312
rect 858 2303 862 2307
rect 865 2303 869 2307
rect 1874 2303 1878 2307
rect 1881 2303 1885 2307
rect 2906 2303 2910 2307
rect 2913 2303 2917 2307
rect 3930 2303 3934 2307
rect 3937 2303 3941 2307
rect 4954 2303 4958 2307
rect 4961 2303 4965 2307
rect 2966 2298 2970 2302
rect 14 2288 18 2292
rect 22 2288 26 2292
rect 118 2288 122 2292
rect 142 2288 146 2292
rect 190 2288 194 2292
rect 270 2288 274 2292
rect 350 2288 354 2292
rect 390 2288 394 2292
rect 414 2288 418 2292
rect 502 2288 506 2292
rect 630 2288 634 2292
rect 670 2288 674 2292
rect 790 2288 794 2292
rect 894 2288 898 2292
rect 966 2288 970 2292
rect 1014 2288 1018 2292
rect 1038 2288 1042 2292
rect 1134 2288 1138 2292
rect 1318 2288 1322 2292
rect 1390 2288 1394 2292
rect 1478 2288 1482 2292
rect 1518 2288 1522 2292
rect 1622 2288 1626 2292
rect 1734 2288 1738 2292
rect 1926 2288 1930 2292
rect 1966 2288 1970 2292
rect 2078 2288 2082 2292
rect 2126 2288 2130 2292
rect 2150 2288 2154 2292
rect 2182 2288 2186 2292
rect 2254 2288 2258 2292
rect 2398 2288 2402 2292
rect 2622 2288 2626 2292
rect 2846 2288 2850 2292
rect 2854 2288 2858 2292
rect 2870 2288 2874 2292
rect 3358 2288 3362 2292
rect 3382 2288 3386 2292
rect 3406 2288 3410 2292
rect 3526 2288 3530 2292
rect 3542 2288 3546 2292
rect 3550 2288 3554 2292
rect 3886 2288 3890 2292
rect 4134 2288 4138 2292
rect 4182 2288 4186 2292
rect 4246 2288 4250 2292
rect 4542 2288 4546 2292
rect 4566 2288 4570 2292
rect 4814 2288 4818 2292
rect 5022 2288 5026 2292
rect 5166 2288 5170 2292
rect 5214 2288 5218 2292
rect 5302 2288 5306 2292
rect 182 2278 186 2282
rect 222 2278 226 2282
rect 318 2278 322 2282
rect 406 2278 410 2282
rect 542 2278 546 2282
rect 710 2278 714 2282
rect 726 2279 730 2283
rect 750 2279 754 2283
rect 1166 2278 1170 2282
rect 1198 2278 1202 2282
rect 6 2268 10 2272
rect 54 2268 58 2272
rect 110 2268 114 2272
rect 158 2268 162 2272
rect 206 2268 210 2272
rect 230 2268 234 2272
rect 238 2268 242 2272
rect 286 2268 290 2272
rect 334 2268 338 2272
rect 374 2268 378 2272
rect 382 2268 386 2272
rect 430 2268 434 2272
rect 486 2268 490 2272
rect 534 2268 538 2272
rect 566 2268 570 2272
rect 646 2268 650 2272
rect 654 2268 658 2272
rect 886 2268 890 2272
rect 918 2268 922 2272
rect 926 2268 930 2272
rect 974 2268 978 2272
rect 982 2268 986 2272
rect 998 2268 1002 2272
rect 1030 2268 1034 2272
rect 1118 2268 1122 2272
rect 1278 2268 1282 2272
rect 1286 2268 1290 2272
rect 1334 2268 1338 2272
rect 1342 2268 1346 2272
rect 1358 2268 1362 2272
rect 1414 2268 1418 2272
rect 1462 2268 1466 2272
rect 1590 2278 1594 2282
rect 1606 2278 1610 2282
rect 1798 2278 1802 2282
rect 1878 2278 1882 2282
rect 1950 2278 1954 2282
rect 2086 2278 2090 2282
rect 2134 2278 2138 2282
rect 2286 2278 2290 2282
rect 2366 2278 2370 2282
rect 2566 2279 2570 2283
rect 2878 2278 2882 2282
rect 2886 2278 2890 2282
rect 2926 2278 2930 2282
rect 2966 2278 2970 2282
rect 3006 2278 3010 2282
rect 3102 2278 3106 2282
rect 3310 2278 3314 2282
rect 3414 2278 3418 2282
rect 3766 2278 3770 2282
rect 3854 2278 3858 2282
rect 3870 2278 3874 2282
rect 3878 2278 3882 2282
rect 3934 2278 3938 2282
rect 4110 2278 4114 2282
rect 4534 2278 4538 2282
rect 4558 2278 4562 2282
rect 4638 2278 4642 2282
rect 4702 2278 4706 2282
rect 4734 2278 4738 2282
rect 5014 2278 5018 2282
rect 5142 2278 5146 2282
rect 5198 2278 5202 2282
rect 5206 2278 5210 2282
rect 1510 2268 1514 2272
rect 1534 2268 1538 2272
rect 1574 2268 1578 2272
rect 1590 2268 1594 2272
rect 1630 2268 1634 2272
rect 1718 2268 1722 2272
rect 1846 2268 1850 2272
rect 1862 2268 1866 2272
rect 1886 2268 1890 2272
rect 1918 2268 1922 2272
rect 1942 2268 1946 2272
rect 2006 2268 2010 2272
rect 2054 2268 2058 2272
rect 2070 2268 2074 2272
rect 2094 2268 2098 2272
rect 2110 2268 2114 2272
rect 2158 2268 2162 2272
rect 2198 2268 2202 2272
rect 2246 2268 2250 2272
rect 2358 2268 2362 2272
rect 2462 2268 2466 2272
rect 2518 2268 2522 2272
rect 2590 2268 2594 2272
rect 2638 2268 2642 2272
rect 2686 2268 2690 2272
rect 2790 2268 2794 2272
rect 2854 2268 2858 2272
rect 2894 2268 2898 2272
rect 2966 2268 2970 2272
rect 2982 2268 2986 2272
rect 3014 2268 3018 2272
rect 3094 2268 3098 2272
rect 3118 2268 3122 2272
rect 3134 2268 3138 2272
rect 3166 2268 3170 2272
rect 3214 2268 3218 2272
rect 3222 2268 3226 2272
rect 3270 2268 3274 2272
rect 3326 2268 3330 2272
rect 3366 2268 3370 2272
rect 3382 2268 3386 2272
rect 3398 2268 3402 2272
rect 3534 2268 3538 2272
rect 3582 2268 3586 2272
rect 3590 2268 3594 2272
rect 3638 2268 3642 2272
rect 3662 2268 3666 2272
rect 3670 2268 3674 2272
rect 3734 2268 3738 2272
rect 3766 2268 3770 2272
rect 3782 2268 3786 2272
rect 3798 2268 3802 2272
rect 3814 2268 3818 2272
rect 62 2258 66 2262
rect 102 2258 106 2262
rect 166 2258 170 2262
rect 310 2258 314 2262
rect 366 2258 370 2262
rect 422 2258 426 2262
rect 446 2258 450 2262
rect 478 2258 482 2262
rect 558 2258 562 2262
rect 598 2258 602 2262
rect 734 2258 738 2262
rect 758 2258 762 2262
rect 766 2258 770 2262
rect 854 2259 858 2263
rect 990 2258 994 2262
rect 1102 2259 1106 2263
rect 1198 2259 1202 2263
rect 1278 2258 1282 2262
rect 1390 2258 1394 2262
rect 1542 2258 1546 2262
rect 1558 2258 1562 2262
rect 1702 2259 1706 2263
rect 1798 2259 1802 2263
rect 1870 2258 1874 2262
rect 1998 2258 2002 2262
rect 2062 2258 2066 2262
rect 2102 2258 2106 2262
rect 2182 2258 2186 2262
rect 2230 2258 2234 2262
rect 2294 2258 2298 2262
rect 2454 2258 2458 2262
rect 2678 2258 2682 2262
rect 2790 2258 2794 2262
rect 2902 2258 2906 2262
rect 2950 2258 2954 2262
rect 2990 2258 2994 2262
rect 3086 2258 3090 2262
rect 3094 2258 3098 2262
rect 3126 2258 3130 2262
rect 3142 2258 3146 2262
rect 3294 2258 3298 2262
rect 3334 2258 3338 2262
rect 3390 2258 3394 2262
rect 3470 2258 3474 2262
rect 3494 2258 3498 2262
rect 3678 2258 3682 2262
rect 3718 2258 3722 2262
rect 3742 2258 3746 2262
rect 3750 2258 3754 2262
rect 3790 2258 3794 2262
rect 3854 2268 3858 2272
rect 3894 2268 3898 2272
rect 3926 2268 3930 2272
rect 3990 2268 3994 2272
rect 4006 2268 4010 2272
rect 4078 2268 4082 2272
rect 4094 2268 4098 2272
rect 4158 2268 4162 2272
rect 4166 2268 4170 2272
rect 4214 2268 4218 2272
rect 4222 2268 4226 2272
rect 4270 2268 4274 2272
rect 4310 2268 4314 2272
rect 4326 2268 4330 2272
rect 4342 2268 4346 2272
rect 4422 2268 4426 2272
rect 4438 2268 4442 2272
rect 4470 2268 4474 2272
rect 4510 2268 4514 2272
rect 4526 2268 4530 2272
rect 4574 2268 4578 2272
rect 4614 2268 4618 2272
rect 4638 2268 4642 2272
rect 4662 2268 4666 2272
rect 4678 2268 4682 2272
rect 4686 2268 4690 2272
rect 4718 2268 4722 2272
rect 4742 2268 4746 2272
rect 4758 2268 4762 2272
rect 4798 2268 4802 2272
rect 4846 2268 4850 2272
rect 4854 2268 4858 2272
rect 4902 2268 4906 2272
rect 4910 2268 4914 2272
rect 4958 2268 4962 2272
rect 4982 2268 4986 2272
rect 5030 2268 5034 2272
rect 5046 2268 5050 2272
rect 5054 2268 5058 2272
rect 5086 2268 5090 2272
rect 5142 2268 5146 2272
rect 5150 2268 5154 2272
rect 5230 2268 5234 2272
rect 5246 2268 5250 2272
rect 3838 2258 3842 2262
rect 3902 2258 3906 2262
rect 3974 2258 3978 2262
rect 4030 2258 4034 2262
rect 4046 2258 4050 2262
rect 4086 2258 4090 2262
rect 4110 2258 4114 2262
rect 4126 2258 4130 2262
rect 4150 2258 4154 2262
rect 4294 2258 4298 2262
rect 4342 2258 4346 2262
rect 4374 2258 4378 2262
rect 4398 2258 4402 2262
rect 4414 2258 4418 2262
rect 4486 2258 4490 2262
rect 4510 2258 4514 2262
rect 4550 2258 4554 2262
rect 4574 2258 4578 2262
rect 4590 2258 4594 2262
rect 4606 2258 4610 2262
rect 4622 2258 4626 2262
rect 4774 2258 4778 2262
rect 4886 2258 4890 2262
rect 4918 2258 4922 2262
rect 4934 2258 4938 2262
rect 4990 2258 4994 2262
rect 5134 2258 5138 2262
rect 5174 2258 5178 2262
rect 5190 2258 5194 2262
rect 5222 2258 5226 2262
rect 190 2248 194 2252
rect 214 2248 218 2252
rect 398 2248 402 2252
rect 590 2248 594 2252
rect 678 2248 682 2252
rect 886 2248 890 2252
rect 1006 2248 1010 2252
rect 1014 2248 1018 2252
rect 1382 2248 1386 2252
rect 1470 2248 1474 2252
rect 1526 2248 1530 2252
rect 1558 2248 1562 2252
rect 1590 2248 1594 2252
rect 1614 2248 1618 2252
rect 1830 2248 1834 2252
rect 1902 2248 1906 2252
rect 1974 2248 1978 2252
rect 2142 2248 2146 2252
rect 2190 2248 2194 2252
rect 2254 2248 2258 2252
rect 2398 2248 2402 2252
rect 2870 2248 2874 2252
rect 3070 2248 3074 2252
rect 3158 2248 3162 2252
rect 3358 2248 3362 2252
rect 3382 2248 3386 2252
rect 3646 2248 3650 2252
rect 3694 2248 3698 2252
rect 3726 2248 3730 2252
rect 3758 2248 3762 2252
rect 3798 2248 3802 2252
rect 3950 2248 3954 2252
rect 3982 2248 3986 2252
rect 3990 2248 3994 2252
rect 4014 2248 4018 2252
rect 4046 2248 4050 2252
rect 4102 2248 4106 2252
rect 4302 2248 4306 2252
rect 4310 2248 4314 2252
rect 4334 2248 4338 2252
rect 4366 2248 4370 2252
rect 4446 2248 4450 2252
rect 4502 2248 4506 2252
rect 4510 2248 4514 2252
rect 4598 2248 4602 2252
rect 4758 2248 4762 2252
rect 4766 2248 4770 2252
rect 4934 2248 4938 2252
rect 4942 2248 4946 2252
rect 5006 2248 5010 2252
rect 5062 2248 5066 2252
rect 5254 2248 5258 2252
rect 5278 2268 5282 2272
rect 5286 2258 5290 2262
rect 5278 2248 5282 2252
rect 558 2238 562 2242
rect 1398 2238 1402 2242
rect 1430 2238 1434 2242
rect 1638 2238 1642 2242
rect 2022 2238 2026 2242
rect 2174 2238 2178 2242
rect 2510 2238 2514 2242
rect 3286 2238 3290 2242
rect 3710 2238 3714 2242
rect 3966 2238 3970 2242
rect 3974 2238 3978 2242
rect 4022 2238 4026 2242
rect 4030 2238 4034 2242
rect 4286 2238 4290 2242
rect 4350 2238 4354 2242
rect 4382 2238 4386 2242
rect 4398 2238 4402 2242
rect 2750 2228 2754 2232
rect 3838 2228 3842 2232
rect 4294 2228 4298 2232
rect 1542 2218 1546 2222
rect 1886 2218 1890 2222
rect 2150 2218 2154 2222
rect 2302 2218 2306 2222
rect 2574 2218 2578 2222
rect 2926 2218 2930 2222
rect 3046 2218 3050 2222
rect 3142 2218 3146 2222
rect 3182 2218 3186 2222
rect 3254 2218 3258 2222
rect 3294 2218 3298 2222
rect 3614 2218 3618 2222
rect 3678 2218 3682 2222
rect 3718 2218 3722 2222
rect 3830 2218 3834 2222
rect 3910 2218 3914 2222
rect 4182 2218 4186 2222
rect 4254 2218 4258 2222
rect 4734 2218 4738 2222
rect 4790 2218 4794 2222
rect 4918 2218 4922 2222
rect 4990 2218 4994 2222
rect 5078 2218 5082 2222
rect 5262 2218 5266 2222
rect 346 2203 350 2207
rect 353 2203 357 2207
rect 1370 2203 1374 2207
rect 1377 2203 1381 2207
rect 2394 2203 2398 2207
rect 2401 2203 2405 2207
rect 3418 2203 3422 2207
rect 3425 2203 3429 2207
rect 4442 2203 4446 2207
rect 4449 2203 4453 2207
rect 326 2188 330 2192
rect 366 2188 370 2192
rect 566 2188 570 2192
rect 886 2188 890 2192
rect 1190 2188 1194 2192
rect 1438 2188 1442 2192
rect 1566 2188 1570 2192
rect 1718 2188 1722 2192
rect 1766 2188 1770 2192
rect 1958 2188 1962 2192
rect 2070 2188 2074 2192
rect 2078 2188 2082 2192
rect 2134 2188 2138 2192
rect 2174 2188 2178 2192
rect 2222 2188 2226 2192
rect 2390 2188 2394 2192
rect 2502 2188 2506 2192
rect 2862 2188 2866 2192
rect 2942 2188 2946 2192
rect 2998 2188 3002 2192
rect 3070 2188 3074 2192
rect 3126 2188 3130 2192
rect 3654 2188 3658 2192
rect 3694 2188 3698 2192
rect 3742 2188 3746 2192
rect 4270 2188 4274 2192
rect 4366 2188 4370 2192
rect 4430 2188 4434 2192
rect 4574 2188 4578 2192
rect 5142 2188 5146 2192
rect 5206 2188 5210 2192
rect 5278 2188 5282 2192
rect 5302 2188 5306 2192
rect 454 2178 458 2182
rect 486 2178 490 2182
rect 662 2178 666 2182
rect 766 2178 770 2182
rect 4222 2178 4226 2182
rect 4238 2178 4242 2182
rect 54 2168 58 2172
rect 150 2168 154 2172
rect 174 2168 178 2172
rect 462 2168 466 2172
rect 670 2168 674 2172
rect 1542 2168 1546 2172
rect 1646 2168 1650 2172
rect 1662 2168 1666 2172
rect 1966 2168 1970 2172
rect 2126 2168 2130 2172
rect 2870 2168 2874 2172
rect 3078 2168 3082 2172
rect 3134 2168 3138 2172
rect 3198 2168 3202 2172
rect 3270 2168 3274 2172
rect 3366 2168 3370 2172
rect 3574 2168 3578 2172
rect 4214 2168 4218 2172
rect 4246 2168 4250 2172
rect 4278 2168 4282 2172
rect 4582 2168 4586 2172
rect 4590 2168 4594 2172
rect 4622 2168 4626 2172
rect 4662 2168 4666 2172
rect 4950 2168 4954 2172
rect 4990 2168 4994 2172
rect 5030 2168 5034 2172
rect 5214 2168 5218 2172
rect 70 2158 74 2162
rect 134 2158 138 2162
rect 158 2158 162 2162
rect 182 2158 186 2162
rect 390 2158 394 2162
rect 422 2158 426 2162
rect 438 2158 442 2162
rect 582 2158 586 2162
rect 614 2158 618 2162
rect 654 2158 658 2162
rect 686 2158 690 2162
rect 6 2148 10 2152
rect 46 2148 50 2152
rect 102 2148 106 2152
rect 142 2148 146 2152
rect 198 2148 202 2152
rect 262 2148 266 2152
rect 366 2148 370 2152
rect 382 2148 386 2152
rect 406 2148 410 2152
rect 454 2148 458 2152
rect 526 2148 530 2152
rect 534 2148 538 2152
rect 598 2148 602 2152
rect 614 2148 618 2152
rect 638 2148 642 2152
rect 662 2148 666 2152
rect 742 2158 746 2162
rect 758 2158 762 2162
rect 878 2158 882 2162
rect 926 2158 930 2162
rect 1294 2158 1298 2162
rect 1558 2158 1562 2162
rect 1646 2158 1650 2162
rect 1694 2158 1698 2162
rect 1702 2158 1706 2162
rect 1886 2158 1890 2162
rect 1950 2158 1954 2162
rect 2158 2158 2162 2162
rect 2214 2158 2218 2162
rect 2430 2158 2434 2162
rect 2446 2158 2450 2162
rect 2574 2158 2578 2162
rect 2694 2158 2698 2162
rect 2766 2158 2770 2162
rect 2854 2158 2858 2162
rect 2902 2158 2906 2162
rect 3054 2158 3058 2162
rect 3062 2158 3066 2162
rect 3150 2158 3154 2162
rect 3206 2158 3210 2162
rect 3238 2158 3242 2162
rect 3382 2158 3386 2162
rect 3406 2158 3410 2162
rect 3934 2158 3938 2162
rect 3982 2158 3986 2162
rect 4030 2158 4034 2162
rect 4038 2158 4042 2162
rect 4078 2158 4082 2162
rect 4230 2158 4234 2162
rect 4262 2158 4266 2162
rect 4294 2158 4298 2162
rect 4310 2158 4314 2162
rect 4542 2158 4546 2162
rect 4550 2158 4554 2162
rect 4654 2158 4658 2162
rect 4830 2158 4834 2162
rect 4894 2158 4898 2162
rect 4934 2158 4938 2162
rect 5014 2158 5018 2162
rect 5070 2158 5074 2162
rect 5102 2158 5106 2162
rect 5118 2158 5122 2162
rect 5198 2158 5202 2162
rect 5230 2158 5234 2162
rect 5286 2158 5290 2162
rect 726 2148 730 2152
rect 782 2148 786 2152
rect 806 2148 810 2152
rect 822 2148 826 2152
rect 854 2148 858 2152
rect 910 2148 914 2152
rect 918 2148 922 2152
rect 942 2148 946 2152
rect 950 2148 954 2152
rect 990 2148 994 2152
rect 54 2138 58 2142
rect 70 2138 74 2142
rect 94 2138 98 2142
rect 110 2138 114 2142
rect 190 2138 194 2142
rect 206 2138 210 2142
rect 270 2138 274 2142
rect 294 2138 298 2142
rect 342 2138 346 2142
rect 1062 2147 1066 2151
rect 1158 2147 1162 2151
rect 1222 2148 1226 2152
rect 1254 2147 1258 2151
rect 1318 2148 1322 2152
rect 1398 2148 1402 2152
rect 1494 2148 1498 2152
rect 1542 2148 1546 2152
rect 1614 2148 1618 2152
rect 1654 2148 1658 2152
rect 1702 2148 1706 2152
rect 1718 2148 1722 2152
rect 1734 2148 1738 2152
rect 1814 2148 1818 2152
rect 1838 2147 1842 2151
rect 1894 2148 1898 2152
rect 1942 2148 1946 2152
rect 1958 2148 1962 2152
rect 2006 2147 2010 2151
rect 2118 2148 2122 2152
rect 2142 2148 2146 2152
rect 2174 2148 2178 2152
rect 2182 2148 2186 2152
rect 2270 2148 2274 2152
rect 2326 2148 2330 2152
rect 2358 2147 2362 2151
rect 2414 2148 2418 2152
rect 2446 2148 2450 2152
rect 2470 2148 2474 2152
rect 2558 2148 2562 2152
rect 2566 2148 2570 2152
rect 2614 2148 2618 2152
rect 2670 2148 2674 2152
rect 2806 2148 2810 2152
rect 2830 2148 2834 2152
rect 2846 2148 2850 2152
rect 2862 2148 2866 2152
rect 3038 2148 3042 2152
rect 3070 2148 3074 2152
rect 3118 2148 3122 2152
rect 3142 2148 3146 2152
rect 3158 2148 3162 2152
rect 3206 2148 3210 2152
rect 3222 2148 3226 2152
rect 3262 2148 3266 2152
rect 3270 2148 3274 2152
rect 3286 2148 3290 2152
rect 3310 2148 3314 2152
rect 3326 2148 3330 2152
rect 3374 2148 3378 2152
rect 3598 2148 3602 2152
rect 3806 2148 3810 2152
rect 3918 2148 3922 2152
rect 3990 2148 3994 2152
rect 4150 2148 4154 2152
rect 4238 2148 4242 2152
rect 4270 2148 4274 2152
rect 4406 2148 4410 2152
rect 4446 2148 4450 2152
rect 4590 2148 4594 2152
rect 4606 2148 4610 2152
rect 4614 2148 4618 2152
rect 4710 2148 4714 2152
rect 4758 2148 4762 2152
rect 4766 2148 4770 2152
rect 4798 2148 4802 2152
rect 4822 2148 4826 2152
rect 4846 2148 4850 2152
rect 4862 2148 4866 2152
rect 4926 2148 4930 2152
rect 4958 2148 4962 2152
rect 4998 2148 5002 2152
rect 5086 2148 5090 2152
rect 5102 2148 5106 2152
rect 5190 2148 5194 2152
rect 5206 2148 5210 2152
rect 5246 2148 5250 2152
rect 5302 2148 5306 2152
rect 414 2138 418 2142
rect 438 2138 442 2142
rect 478 2138 482 2142
rect 534 2138 538 2142
rect 558 2138 562 2142
rect 590 2138 594 2142
rect 606 2138 610 2142
rect 646 2138 650 2142
rect 686 2138 690 2142
rect 702 2138 706 2142
rect 726 2138 730 2142
rect 878 2138 882 2142
rect 894 2138 898 2142
rect 902 2138 906 2142
rect 1078 2138 1082 2142
rect 1150 2138 1154 2142
rect 1422 2138 1426 2142
rect 1502 2138 1506 2142
rect 1534 2138 1538 2142
rect 1590 2138 1594 2142
rect 1678 2138 1682 2142
rect 1878 2138 1882 2142
rect 1910 2138 1914 2142
rect 1934 2138 1938 2142
rect 2270 2138 2274 2142
rect 2286 2138 2290 2142
rect 2398 2138 2402 2142
rect 2422 2138 2426 2142
rect 2462 2138 2466 2142
rect 2534 2138 2538 2142
rect 2590 2138 2594 2142
rect 2598 2138 2602 2142
rect 2646 2138 2650 2142
rect 2678 2138 2682 2142
rect 2694 2138 2698 2142
rect 2718 2138 2722 2142
rect 2782 2138 2786 2142
rect 2814 2138 2818 2142
rect 2838 2138 2842 2142
rect 2886 2138 2890 2142
rect 2926 2138 2930 2142
rect 2974 2138 2978 2142
rect 2982 2138 2986 2142
rect 3030 2138 3034 2142
rect 3038 2138 3042 2142
rect 3102 2138 3106 2142
rect 3166 2138 3170 2142
rect 3230 2138 3234 2142
rect 3246 2138 3250 2142
rect 3262 2138 3266 2142
rect 3326 2138 3330 2142
rect 3334 2138 3338 2142
rect 3406 2138 3410 2142
rect 3478 2138 3482 2142
rect 3486 2138 3490 2142
rect 3534 2138 3538 2142
rect 3622 2138 3626 2142
rect 3670 2138 3674 2142
rect 3726 2138 3730 2142
rect 3798 2138 3802 2142
rect 3854 2138 3858 2142
rect 3902 2138 3906 2142
rect 3958 2138 3962 2142
rect 3998 2138 4002 2142
rect 4030 2138 4034 2142
rect 4062 2138 4066 2142
rect 4094 2138 4098 2142
rect 4294 2138 4298 2142
rect 4310 2138 4314 2142
rect 4334 2138 4338 2142
rect 4350 2138 4354 2142
rect 4414 2138 4418 2142
rect 4462 2138 4466 2142
rect 4470 2138 4474 2142
rect 4526 2138 4530 2142
rect 4550 2138 4554 2142
rect 4566 2138 4570 2142
rect 4638 2138 4642 2142
rect 4654 2138 4658 2142
rect 4678 2138 4682 2142
rect 4734 2138 4738 2142
rect 4758 2138 4762 2142
rect 4774 2138 4778 2142
rect 4862 2138 4866 2142
rect 4870 2138 4874 2142
rect 4886 2138 4890 2142
rect 4910 2138 4914 2142
rect 4958 2138 4962 2142
rect 5014 2138 5018 2142
rect 5030 2138 5034 2142
rect 5054 2138 5058 2142
rect 5086 2138 5090 2142
rect 5094 2138 5098 2142
rect 5182 2138 5186 2142
rect 5254 2138 5258 2142
rect 5310 2138 5314 2142
rect 30 2128 34 2132
rect 118 2128 122 2132
rect 126 2128 130 2132
rect 174 2128 178 2132
rect 214 2128 218 2132
rect 278 2128 282 2132
rect 542 2128 546 2132
rect 710 2128 714 2132
rect 774 2128 778 2132
rect 782 2128 786 2132
rect 798 2128 802 2132
rect 838 2128 842 2132
rect 862 2128 866 2132
rect 942 2128 946 2132
rect 1294 2128 1298 2132
rect 1310 2127 1314 2131
rect 1574 2128 1578 2132
rect 1582 2128 1586 2132
rect 1638 2128 1642 2132
rect 1654 2128 1658 2132
rect 1750 2128 1754 2132
rect 1758 2128 1762 2132
rect 1918 2128 1922 2132
rect 2006 2128 2010 2132
rect 2086 2128 2090 2132
rect 2094 2128 2098 2132
rect 2142 2128 2146 2132
rect 2206 2128 2210 2132
rect 2246 2128 2250 2132
rect 2254 2128 2258 2132
rect 2478 2128 2482 2132
rect 2726 2128 2730 2132
rect 2822 2128 2826 2132
rect 3094 2128 3098 2132
rect 3190 2128 3194 2132
rect 3286 2128 3290 2132
rect 3350 2128 3354 2132
rect 3822 2128 3826 2132
rect 3846 2128 3850 2132
rect 4014 2128 4018 2132
rect 4086 2128 4090 2132
rect 4142 2128 4146 2132
rect 4342 2128 4346 2132
rect 4430 2128 4434 2132
rect 4550 2128 4554 2132
rect 4686 2128 4690 2132
rect 4694 2128 4698 2132
rect 4702 2128 4706 2132
rect 4750 2128 4754 2132
rect 4806 2128 4810 2132
rect 4894 2128 4898 2132
rect 5062 2128 5066 2132
rect 5126 2128 5130 2132
rect 5166 2128 5170 2132
rect 5238 2128 5242 2132
rect 5254 2128 5258 2132
rect 86 2118 90 2122
rect 230 2118 234 2122
rect 246 2118 250 2122
rect 494 2118 498 2122
rect 726 2118 730 2122
rect 910 2118 914 2122
rect 998 2118 1002 2122
rect 1094 2118 1098 2122
rect 1342 2118 1346 2122
rect 1774 2118 1778 2122
rect 2262 2118 2266 2122
rect 2294 2118 2298 2122
rect 2542 2118 2546 2122
rect 2574 2118 2578 2122
rect 2590 2118 2594 2122
rect 2686 2118 2690 2122
rect 2790 2118 2794 2122
rect 2918 2118 2922 2122
rect 3038 2118 3042 2122
rect 3174 2118 3178 2122
rect 3326 2118 3330 2122
rect 3342 2118 3346 2122
rect 3374 2118 3378 2122
rect 3422 2118 3426 2122
rect 3446 2118 3450 2122
rect 3526 2118 3530 2122
rect 3838 2118 3842 2122
rect 3870 2118 3874 2122
rect 3982 2118 3986 2122
rect 4006 2118 4010 2122
rect 4110 2118 4114 2122
rect 4486 2118 4490 2122
rect 4726 2118 4730 2122
rect 4862 2118 4866 2122
rect 4990 2118 4994 2122
rect 5070 2118 5074 2122
rect 5286 2118 5290 2122
rect 30 2108 34 2112
rect 542 2108 546 2112
rect 710 2108 714 2112
rect 742 2108 746 2112
rect 838 2108 842 2112
rect 3094 2108 3098 2112
rect 3286 2108 3290 2112
rect 4638 2108 4642 2112
rect 4686 2108 4690 2112
rect 4806 2108 4810 2112
rect 858 2103 862 2107
rect 865 2103 869 2107
rect 1874 2103 1878 2107
rect 1881 2103 1885 2107
rect 2906 2103 2910 2107
rect 2913 2103 2917 2107
rect 3930 2103 3934 2107
rect 3937 2103 3941 2107
rect 4954 2103 4958 2107
rect 4961 2103 4965 2107
rect 374 2098 378 2102
rect 982 2098 986 2102
rect 1846 2098 1850 2102
rect 2598 2098 2602 2102
rect 3030 2098 3034 2102
rect 3558 2098 3562 2102
rect 3694 2098 3698 2102
rect 14 2088 18 2092
rect 30 2088 34 2092
rect 46 2088 50 2092
rect 70 2088 74 2092
rect 110 2088 114 2092
rect 238 2088 242 2092
rect 342 2088 346 2092
rect 406 2088 410 2092
rect 430 2088 434 2092
rect 478 2088 482 2092
rect 566 2088 570 2092
rect 622 2088 626 2092
rect 718 2088 722 2092
rect 766 2088 770 2092
rect 830 2088 834 2092
rect 846 2088 850 2092
rect 886 2088 890 2092
rect 1046 2088 1050 2092
rect 1086 2088 1090 2092
rect 1278 2088 1282 2092
rect 1422 2088 1426 2092
rect 1470 2088 1474 2092
rect 1486 2088 1490 2092
rect 1502 2088 1506 2092
rect 1590 2088 1594 2092
rect 1702 2088 1706 2092
rect 1766 2088 1770 2092
rect 1902 2088 1906 2092
rect 1918 2088 1922 2092
rect 1958 2088 1962 2092
rect 1998 2088 2002 2092
rect 2062 2088 2066 2092
rect 2110 2088 2114 2092
rect 2134 2088 2138 2092
rect 2190 2088 2194 2092
rect 2294 2088 2298 2092
rect 2670 2088 2674 2092
rect 2838 2088 2842 2092
rect 2854 2088 2858 2092
rect 2894 2088 2898 2092
rect 3046 2088 3050 2092
rect 3382 2088 3386 2092
rect 3502 2088 3506 2092
rect 3646 2088 3650 2092
rect 3718 2088 3722 2092
rect 3910 2088 3914 2092
rect 4014 2088 4018 2092
rect 4206 2088 4210 2092
rect 4286 2088 4290 2092
rect 4470 2088 4474 2092
rect 4526 2088 4530 2092
rect 4622 2088 4626 2092
rect 4670 2088 4674 2092
rect 4678 2088 4682 2092
rect 4750 2088 4754 2092
rect 4790 2088 4794 2092
rect 4846 2088 4850 2092
rect 4902 2088 4906 2092
rect 4926 2088 4930 2092
rect 5086 2088 5090 2092
rect 78 2078 82 2082
rect 190 2078 194 2082
rect 254 2078 258 2082
rect 318 2078 322 2082
rect 350 2078 354 2082
rect 374 2078 378 2082
rect 470 2078 474 2082
rect 582 2078 586 2082
rect 982 2078 986 2082
rect 1014 2078 1018 2082
rect 1078 2078 1082 2082
rect 1150 2078 1154 2082
rect 1310 2078 1314 2082
rect 1494 2078 1498 2082
rect 1566 2078 1570 2082
rect 1582 2078 1586 2082
rect 1654 2078 1658 2082
rect 1726 2078 1730 2082
rect 1742 2078 1746 2082
rect 1758 2078 1762 2082
rect 1846 2078 1850 2082
rect 1910 2078 1914 2082
rect 1926 2078 1930 2082
rect 1990 2078 1994 2082
rect 2070 2078 2074 2082
rect 2094 2078 2098 2082
rect 2302 2078 2306 2082
rect 6 2068 10 2072
rect 38 2068 42 2072
rect 86 2068 90 2072
rect 134 2068 138 2072
rect 150 2068 154 2072
rect 2478 2078 2482 2082
rect 2630 2078 2634 2082
rect 2726 2078 2730 2082
rect 2806 2078 2810 2082
rect 3094 2078 3098 2082
rect 3174 2078 3178 2082
rect 3206 2078 3210 2082
rect 3390 2078 3394 2082
rect 3750 2078 3754 2082
rect 3990 2078 3994 2082
rect 4054 2078 4058 2082
rect 4142 2078 4146 2082
rect 4254 2078 4258 2082
rect 4886 2078 4890 2082
rect 5030 2078 5034 2082
rect 5110 2078 5114 2082
rect 5286 2079 5290 2083
rect 246 2068 250 2072
rect 270 2068 274 2072
rect 414 2068 418 2072
rect 438 2068 442 2072
rect 454 2068 458 2072
rect 502 2068 506 2072
rect 542 2068 546 2072
rect 590 2068 594 2072
rect 638 2068 642 2072
rect 694 2068 698 2072
rect 742 2068 746 2072
rect 798 2068 802 2072
rect 806 2068 810 2072
rect 854 2068 858 2072
rect 878 2068 882 2072
rect 926 2068 930 2072
rect 1006 2068 1010 2072
rect 1030 2068 1034 2072
rect 1038 2068 1042 2072
rect 1054 2068 1058 2072
rect 1070 2068 1074 2072
rect 1214 2068 1218 2072
rect 1262 2068 1266 2072
rect 1358 2068 1362 2072
rect 1390 2068 1394 2072
rect 1438 2068 1442 2072
rect 1446 2068 1450 2072
rect 14 2058 18 2062
rect 30 2058 34 2062
rect 62 2058 66 2062
rect 158 2058 162 2062
rect 174 2058 178 2062
rect 206 2058 210 2062
rect 278 2058 282 2062
rect 294 2058 298 2062
rect 318 2058 322 2062
rect 398 2058 402 2062
rect 446 2058 450 2062
rect 494 2058 498 2062
rect 510 2058 514 2062
rect 526 2058 530 2062
rect 646 2058 650 2062
rect 694 2058 698 2062
rect 894 2058 898 2062
rect 950 2058 954 2062
rect 966 2058 970 2062
rect 1030 2058 1034 2062
rect 1118 2058 1122 2062
rect 1150 2059 1154 2063
rect 1246 2059 1250 2063
rect 1334 2058 1338 2062
rect 1454 2058 1458 2062
rect 1478 2058 1482 2062
rect 1518 2058 1522 2062
rect 1558 2068 1562 2072
rect 1694 2068 1698 2072
rect 1766 2068 1770 2072
rect 1838 2068 1842 2072
rect 1854 2068 1858 2072
rect 1886 2068 1890 2072
rect 1934 2068 1938 2072
rect 1982 2068 1986 2072
rect 2006 2068 2010 2072
rect 2038 2068 2042 2072
rect 1550 2058 1554 2062
rect 1566 2058 1570 2062
rect 1654 2059 1658 2063
rect 1686 2058 1690 2062
rect 1782 2058 1786 2062
rect 1798 2058 1802 2062
rect 2086 2068 2090 2072
rect 2118 2068 2122 2072
rect 2126 2068 2130 2072
rect 2174 2068 2178 2072
rect 2198 2068 2202 2072
rect 2318 2068 2322 2072
rect 2326 2068 2330 2072
rect 2366 2068 2370 2072
rect 2494 2068 2498 2072
rect 2582 2068 2586 2072
rect 2646 2068 2650 2072
rect 2230 2059 2234 2063
rect 2766 2068 2770 2072
rect 2798 2068 2802 2072
rect 2830 2068 2834 2072
rect 2870 2068 2874 2072
rect 2878 2068 2882 2072
rect 2926 2068 2930 2072
rect 3030 2068 3034 2072
rect 3070 2068 3074 2072
rect 3102 2068 3106 2072
rect 3134 2068 3138 2072
rect 3238 2068 3242 2072
rect 3342 2068 3346 2072
rect 3358 2068 3362 2072
rect 3374 2068 3378 2072
rect 3422 2068 3426 2072
rect 3438 2068 3442 2072
rect 3462 2068 3466 2072
rect 3470 2068 3474 2072
rect 3518 2068 3522 2072
rect 3566 2068 3570 2072
rect 3574 2068 3578 2072
rect 3622 2068 3626 2072
rect 3630 2068 3634 2072
rect 3678 2068 3682 2072
rect 3686 2068 3690 2072
rect 3734 2068 3738 2072
rect 3806 2068 3810 2072
rect 3822 2068 3826 2072
rect 3990 2068 3994 2072
rect 3998 2068 4002 2072
rect 4054 2068 4058 2072
rect 4070 2068 4074 2072
rect 4206 2068 4210 2072
rect 4222 2068 4226 2072
rect 4246 2068 4250 2072
rect 4278 2068 4282 2072
rect 4494 2068 4498 2072
rect 4542 2068 4546 2072
rect 4550 2068 4554 2072
rect 4598 2068 4602 2072
rect 4654 2068 4658 2072
rect 4662 2068 4666 2072
rect 4710 2068 4714 2072
rect 4718 2068 4722 2072
rect 4766 2068 4770 2072
rect 4774 2068 4778 2072
rect 4822 2068 4826 2072
rect 4830 2068 4834 2072
rect 4902 2068 4906 2072
rect 4958 2068 4962 2072
rect 5006 2068 5010 2072
rect 5046 2068 5050 2072
rect 2262 2058 2266 2062
rect 2374 2058 2378 2062
rect 2422 2058 2426 2062
rect 2454 2058 2458 2062
rect 2486 2058 2490 2062
rect 2502 2058 2506 2062
rect 2526 2058 2530 2062
rect 2542 2058 2546 2062
rect 2558 2058 2562 2062
rect 2566 2058 2570 2062
rect 2606 2058 2610 2062
rect 2654 2058 2658 2062
rect 2670 2058 2674 2062
rect 2710 2058 2714 2062
rect 2742 2058 2746 2062
rect 2758 2058 2762 2062
rect 2782 2058 2786 2062
rect 2790 2058 2794 2062
rect 2822 2058 2826 2062
rect 2982 2058 2986 2062
rect 3006 2058 3010 2062
rect 3062 2058 3066 2062
rect 3078 2058 3082 2062
rect 3110 2058 3114 2062
rect 3142 2058 3146 2062
rect 3158 2058 3162 2062
rect 3190 2058 3194 2062
rect 3222 2058 3226 2062
rect 3254 2058 3258 2062
rect 3294 2058 3298 2062
rect 3318 2058 3322 2062
rect 3342 2058 3346 2062
rect 3366 2058 3370 2062
rect 3414 2058 3418 2062
rect 3478 2058 3482 2062
rect 3502 2058 3506 2062
rect 3558 2058 3562 2062
rect 3590 2058 3594 2062
rect 3838 2059 3842 2063
rect 4086 2058 4090 2062
rect 4110 2058 4114 2062
rect 4222 2058 4226 2062
rect 4318 2058 4322 2062
rect 4342 2058 4346 2062
rect 4406 2059 4410 2063
rect 4910 2058 4914 2062
rect 4982 2058 4986 2062
rect 5070 2058 5074 2062
rect 5118 2068 5122 2072
rect 5166 2068 5170 2072
rect 5174 2068 5178 2072
rect 5222 2068 5226 2072
rect 5094 2058 5098 2062
rect 5110 2058 5114 2062
rect 5230 2058 5234 2062
rect 5254 2058 5258 2062
rect 5278 2058 5282 2062
rect 30 2048 34 2052
rect 166 2048 170 2052
rect 222 2048 226 2052
rect 230 2048 234 2052
rect 286 2048 290 2052
rect 422 2048 426 2052
rect 510 2048 514 2052
rect 566 2048 570 2052
rect 582 2048 586 2052
rect 1062 2048 1066 2052
rect 1502 2048 1506 2052
rect 1766 2048 1770 2052
rect 1782 2048 1786 2052
rect 1854 2048 1858 2052
rect 2022 2048 2026 2052
rect 2102 2048 2106 2052
rect 2182 2048 2186 2052
rect 2334 2048 2338 2052
rect 2390 2048 2394 2052
rect 2446 2048 2450 2052
rect 2534 2048 2538 2052
rect 2598 2048 2602 2052
rect 2662 2048 2666 2052
rect 2774 2048 2778 2052
rect 2846 2048 2850 2052
rect 2854 2048 2858 2052
rect 3126 2048 3130 2052
rect 3214 2048 3218 2052
rect 3246 2048 3250 2052
rect 3302 2048 3306 2052
rect 3358 2048 3362 2052
rect 3398 2048 3402 2052
rect 3446 2048 3450 2052
rect 3542 2048 3546 2052
rect 4094 2048 4098 2052
rect 4102 2048 4106 2052
rect 4142 2048 4146 2052
rect 4206 2048 4210 2052
rect 4278 2048 4282 2052
rect 5022 2048 5026 2052
rect 5078 2048 5082 2052
rect 5094 2048 5098 2052
rect 150 2038 154 2042
rect 166 2038 170 2042
rect 302 2038 306 2042
rect 398 2038 402 2042
rect 1006 2038 1010 2042
rect 1182 2038 1186 2042
rect 1742 2038 1746 2042
rect 1806 2038 1810 2042
rect 1822 2038 1826 2042
rect 2430 2038 2434 2042
rect 2462 2038 2466 2042
rect 2518 2038 2522 2042
rect 2614 2038 2618 2042
rect 2670 2038 2674 2042
rect 2678 2038 2682 2042
rect 2702 2038 2706 2042
rect 3110 2038 3114 2042
rect 3174 2038 3178 2042
rect 3198 2038 3202 2042
rect 3222 2038 3226 2042
rect 3262 2038 3266 2042
rect 3286 2038 3290 2042
rect 3326 2038 3330 2042
rect 3558 2038 3562 2042
rect 4110 2038 4114 2042
rect 4166 2038 4170 2042
rect 4566 2038 4570 2042
rect 5190 2038 5194 2042
rect 470 2028 474 2032
rect 2142 2028 2146 2032
rect 3294 2028 3298 2032
rect 3414 2028 3418 2032
rect 3534 2028 3538 2032
rect 5054 2028 5058 2032
rect 14 2018 18 2022
rect 206 2018 210 2022
rect 254 2018 258 2022
rect 294 2018 298 2022
rect 934 2018 938 2022
rect 1718 2018 1722 2022
rect 1734 2018 1738 2022
rect 1814 2018 1818 2022
rect 1918 2018 1922 2022
rect 2310 2018 2314 2022
rect 2350 2018 2354 2022
rect 2374 2018 2378 2022
rect 2422 2018 2426 2022
rect 2470 2018 2474 2022
rect 2510 2018 2514 2022
rect 2606 2018 2610 2022
rect 2630 2018 2634 2022
rect 2694 2018 2698 2022
rect 2950 2018 2954 2022
rect 3254 2018 3258 2022
rect 3750 2018 3754 2022
rect 3934 2018 3938 2022
rect 4110 2018 4114 2022
rect 5014 2018 5018 2022
rect 346 2003 350 2007
rect 353 2003 357 2007
rect 1370 2003 1374 2007
rect 1377 2003 1381 2007
rect 2394 2003 2398 2007
rect 2401 2003 2405 2007
rect 3418 2003 3422 2007
rect 3425 2003 3429 2007
rect 4442 2003 4446 2007
rect 4449 2003 4453 2007
rect 174 1988 178 1992
rect 398 1988 402 1992
rect 470 1988 474 1992
rect 646 1988 650 1992
rect 758 1988 762 1992
rect 1142 1988 1146 1992
rect 1278 1988 1282 1992
rect 1358 1988 1362 1992
rect 1478 1988 1482 1992
rect 1502 1988 1506 1992
rect 1582 1988 1586 1992
rect 1622 1988 1626 1992
rect 1806 1988 1810 1992
rect 1926 1988 1930 1992
rect 2030 1988 2034 1992
rect 2798 1988 2802 1992
rect 2870 1988 2874 1992
rect 2894 1988 2898 1992
rect 3150 1988 3154 1992
rect 3366 1988 3370 1992
rect 3750 1988 3754 1992
rect 4118 1988 4122 1992
rect 4166 1988 4170 1992
rect 4206 1988 4210 1992
rect 4950 1988 4954 1992
rect 5006 1988 5010 1992
rect 5038 1988 5042 1992
rect 5078 1988 5082 1992
rect 5174 1988 5178 1992
rect 5254 1988 5258 1992
rect 5262 1988 5266 1992
rect 38 1978 42 1982
rect 1422 1978 1426 1982
rect 1774 1978 1778 1982
rect 2270 1978 2274 1982
rect 2606 1978 2610 1982
rect 6 1968 10 1972
rect 30 1968 34 1972
rect 222 1968 226 1972
rect 246 1968 250 1972
rect 262 1968 266 1972
rect 462 1968 466 1972
rect 534 1968 538 1972
rect 574 1968 578 1972
rect 998 1968 1002 1972
rect 1062 1968 1066 1972
rect 1110 1968 1114 1972
rect 1158 1968 1162 1972
rect 1574 1968 1578 1972
rect 1830 1968 1834 1972
rect 1838 1968 1842 1972
rect 2022 1968 2026 1972
rect 2054 1968 2058 1972
rect 2262 1968 2266 1972
rect 3142 1968 3146 1972
rect 3406 1968 3410 1972
rect 4006 1968 4010 1972
rect 4318 1968 4322 1972
rect 5270 1968 5274 1972
rect 46 1958 50 1962
rect 134 1958 138 1962
rect 214 1958 218 1962
rect 262 1958 266 1962
rect 358 1958 362 1962
rect 446 1958 450 1962
rect 478 1958 482 1962
rect 518 1958 522 1962
rect 582 1958 586 1962
rect 630 1958 634 1962
rect 638 1958 642 1962
rect 854 1958 858 1962
rect 870 1958 874 1962
rect 926 1958 930 1962
rect 982 1958 986 1962
rect 1046 1958 1050 1962
rect 1062 1958 1066 1962
rect 1294 1958 1298 1962
rect 1558 1958 1562 1962
rect 1590 1958 1594 1962
rect 38 1948 42 1952
rect 62 1948 66 1952
rect 78 1948 82 1952
rect 86 1948 90 1952
rect 102 1948 106 1952
rect 254 1948 258 1952
rect 294 1948 298 1952
rect 302 1948 306 1952
rect 318 1948 322 1952
rect 342 1948 346 1952
rect 374 1948 378 1952
rect 390 1948 394 1952
rect 470 1948 474 1952
rect 518 1948 522 1952
rect 566 1948 570 1952
rect 598 1948 602 1952
rect 614 1948 618 1952
rect 638 1948 642 1952
rect 70 1938 74 1942
rect 110 1938 114 1942
rect 190 1938 194 1942
rect 214 1938 218 1942
rect 286 1938 290 1942
rect 310 1938 314 1942
rect 326 1938 330 1942
rect 382 1938 386 1942
rect 390 1938 394 1942
rect 494 1938 498 1942
rect 510 1938 514 1942
rect 534 1938 538 1942
rect 598 1938 602 1942
rect 726 1947 730 1951
rect 774 1948 778 1952
rect 822 1948 826 1952
rect 838 1948 842 1952
rect 886 1948 890 1952
rect 910 1948 914 1952
rect 926 1948 930 1952
rect 974 1948 978 1952
rect 990 1948 994 1952
rect 1014 1948 1018 1952
rect 1030 1948 1034 1952
rect 1670 1957 1674 1961
rect 1742 1958 1746 1962
rect 1846 1958 1850 1962
rect 1870 1958 1874 1962
rect 1894 1958 1898 1962
rect 2038 1958 2042 1962
rect 2070 1958 2074 1962
rect 2094 1958 2098 1962
rect 2102 1958 2106 1962
rect 2134 1958 2138 1962
rect 2278 1958 2282 1962
rect 2310 1958 2314 1962
rect 2582 1958 2586 1962
rect 2782 1958 2786 1962
rect 2886 1958 2890 1962
rect 3126 1958 3130 1962
rect 3286 1958 3290 1962
rect 3350 1958 3354 1962
rect 4046 1958 4050 1962
rect 4078 1958 4082 1962
rect 4086 1958 4090 1962
rect 4126 1958 4130 1962
rect 1086 1948 1090 1952
rect 1102 1948 1106 1952
rect 1110 1948 1114 1952
rect 1126 1948 1130 1952
rect 654 1938 658 1942
rect 742 1938 746 1942
rect 782 1938 786 1942
rect 830 1938 834 1942
rect 902 1938 906 1942
rect 918 1938 922 1942
rect 942 1938 946 1942
rect 966 1938 970 1942
rect 1038 1938 1042 1942
rect 1222 1947 1226 1951
rect 1254 1948 1258 1952
rect 1278 1948 1282 1952
rect 1302 1948 1306 1952
rect 1318 1948 1322 1952
rect 1350 1948 1354 1952
rect 1542 1948 1546 1952
rect 1558 1948 1562 1952
rect 1582 1948 1586 1952
rect 1598 1948 1602 1952
rect 1686 1948 1690 1952
rect 1726 1948 1730 1952
rect 1750 1948 1754 1952
rect 1766 1948 1770 1952
rect 1790 1948 1794 1952
rect 1838 1948 1842 1952
rect 1910 1948 1914 1952
rect 1958 1948 1962 1952
rect 2030 1948 2034 1952
rect 2062 1948 2066 1952
rect 2118 1948 2122 1952
rect 2142 1948 2146 1952
rect 2150 1948 2154 1952
rect 2166 1948 2170 1952
rect 2214 1948 2218 1952
rect 2222 1948 2226 1952
rect 2270 1948 2274 1952
rect 2294 1948 2298 1952
rect 2350 1948 2354 1952
rect 2454 1948 2458 1952
rect 2462 1948 2466 1952
rect 2638 1948 2642 1952
rect 1134 1938 1138 1942
rect 1238 1938 1242 1942
rect 1270 1938 1274 1942
rect 1310 1938 1314 1942
rect 1326 1938 1330 1942
rect 1390 1938 1394 1942
rect 1438 1938 1442 1942
rect 1446 1938 1450 1942
rect 1494 1938 1498 1942
rect 1518 1938 1522 1942
rect 1534 1938 1538 1942
rect 1598 1938 1602 1942
rect 1654 1938 1658 1942
rect 1718 1938 1722 1942
rect 1750 1938 1754 1942
rect 1798 1938 1802 1942
rect 1854 1938 1858 1942
rect 1902 1938 1906 1942
rect 1918 1938 1922 1942
rect 1942 1938 1946 1942
rect 2006 1938 2010 1942
rect 2062 1938 2066 1942
rect 2078 1938 2082 1942
rect 2126 1938 2130 1942
rect 2158 1938 2162 1942
rect 2174 1938 2178 1942
rect 2190 1938 2194 1942
rect 2230 1938 2234 1942
rect 2286 1938 2290 1942
rect 2302 1938 2306 1942
rect 2334 1938 2338 1942
rect 2350 1938 2354 1942
rect 2726 1947 2730 1951
rect 2758 1948 2762 1952
rect 2798 1948 2802 1952
rect 2814 1948 2818 1952
rect 3022 1947 3026 1951
rect 3134 1948 3138 1952
rect 3158 1948 3162 1952
rect 3222 1948 3226 1952
rect 3246 1948 3250 1952
rect 3262 1948 3266 1952
rect 3310 1948 3314 1952
rect 3334 1948 3338 1952
rect 3358 1948 3362 1952
rect 3374 1948 3378 1952
rect 3454 1948 3458 1952
rect 2366 1938 2370 1942
rect 2446 1938 2450 1942
rect 2462 1938 2466 1942
rect 2478 1938 2482 1942
rect 2534 1938 2538 1942
rect 2566 1938 2570 1942
rect 2590 1938 2594 1942
rect 2638 1938 2642 1942
rect 2718 1938 2722 1942
rect 2806 1938 2810 1942
rect 2830 1938 2834 1942
rect 2854 1940 2858 1944
rect 2862 1938 2866 1942
rect 2942 1938 2946 1942
rect 2990 1938 2994 1942
rect 3030 1938 3034 1942
rect 3102 1938 3106 1942
rect 3118 1938 3122 1942
rect 3166 1938 3170 1942
rect 3198 1938 3202 1942
rect 3230 1938 3234 1942
rect 3254 1938 3258 1942
rect 3302 1938 3306 1942
rect 3318 1938 3322 1942
rect 3326 1938 3330 1942
rect 3382 1938 3386 1942
rect 3502 1948 3506 1952
rect 3630 1948 3634 1952
rect 3654 1948 3658 1952
rect 3742 1948 3746 1952
rect 3790 1948 3794 1952
rect 3870 1947 3874 1951
rect 3902 1948 3906 1952
rect 3974 1948 3978 1952
rect 4046 1948 4050 1952
rect 4110 1948 4114 1952
rect 3486 1938 3490 1942
rect 3534 1938 3538 1942
rect 3542 1938 3546 1942
rect 3694 1938 3698 1942
rect 3742 1938 3746 1942
rect 3974 1938 3978 1942
rect 4022 1938 4026 1942
rect 4030 1938 4034 1942
rect 4062 1938 4066 1942
rect 4270 1947 4274 1951
rect 4414 1948 4418 1952
rect 4486 1948 4490 1952
rect 4510 1958 4514 1962
rect 4838 1958 4842 1962
rect 5046 1958 5050 1962
rect 5206 1958 5210 1962
rect 5286 1958 5290 1962
rect 4622 1948 4626 1952
rect 4886 1947 4890 1951
rect 4918 1948 4922 1952
rect 5110 1947 5114 1951
rect 5142 1948 5146 1952
rect 5198 1948 5202 1952
rect 5270 1948 5274 1952
rect 4110 1938 4114 1942
rect 4126 1938 4130 1942
rect 4182 1938 4186 1942
rect 4190 1938 4194 1942
rect 4238 1938 4242 1942
rect 4254 1938 4258 1942
rect 4382 1938 4386 1942
rect 4406 1938 4410 1942
rect 4446 1938 4450 1942
rect 4510 1938 4514 1942
rect 4534 1940 4538 1944
rect 4550 1938 4554 1942
rect 4598 1938 4602 1942
rect 4630 1938 4634 1942
rect 4638 1938 4642 1942
rect 4686 1938 4690 1942
rect 4694 1938 4698 1942
rect 4742 1938 4746 1942
rect 4798 1938 4802 1942
rect 4806 1938 4810 1942
rect 4854 1938 4858 1942
rect 4974 1938 4978 1942
rect 5030 1938 5034 1942
rect 5062 1938 5066 1942
rect 5094 1938 5098 1942
rect 5222 1938 5226 1942
rect 5238 1940 5242 1944
rect 14 1928 18 1932
rect 54 1928 58 1932
rect 86 1928 90 1932
rect 222 1928 226 1932
rect 270 1928 274 1932
rect 430 1928 434 1932
rect 438 1928 442 1932
rect 550 1928 554 1932
rect 598 1928 602 1932
rect 726 1928 730 1932
rect 854 1928 858 1932
rect 1078 1928 1082 1932
rect 1086 1928 1090 1932
rect 1150 1928 1154 1932
rect 1262 1928 1266 1932
rect 1326 1928 1330 1932
rect 1342 1928 1346 1932
rect 1366 1928 1370 1932
rect 1502 1928 1506 1932
rect 1702 1928 1706 1932
rect 1750 1928 1754 1932
rect 1814 1928 1818 1932
rect 1926 1928 1930 1932
rect 2182 1928 2186 1932
rect 2190 1928 2194 1932
rect 2198 1928 2202 1932
rect 2238 1928 2242 1932
rect 2246 1928 2250 1932
rect 2318 1928 2322 1932
rect 2358 1928 2362 1932
rect 2430 1928 2434 1932
rect 2478 1928 2482 1932
rect 2814 1928 2818 1932
rect 2830 1928 2834 1932
rect 2878 1928 2882 1932
rect 2934 1928 2938 1932
rect 3094 1928 3098 1932
rect 3182 1928 3186 1932
rect 3190 1928 3194 1932
rect 3214 1928 3218 1932
rect 3254 1928 3258 1932
rect 3286 1928 3290 1932
rect 3398 1928 3402 1932
rect 3478 1928 3482 1932
rect 3622 1928 3626 1932
rect 4054 1928 4058 1932
rect 4342 1928 4346 1932
rect 4350 1928 4354 1932
rect 4398 1928 4402 1932
rect 4470 1928 4474 1932
rect 5054 1928 5058 1932
rect 238 1918 242 1922
rect 662 1918 666 1922
rect 806 1918 810 1922
rect 958 1918 962 1922
rect 998 1918 1002 1922
rect 1294 1918 1298 1922
rect 1862 1918 1866 1922
rect 1974 1918 1978 1922
rect 2086 1918 2090 1922
rect 2102 1918 2106 1922
rect 2326 1918 2330 1922
rect 2366 1918 2370 1922
rect 2438 1918 2442 1922
rect 2502 1918 2506 1922
rect 2574 1918 2578 1922
rect 2598 1918 2602 1922
rect 2958 1918 2962 1922
rect 3086 1918 3090 1922
rect 3350 1918 3354 1922
rect 3390 1918 3394 1922
rect 3518 1918 3522 1922
rect 3574 1918 3578 1922
rect 3686 1918 3690 1922
rect 4086 1918 4090 1922
rect 4358 1918 4362 1922
rect 4406 1918 4410 1922
rect 4494 1918 4498 1922
rect 4510 1918 4514 1922
rect 4566 1918 4570 1922
rect 4606 1918 4610 1922
rect 4654 1918 4658 1922
rect 4702 1918 4706 1922
rect 4710 1918 4714 1922
rect 4766 1918 4770 1922
rect 5206 1918 5210 1922
rect 5262 1918 5266 1922
rect 1086 1908 1090 1912
rect 1750 1908 1754 1912
rect 2478 1908 2482 1912
rect 4470 1908 4474 1912
rect 4758 1908 4762 1912
rect 858 1903 862 1907
rect 865 1903 869 1907
rect 1874 1903 1878 1907
rect 1881 1903 1885 1907
rect 2906 1903 2910 1907
rect 2913 1903 2917 1907
rect 3930 1903 3934 1907
rect 3937 1903 3941 1907
rect 4954 1903 4958 1907
rect 4961 1903 4965 1907
rect 990 1898 994 1902
rect 1134 1898 1138 1902
rect 1806 1898 1810 1902
rect 1990 1898 1994 1902
rect 2198 1898 2202 1902
rect 4246 1898 4250 1902
rect 4414 1898 4418 1902
rect 4526 1898 4530 1902
rect 4550 1898 4554 1902
rect 4614 1898 4618 1902
rect 4630 1898 4634 1902
rect 4638 1898 4642 1902
rect 4718 1898 4722 1902
rect 14 1888 18 1892
rect 22 1888 26 1892
rect 70 1888 74 1892
rect 158 1888 162 1892
rect 190 1888 194 1892
rect 398 1888 402 1892
rect 406 1888 410 1892
rect 454 1888 458 1892
rect 502 1888 506 1892
rect 534 1888 538 1892
rect 878 1888 882 1892
rect 966 1888 970 1892
rect 1014 1888 1018 1892
rect 1030 1888 1034 1892
rect 1102 1888 1106 1892
rect 1166 1888 1170 1892
rect 1190 1888 1194 1892
rect 1206 1888 1210 1892
rect 1318 1888 1322 1892
rect 1430 1888 1434 1892
rect 1558 1888 1562 1892
rect 1606 1888 1610 1892
rect 1646 1888 1650 1892
rect 1702 1888 1706 1892
rect 1718 1888 1722 1892
rect 1830 1888 1834 1892
rect 2182 1888 2186 1892
rect 2222 1888 2226 1892
rect 2238 1888 2242 1892
rect 2246 1888 2250 1892
rect 2278 1888 2282 1892
rect 2302 1888 2306 1892
rect 2430 1888 2434 1892
rect 2462 1888 2466 1892
rect 2694 1888 2698 1892
rect 2766 1888 2770 1892
rect 2814 1888 2818 1892
rect 2838 1888 2842 1892
rect 2958 1888 2962 1892
rect 2998 1888 3002 1892
rect 3110 1888 3114 1892
rect 3214 1888 3218 1892
rect 3486 1888 3490 1892
rect 3598 1888 3602 1892
rect 3606 1888 3610 1892
rect 3742 1888 3746 1892
rect 3838 1888 3842 1892
rect 3934 1888 3938 1892
rect 4070 1888 4074 1892
rect 4142 1888 4146 1892
rect 4166 1888 4170 1892
rect 4310 1888 4314 1892
rect 4686 1888 4690 1892
rect 4790 1888 4794 1892
rect 4798 1888 4802 1892
rect 4854 1888 4858 1892
rect 4926 1888 4930 1892
rect 4998 1888 5002 1892
rect 5054 1888 5058 1892
rect 5230 1888 5234 1892
rect 62 1878 66 1882
rect 110 1878 114 1882
rect 302 1878 306 1882
rect 334 1878 338 1882
rect 374 1878 378 1882
rect 382 1878 386 1882
rect 550 1878 554 1882
rect 566 1878 570 1882
rect 750 1878 754 1882
rect 838 1878 842 1882
rect 878 1878 882 1882
rect 990 1878 994 1882
rect 1054 1878 1058 1882
rect 1310 1878 1314 1882
rect 1582 1878 1586 1882
rect 1598 1878 1602 1882
rect 1614 1878 1618 1882
rect 1662 1879 1666 1883
rect 1710 1878 1714 1882
rect 6 1868 10 1872
rect 54 1868 58 1872
rect 78 1868 82 1872
rect 126 1868 130 1872
rect 166 1868 170 1872
rect 182 1868 186 1872
rect 238 1868 242 1872
rect 270 1868 274 1872
rect 286 1868 290 1872
rect 326 1868 330 1872
rect 390 1868 394 1872
rect 438 1868 442 1872
rect 446 1868 450 1872
rect 470 1868 474 1872
rect 518 1868 522 1872
rect 526 1868 530 1872
rect 654 1868 658 1872
rect 742 1868 746 1872
rect 782 1868 786 1872
rect 86 1858 90 1862
rect 110 1858 114 1862
rect 182 1858 186 1862
rect 214 1858 218 1862
rect 246 1858 250 1862
rect 254 1858 258 1862
rect 350 1858 354 1862
rect 550 1858 554 1862
rect 638 1859 642 1863
rect 790 1858 794 1862
rect 814 1858 818 1862
rect 942 1868 946 1872
rect 958 1868 962 1872
rect 982 1868 986 1872
rect 1038 1868 1042 1872
rect 1094 1868 1098 1872
rect 1142 1868 1146 1872
rect 1150 1868 1154 1872
rect 1198 1868 1202 1872
rect 1238 1868 1242 1872
rect 1254 1868 1258 1872
rect 1526 1868 1530 1872
rect 1574 1868 1578 1872
rect 1622 1868 1626 1872
rect 1678 1868 1682 1872
rect 1726 1868 1730 1872
rect 1742 1868 1746 1872
rect 1758 1868 1762 1872
rect 1766 1868 1770 1872
rect 1822 1868 1826 1872
rect 2094 1878 2098 1882
rect 2102 1878 2106 1882
rect 2166 1878 2170 1882
rect 2190 1878 2194 1882
rect 2198 1878 2202 1882
rect 2342 1878 2346 1882
rect 2470 1878 2474 1882
rect 2598 1878 2602 1882
rect 2686 1878 2690 1882
rect 2758 1878 2762 1882
rect 2798 1878 2802 1882
rect 2806 1878 2810 1882
rect 2910 1878 2914 1882
rect 2926 1878 2930 1882
rect 3166 1878 3170 1882
rect 3238 1878 3242 1882
rect 3254 1878 3258 1882
rect 3334 1878 3338 1882
rect 3350 1878 3354 1882
rect 3366 1878 3370 1882
rect 3982 1878 3986 1882
rect 4246 1878 4250 1882
rect 4254 1878 4258 1882
rect 4342 1878 4346 1882
rect 4414 1878 4418 1882
rect 4422 1878 4426 1882
rect 4526 1878 4530 1882
rect 4534 1878 4538 1882
rect 4614 1878 4618 1882
rect 4638 1878 4642 1882
rect 4718 1878 4722 1882
rect 5158 1878 5162 1882
rect 5214 1878 5218 1882
rect 5294 1878 5298 1882
rect 1934 1868 1938 1872
rect 1950 1868 1954 1872
rect 1998 1868 2002 1872
rect 918 1858 922 1862
rect 1014 1858 1018 1862
rect 1030 1858 1034 1862
rect 1078 1858 1082 1862
rect 1270 1859 1274 1863
rect 1302 1858 1306 1862
rect 1350 1858 1354 1862
rect 1382 1859 1386 1863
rect 1462 1858 1466 1862
rect 1494 1859 1498 1863
rect 1598 1858 1602 1862
rect 1630 1858 1634 1862
rect 1670 1858 1674 1862
rect 1686 1858 1690 1862
rect 1734 1858 1738 1862
rect 1926 1858 1930 1862
rect 1942 1858 1946 1862
rect 2014 1858 2018 1862
rect 2054 1858 2058 1862
rect 2070 1868 2074 1872
rect 2110 1868 2114 1872
rect 2150 1868 2154 1872
rect 2206 1868 2210 1872
rect 2246 1868 2250 1872
rect 2262 1866 2266 1870
rect 2286 1868 2290 1872
rect 2326 1868 2330 1872
rect 2374 1868 2378 1872
rect 2382 1868 2386 1872
rect 2414 1868 2418 1872
rect 2438 1868 2442 1872
rect 2590 1868 2594 1872
rect 2598 1868 2602 1872
rect 2630 1868 2634 1872
rect 2662 1868 2666 1872
rect 2710 1866 2714 1870
rect 2718 1868 2722 1872
rect 2734 1868 2738 1872
rect 2750 1868 2754 1872
rect 2774 1868 2778 1872
rect 2838 1868 2842 1872
rect 2854 1868 2858 1872
rect 2862 1868 2866 1872
rect 2918 1868 2922 1872
rect 2966 1868 2970 1872
rect 2094 1858 2098 1862
rect 2118 1858 2122 1862
rect 2142 1858 2146 1862
rect 2174 1858 2178 1862
rect 2246 1858 2250 1862
rect 3094 1868 3098 1872
rect 3118 1868 3122 1872
rect 3134 1868 3138 1872
rect 3174 1868 3178 1872
rect 3198 1868 3202 1872
rect 3302 1868 3306 1872
rect 3406 1868 3410 1872
rect 3430 1868 3434 1872
rect 3502 1868 3506 1872
rect 3686 1868 3690 1872
rect 3702 1868 3706 1872
rect 3718 1868 3722 1872
rect 3854 1868 3858 1872
rect 4054 1868 4058 1872
rect 4102 1868 4106 1872
rect 4110 1868 4114 1872
rect 4158 1868 4162 1872
rect 4166 1868 4170 1872
rect 4182 1868 4186 1872
rect 4238 1868 4242 1872
rect 4270 1868 4274 1872
rect 4278 1866 4282 1870
rect 4302 1868 4306 1872
rect 4350 1868 4354 1872
rect 4366 1868 4370 1872
rect 4390 1868 4394 1872
rect 4462 1868 4466 1872
rect 4518 1868 4522 1872
rect 4670 1868 4674 1872
rect 4686 1868 4690 1872
rect 4694 1868 4698 1872
rect 4710 1868 4714 1872
rect 4774 1868 4778 1872
rect 4782 1868 4786 1872
rect 2326 1858 2330 1862
rect 2342 1858 2346 1862
rect 2366 1858 2370 1862
rect 2446 1858 2450 1862
rect 2494 1858 2498 1862
rect 2526 1858 2530 1862
rect 2558 1858 2562 1862
rect 2622 1858 2626 1862
rect 2630 1858 2634 1862
rect 2654 1858 2658 1862
rect 2670 1858 2674 1862
rect 2742 1858 2746 1862
rect 2782 1858 2786 1862
rect 2830 1858 2834 1862
rect 2870 1858 2874 1862
rect 2886 1858 2890 1862
rect 2894 1858 2898 1862
rect 2942 1858 2946 1862
rect 2974 1858 2978 1862
rect 2990 1858 2994 1862
rect 3030 1858 3034 1862
rect 3046 1858 3050 1862
rect 3142 1858 3146 1862
rect 3158 1858 3162 1862
rect 3198 1858 3202 1862
rect 3286 1859 3290 1863
rect 3334 1858 3338 1862
rect 3350 1858 3354 1862
rect 3398 1858 3402 1862
rect 3550 1858 3554 1862
rect 3566 1858 3570 1862
rect 3670 1859 3674 1863
rect 3726 1858 3730 1862
rect 3774 1859 3778 1863
rect 3806 1858 3810 1862
rect 3870 1859 3874 1863
rect 3902 1858 3906 1862
rect 3982 1859 3986 1863
rect 4190 1858 4194 1862
rect 4198 1858 4202 1862
rect 4254 1858 4258 1862
rect 4310 1858 4314 1862
rect 4358 1858 4362 1862
rect 4398 1858 4402 1862
rect 4446 1858 4450 1862
rect 4478 1858 4482 1862
rect 4558 1858 4562 1862
rect 4590 1858 4594 1862
rect 4614 1858 4618 1862
rect 4630 1858 4634 1862
rect 4662 1858 4666 1862
rect 4838 1868 4842 1872
rect 4886 1868 4890 1872
rect 4894 1868 4898 1872
rect 4942 1868 4946 1872
rect 4950 1868 4954 1872
rect 5014 1868 5018 1872
rect 5022 1868 5026 1872
rect 5070 1868 5074 1872
rect 5078 1868 5082 1872
rect 5126 1868 5130 1872
rect 5166 1868 5170 1872
rect 4838 1858 4842 1862
rect 5134 1858 5138 1862
rect 5190 1858 5194 1862
rect 5238 1858 5242 1862
rect 5270 1858 5274 1862
rect 5278 1858 5282 1862
rect 118 1848 122 1852
rect 142 1848 146 1852
rect 198 1848 202 1852
rect 206 1848 210 1852
rect 262 1848 266 1852
rect 270 1848 274 1852
rect 286 1848 290 1852
rect 326 1848 330 1852
rect 462 1848 466 1852
rect 542 1848 546 1852
rect 726 1848 730 1852
rect 886 1848 890 1852
rect 910 1848 914 1852
rect 942 1848 946 1852
rect 966 1848 970 1852
rect 998 1848 1002 1852
rect 1014 1848 1018 1852
rect 1046 1848 1050 1852
rect 1054 1848 1058 1852
rect 1758 1848 1762 1852
rect 1838 1848 1842 1852
rect 2006 1848 2010 1852
rect 2038 1848 2042 1852
rect 2086 1848 2090 1852
rect 2134 1848 2138 1852
rect 2230 1848 2234 1852
rect 2302 1848 2306 1852
rect 2422 1848 2426 1852
rect 2438 1848 2442 1852
rect 2502 1848 2506 1852
rect 2534 1848 2538 1852
rect 2566 1848 2570 1852
rect 2606 1848 2610 1852
rect 2638 1848 2642 1852
rect 2726 1848 2730 1852
rect 2838 1848 2842 1852
rect 2958 1848 2962 1852
rect 2990 1848 2994 1852
rect 3110 1848 3114 1852
rect 3134 1848 3138 1852
rect 3158 1848 3162 1852
rect 3214 1848 3218 1852
rect 3342 1848 3346 1852
rect 3398 1848 3402 1852
rect 3446 1848 3450 1852
rect 3718 1848 3722 1852
rect 4182 1848 4186 1852
rect 4326 1848 4330 1852
rect 4470 1848 4474 1852
rect 4582 1848 4586 1852
rect 4670 1848 4674 1852
rect 5246 1848 5250 1852
rect 102 1838 106 1842
rect 214 1838 218 1842
rect 222 1838 226 1842
rect 806 1838 810 1842
rect 926 1838 930 1842
rect 2022 1838 2026 1842
rect 2518 1838 2522 1842
rect 2550 1838 2554 1842
rect 2670 1838 2674 1842
rect 3326 1838 3330 1842
rect 4046 1838 4050 1842
rect 4206 1838 4210 1842
rect 4222 1838 4226 1842
rect 4462 1838 4466 1842
rect 4486 1838 4490 1842
rect 4502 1838 4506 1842
rect 4566 1838 4570 1842
rect 4598 1838 4602 1842
rect 5182 1838 5186 1842
rect 5230 1838 5234 1842
rect 5262 1838 5266 1842
rect 574 1818 578 1822
rect 686 1818 690 1822
rect 766 1818 770 1822
rect 798 1818 802 1822
rect 846 1818 850 1822
rect 918 1818 922 1822
rect 1078 1818 1082 1822
rect 1790 1818 1794 1822
rect 1862 1818 1866 1822
rect 1966 1818 1970 1822
rect 2030 1818 2034 1822
rect 2054 1818 2058 1822
rect 2118 1818 2122 1822
rect 2166 1818 2170 1822
rect 2310 1818 2314 1822
rect 2326 1818 2330 1822
rect 2390 1818 2394 1822
rect 2478 1818 2482 1822
rect 2558 1818 2562 1822
rect 2742 1818 2746 1822
rect 4086 1818 4090 1822
rect 4214 1818 4218 1822
rect 4310 1818 4314 1822
rect 4422 1818 4426 1822
rect 4478 1818 4482 1822
rect 4542 1818 4546 1822
rect 4558 1818 4562 1822
rect 4590 1818 4594 1822
rect 4638 1818 4642 1822
rect 4742 1818 4746 1822
rect 5094 1818 5098 1822
rect 5214 1818 5218 1822
rect 5270 1818 5274 1822
rect 346 1803 350 1807
rect 353 1803 357 1807
rect 1370 1803 1374 1807
rect 1377 1803 1381 1807
rect 2394 1803 2398 1807
rect 2401 1803 2405 1807
rect 3418 1803 3422 1807
rect 3425 1803 3429 1807
rect 4442 1803 4446 1807
rect 4449 1803 4453 1807
rect 38 1788 42 1792
rect 78 1788 82 1792
rect 118 1788 122 1792
rect 158 1788 162 1792
rect 198 1788 202 1792
rect 326 1788 330 1792
rect 470 1788 474 1792
rect 518 1788 522 1792
rect 582 1788 586 1792
rect 670 1788 674 1792
rect 1006 1788 1010 1792
rect 1254 1788 1258 1792
rect 1318 1788 1322 1792
rect 1582 1788 1586 1792
rect 1606 1788 1610 1792
rect 1686 1788 1690 1792
rect 1710 1788 1714 1792
rect 1742 1788 1746 1792
rect 1806 1788 1810 1792
rect 1894 1788 1898 1792
rect 1934 1788 1938 1792
rect 1998 1788 2002 1792
rect 2014 1788 2018 1792
rect 2102 1788 2106 1792
rect 2134 1788 2138 1792
rect 2614 1788 2618 1792
rect 2638 1788 2642 1792
rect 2830 1788 2834 1792
rect 2870 1788 2874 1792
rect 2990 1788 2994 1792
rect 3022 1788 3026 1792
rect 3054 1788 3058 1792
rect 3270 1788 3274 1792
rect 3550 1788 3554 1792
rect 4062 1788 4066 1792
rect 4910 1788 4914 1792
rect 4358 1778 4362 1782
rect 6 1768 10 1772
rect 30 1768 34 1772
rect 78 1768 82 1772
rect 86 1768 90 1772
rect 142 1768 146 1772
rect 174 1768 178 1772
rect 286 1768 290 1772
rect 398 1768 402 1772
rect 422 1768 426 1772
rect 894 1768 898 1772
rect 902 1768 906 1772
rect 1014 1768 1018 1772
rect 1150 1768 1154 1772
rect 1430 1768 1434 1772
rect 1718 1768 1722 1772
rect 1990 1768 1994 1772
rect 2110 1768 2114 1772
rect 2270 1768 2274 1772
rect 2318 1768 2322 1772
rect 2558 1768 2562 1772
rect 2646 1768 2650 1772
rect 3014 1768 3018 1772
rect 3046 1768 3050 1772
rect 3614 1768 3618 1772
rect 4190 1768 4194 1772
rect 4270 1768 4274 1772
rect 4350 1768 4354 1772
rect 4366 1768 4370 1772
rect 4710 1768 4714 1772
rect 4742 1768 4746 1772
rect 4750 1768 4754 1772
rect 4854 1768 4858 1772
rect 4878 1768 4882 1772
rect 4886 1768 4890 1772
rect 4918 1768 4922 1772
rect 5014 1768 5018 1772
rect 70 1758 74 1762
rect 102 1758 106 1762
rect 262 1758 266 1762
rect 318 1758 322 1762
rect 382 1758 386 1762
rect 454 1758 458 1762
rect 462 1758 466 1762
rect 742 1758 746 1762
rect 38 1748 42 1752
rect 78 1748 82 1752
rect 118 1748 122 1752
rect 142 1748 146 1752
rect 254 1748 258 1752
rect 294 1748 298 1752
rect 366 1748 370 1752
rect 438 1748 442 1752
rect 446 1748 450 1752
rect 702 1748 706 1752
rect 734 1748 738 1752
rect 758 1748 762 1752
rect 886 1758 890 1762
rect 926 1758 930 1762
rect 974 1758 978 1762
rect 990 1758 994 1762
rect 998 1758 1002 1762
rect 1038 1758 1042 1762
rect 1094 1758 1098 1762
rect 822 1748 826 1752
rect 830 1748 834 1752
rect 894 1748 898 1752
rect 966 1748 970 1752
rect 974 1748 978 1752
rect 1006 1748 1010 1752
rect 1030 1748 1034 1752
rect 1086 1748 1090 1752
rect 1102 1748 1106 1752
rect 1678 1758 1682 1762
rect 1694 1758 1698 1762
rect 1702 1758 1706 1762
rect 1734 1758 1738 1762
rect 1782 1758 1786 1762
rect 1974 1758 1978 1762
rect 2006 1758 2010 1762
rect 2182 1758 2186 1762
rect 2286 1758 2290 1762
rect 1182 1748 1186 1752
rect 126 1738 130 1742
rect 150 1738 154 1742
rect 182 1738 186 1742
rect 238 1738 242 1742
rect 262 1738 266 1742
rect 278 1738 282 1742
rect 286 1738 290 1742
rect 334 1738 338 1742
rect 342 1738 346 1742
rect 374 1738 378 1742
rect 430 1738 434 1742
rect 502 1738 506 1742
rect 550 1738 554 1742
rect 558 1738 562 1742
rect 606 1738 610 1742
rect 614 1738 618 1742
rect 726 1738 730 1742
rect 750 1738 754 1742
rect 766 1738 770 1742
rect 774 1738 778 1742
rect 798 1738 802 1742
rect 822 1738 826 1742
rect 934 1738 938 1742
rect 950 1738 954 1742
rect 958 1738 962 1742
rect 1030 1738 1034 1742
rect 1070 1738 1074 1742
rect 1214 1747 1218 1751
rect 1350 1748 1354 1752
rect 1382 1747 1386 1751
rect 1462 1748 1466 1752
rect 1494 1747 1498 1751
rect 1542 1748 1546 1752
rect 1710 1748 1714 1752
rect 1870 1748 1874 1752
rect 1950 1748 1954 1752
rect 1982 1748 1986 1752
rect 2118 1748 2122 1752
rect 2150 1748 2154 1752
rect 2278 1748 2282 1752
rect 2318 1748 2322 1752
rect 2374 1758 2378 1762
rect 2462 1758 2466 1762
rect 2550 1758 2554 1762
rect 2574 1758 2578 1762
rect 2582 1758 2586 1762
rect 2630 1758 2634 1762
rect 2718 1758 2722 1762
rect 2862 1758 2866 1762
rect 2942 1758 2946 1762
rect 2998 1758 3002 1762
rect 3030 1758 3034 1762
rect 3190 1758 3194 1762
rect 3606 1758 3610 1762
rect 3742 1758 3746 1762
rect 3774 1758 3778 1762
rect 4198 1758 4202 1762
rect 4238 1758 4242 1762
rect 4278 1758 4282 1762
rect 4294 1758 4298 1762
rect 4342 1758 4346 1762
rect 4350 1758 4354 1762
rect 4382 1758 4386 1762
rect 4414 1758 4418 1762
rect 4430 1758 4434 1762
rect 4582 1758 4586 1762
rect 4598 1758 4602 1762
rect 4622 1758 4626 1762
rect 4638 1758 4642 1762
rect 4678 1758 4682 1762
rect 4702 1758 4706 1762
rect 4726 1758 4730 1762
rect 4734 1758 4738 1762
rect 4766 1758 4770 1762
rect 4806 1758 4810 1762
rect 4822 1758 4826 1762
rect 4902 1758 4906 1762
rect 5222 1758 5226 1762
rect 5302 1758 5306 1762
rect 2350 1748 2354 1752
rect 2454 1748 2458 1752
rect 2542 1748 2546 1752
rect 2566 1748 2570 1752
rect 2582 1748 2586 1752
rect 2614 1748 2618 1752
rect 2678 1748 2682 1752
rect 2726 1748 2730 1752
rect 2750 1748 2754 1752
rect 2766 1748 2770 1752
rect 2918 1748 2922 1752
rect 2974 1748 2978 1752
rect 3006 1748 3010 1752
rect 3038 1748 3042 1752
rect 1094 1738 1098 1742
rect 1142 1738 1146 1742
rect 1310 1738 1314 1742
rect 1422 1738 1426 1742
rect 1598 1738 1602 1742
rect 1670 1738 1674 1742
rect 1838 1738 1842 1742
rect 1926 1738 1930 1742
rect 1942 1738 1946 1742
rect 2046 1738 2050 1742
rect 2094 1738 2098 1742
rect 2158 1738 2162 1742
rect 2198 1738 2202 1742
rect 2206 1738 2210 1742
rect 2254 1738 2258 1742
rect 2294 1738 2298 1742
rect 2302 1738 2306 1742
rect 2310 1738 2314 1742
rect 2342 1738 2346 1742
rect 2358 1738 2362 1742
rect 2422 1738 2426 1742
rect 2446 1738 2450 1742
rect 2478 1738 2482 1742
rect 2502 1738 2506 1742
rect 2534 1738 2538 1742
rect 3238 1747 3242 1751
rect 3302 1748 3306 1752
rect 3334 1747 3338 1751
rect 3390 1747 3394 1751
rect 3494 1748 3498 1752
rect 3518 1748 3522 1752
rect 3534 1748 3538 1752
rect 3558 1748 3562 1752
rect 3566 1748 3570 1752
rect 2598 1738 2602 1742
rect 2606 1738 2610 1742
rect 2710 1738 2714 1742
rect 2742 1738 2746 1742
rect 2774 1738 2778 1742
rect 2822 1738 2826 1742
rect 2846 1738 2850 1742
rect 2862 1738 2866 1742
rect 2878 1738 2882 1742
rect 2926 1738 2930 1742
rect 2934 1738 2938 1742
rect 2942 1738 2946 1742
rect 3062 1738 3066 1742
rect 3110 1738 3114 1742
rect 3118 1738 3122 1742
rect 3166 1738 3170 1742
rect 3254 1738 3258 1742
rect 3406 1738 3410 1742
rect 3462 1738 3466 1742
rect 3502 1738 3506 1742
rect 3678 1747 3682 1751
rect 3710 1748 3714 1752
rect 3758 1748 3762 1752
rect 3894 1747 3898 1751
rect 3982 1748 3986 1752
rect 4206 1748 4210 1752
rect 4278 1748 4282 1752
rect 4334 1748 4338 1752
rect 4358 1748 4362 1752
rect 4414 1748 4418 1752
rect 4430 1748 4434 1752
rect 4486 1748 4490 1752
rect 4510 1748 4514 1752
rect 4542 1748 4546 1752
rect 4614 1748 4618 1752
rect 4662 1748 4666 1752
rect 4718 1748 4722 1752
rect 4742 1748 4746 1752
rect 4766 1748 4770 1752
rect 4806 1748 4810 1752
rect 4830 1748 4834 1752
rect 4846 1748 4850 1752
rect 4878 1748 4882 1752
rect 4910 1748 4914 1752
rect 4934 1748 4938 1752
rect 4974 1748 4978 1752
rect 5046 1748 5050 1752
rect 5070 1748 5074 1752
rect 5238 1748 5242 1752
rect 5270 1748 5274 1752
rect 3590 1738 3594 1742
rect 3694 1738 3698 1742
rect 3718 1738 3722 1742
rect 3766 1738 3770 1742
rect 3782 1738 3786 1742
rect 3790 1738 3794 1742
rect 3814 1738 3818 1742
rect 3862 1738 3866 1742
rect 3902 1738 3906 1742
rect 3910 1738 3914 1742
rect 3974 1738 3978 1742
rect 4046 1738 4050 1742
rect 4070 1738 4074 1742
rect 4118 1738 4122 1742
rect 4126 1738 4130 1742
rect 4182 1738 4186 1742
rect 4214 1738 4218 1742
rect 4254 1738 4258 1742
rect 4406 1738 4410 1742
rect 4438 1738 4442 1742
rect 4550 1738 4554 1742
rect 4566 1738 4570 1742
rect 4606 1738 4610 1742
rect 4678 1738 4682 1742
rect 4694 1738 4698 1742
rect 4798 1738 4802 1742
rect 4942 1738 4946 1742
rect 5006 1738 5010 1742
rect 5110 1738 5114 1742
rect 5166 1738 5170 1742
rect 5246 1738 5250 1742
rect 5262 1738 5266 1742
rect 14 1728 18 1732
rect 62 1728 66 1732
rect 142 1728 146 1732
rect 238 1728 242 1732
rect 398 1728 402 1732
rect 406 1728 410 1732
rect 494 1728 498 1732
rect 686 1728 690 1732
rect 702 1728 706 1732
rect 918 1728 922 1732
rect 1118 1728 1122 1732
rect 1614 1728 1618 1732
rect 1766 1728 1770 1732
rect 1782 1728 1786 1732
rect 1846 1728 1850 1732
rect 2038 1728 2042 1732
rect 2142 1728 2146 1732
rect 2174 1728 2178 1732
rect 2374 1728 2378 1732
rect 2422 1728 2426 1732
rect 2430 1728 2434 1732
rect 2486 1728 2490 1732
rect 2510 1728 2514 1732
rect 2518 1728 2522 1732
rect 2526 1728 2530 1732
rect 2646 1728 2650 1732
rect 2654 1728 2658 1732
rect 2710 1728 2714 1732
rect 2750 1728 2754 1732
rect 2854 1728 2858 1732
rect 2950 1728 2954 1732
rect 2982 1728 2986 1732
rect 3478 1728 3482 1732
rect 3518 1728 3522 1732
rect 3542 1728 3546 1732
rect 3798 1728 3802 1732
rect 3830 1728 3834 1732
rect 3862 1728 3866 1732
rect 4054 1728 4058 1732
rect 4230 1728 4234 1732
rect 4382 1728 4386 1732
rect 4462 1728 4466 1732
rect 4494 1728 4498 1732
rect 4510 1728 4514 1732
rect 4550 1728 4554 1732
rect 4830 1728 4834 1732
rect 4854 1728 4858 1732
rect 4958 1728 4962 1732
rect 5006 1728 5010 1732
rect 5278 1728 5282 1732
rect 262 1718 266 1722
rect 310 1718 314 1722
rect 342 1718 346 1722
rect 694 1718 698 1722
rect 718 1718 722 1722
rect 822 1718 826 1722
rect 958 1718 962 1722
rect 1126 1718 1130 1722
rect 1254 1718 1258 1722
rect 1934 1718 1938 1722
rect 2078 1718 2082 1722
rect 2166 1718 2170 1722
rect 2182 1718 2186 1722
rect 2222 1718 2226 1722
rect 2278 1718 2282 1722
rect 2414 1718 2418 1722
rect 2462 1718 2466 1722
rect 2758 1718 2762 1722
rect 2790 1718 2794 1722
rect 2918 1718 2922 1722
rect 3078 1718 3082 1722
rect 3134 1718 3138 1722
rect 3454 1718 3458 1722
rect 3526 1718 3530 1722
rect 3598 1718 3602 1722
rect 3726 1718 3730 1722
rect 3806 1718 3810 1722
rect 4086 1718 4090 1722
rect 4142 1718 4146 1722
rect 4222 1718 4226 1722
rect 4270 1718 4274 1722
rect 4294 1718 4298 1722
rect 4470 1718 4474 1722
rect 4526 1718 4530 1722
rect 4558 1718 4562 1722
rect 4646 1718 4650 1722
rect 4678 1718 4682 1722
rect 4950 1718 4954 1722
rect 5134 1718 5138 1722
rect 238 1708 242 1712
rect 422 1708 426 1712
rect 1118 1708 1122 1712
rect 2878 1708 2882 1712
rect 858 1703 862 1707
rect 865 1703 869 1707
rect 1874 1703 1878 1707
rect 1881 1703 1885 1707
rect 2906 1703 2910 1707
rect 2913 1703 2917 1707
rect 3930 1703 3934 1707
rect 3937 1703 3941 1707
rect 4954 1703 4958 1707
rect 4961 1703 4965 1707
rect 374 1698 378 1702
rect 1030 1698 1034 1702
rect 86 1688 90 1692
rect 142 1688 146 1692
rect 198 1688 202 1692
rect 206 1688 210 1692
rect 222 1688 226 1692
rect 438 1688 442 1692
rect 542 1688 546 1692
rect 598 1688 602 1692
rect 670 1688 674 1692
rect 934 1688 938 1692
rect 998 1688 1002 1692
rect 1022 1688 1026 1692
rect 1222 1688 1226 1692
rect 1358 1688 1362 1692
rect 1502 1688 1506 1692
rect 1614 1688 1618 1692
rect 1758 1688 1762 1692
rect 1806 1688 1810 1692
rect 1838 1688 1842 1692
rect 1902 1688 1906 1692
rect 1958 1688 1962 1692
rect 1982 1688 1986 1692
rect 2006 1688 2010 1692
rect 2046 1688 2050 1692
rect 2102 1688 2106 1692
rect 2390 1688 2394 1692
rect 2446 1688 2450 1692
rect 2534 1688 2538 1692
rect 2558 1688 2562 1692
rect 2574 1688 2578 1692
rect 2606 1688 2610 1692
rect 2694 1688 2698 1692
rect 2806 1688 2810 1692
rect 2846 1688 2850 1692
rect 2974 1688 2978 1692
rect 2982 1688 2986 1692
rect 3078 1688 3082 1692
rect 3286 1688 3290 1692
rect 3342 1688 3346 1692
rect 3510 1688 3514 1692
rect 3654 1688 3658 1692
rect 3694 1688 3698 1692
rect 3710 1688 3714 1692
rect 4006 1688 4010 1692
rect 4014 1688 4018 1692
rect 4254 1688 4258 1692
rect 4462 1688 4466 1692
rect 4814 1688 4818 1692
rect 4878 1688 4882 1692
rect 4990 1688 4994 1692
rect 5038 1688 5042 1692
rect 5150 1688 5154 1692
rect 5190 1688 5194 1692
rect 5278 1688 5282 1692
rect 5286 1688 5290 1692
rect 366 1678 370 1682
rect 374 1678 378 1682
rect 694 1678 698 1682
rect 702 1678 706 1682
rect 782 1678 786 1682
rect 814 1678 818 1682
rect 822 1678 826 1682
rect 838 1678 842 1682
rect 870 1678 874 1682
rect 926 1678 930 1682
rect 1046 1678 1050 1682
rect 1134 1678 1138 1682
rect 1182 1678 1186 1682
rect 1326 1678 1330 1682
rect 1654 1678 1658 1682
rect 1814 1678 1818 1682
rect 1894 1678 1898 1682
rect 1966 1678 1970 1682
rect 1974 1678 1978 1682
rect 2214 1678 2218 1682
rect 2254 1678 2258 1682
rect 2262 1678 2266 1682
rect 2294 1678 2298 1682
rect 2374 1678 2378 1682
rect 2406 1678 2410 1682
rect 2502 1678 2506 1682
rect 2550 1678 2554 1682
rect 2598 1678 2602 1682
rect 3254 1678 3258 1682
rect 3334 1678 3338 1682
rect 3374 1678 3378 1682
rect 3446 1678 3450 1682
rect 54 1668 58 1672
rect 102 1668 106 1672
rect 110 1668 114 1672
rect 158 1668 162 1672
rect 166 1668 170 1672
rect 214 1668 218 1672
rect 246 1668 250 1672
rect 302 1668 306 1672
rect 310 1668 314 1672
rect 318 1666 322 1670
rect 350 1668 354 1672
rect 422 1668 426 1672
rect 430 1668 434 1672
rect 478 1668 482 1672
rect 486 1668 490 1672
rect 534 1668 538 1672
rect 558 1668 562 1672
rect 566 1668 570 1672
rect 614 1668 618 1672
rect 622 1668 626 1672
rect 654 1668 658 1672
rect 670 1668 674 1672
rect 702 1668 706 1672
rect 750 1668 754 1672
rect 782 1668 786 1672
rect 798 1668 802 1672
rect 846 1668 850 1672
rect 886 1668 890 1672
rect 902 1668 906 1672
rect 918 1668 922 1672
rect 942 1668 946 1672
rect 990 1668 994 1672
rect 1038 1668 1042 1672
rect 1166 1668 1170 1672
rect 1214 1668 1218 1672
rect 1254 1668 1258 1672
rect 1326 1668 1330 1672
rect 1398 1668 1402 1672
rect 1462 1668 1466 1672
rect 1486 1668 1490 1672
rect 1598 1668 1602 1672
rect 1646 1668 1650 1672
rect 1670 1668 1674 1672
rect 22 1658 26 1662
rect 46 1658 50 1662
rect 238 1658 242 1662
rect 262 1658 266 1662
rect 374 1658 378 1662
rect 390 1658 394 1662
rect 414 1658 418 1662
rect 630 1658 634 1662
rect 678 1658 682 1662
rect 718 1658 722 1662
rect 742 1658 746 1662
rect 758 1658 762 1662
rect 774 1658 778 1662
rect 806 1658 810 1662
rect 894 1658 898 1662
rect 950 1658 954 1662
rect 974 1658 978 1662
rect 1046 1658 1050 1662
rect 1078 1658 1082 1662
rect 1102 1658 1106 1662
rect 1142 1658 1146 1662
rect 1158 1658 1162 1662
rect 1166 1658 1170 1662
rect 1206 1658 1210 1662
rect 1286 1659 1290 1663
rect 1470 1659 1474 1663
rect 1534 1658 1538 1662
rect 1566 1659 1570 1663
rect 1670 1658 1674 1662
rect 1686 1658 1690 1662
rect 1742 1668 1746 1672
rect 1790 1668 1794 1672
rect 1822 1668 1826 1672
rect 1894 1668 1898 1672
rect 1910 1668 1914 1672
rect 1942 1668 1946 1672
rect 1990 1668 1994 1672
rect 2022 1668 2026 1672
rect 2030 1668 2034 1672
rect 2086 1668 2090 1672
rect 2134 1668 2138 1672
rect 2158 1668 2162 1672
rect 2166 1668 2170 1672
rect 2214 1668 2218 1672
rect 2278 1668 2282 1672
rect 2342 1668 2346 1672
rect 2366 1668 2370 1672
rect 2398 1668 2402 1672
rect 2406 1668 2410 1672
rect 2470 1668 2474 1672
rect 2510 1668 2514 1672
rect 2526 1668 2530 1672
rect 2590 1668 2594 1672
rect 2614 1668 2618 1672
rect 2678 1668 2682 1672
rect 2814 1668 2818 1672
rect 2878 1668 2882 1672
rect 3102 1668 3106 1672
rect 3134 1668 3138 1672
rect 3182 1668 3186 1672
rect 3310 1668 3314 1672
rect 3318 1668 3322 1672
rect 3366 1668 3370 1672
rect 3430 1668 3434 1672
rect 3526 1678 3530 1682
rect 3590 1678 3594 1682
rect 3606 1678 3610 1682
rect 3614 1678 3618 1682
rect 4342 1678 4346 1682
rect 4382 1678 4386 1682
rect 4590 1678 4594 1682
rect 4750 1678 4754 1682
rect 4758 1678 4762 1682
rect 5110 1678 5114 1682
rect 5142 1678 5146 1682
rect 5174 1678 5178 1682
rect 5182 1678 5186 1682
rect 5214 1678 5218 1682
rect 3518 1668 3522 1672
rect 3558 1668 3562 1672
rect 3630 1668 3634 1672
rect 3662 1668 3666 1672
rect 3702 1668 3706 1672
rect 3790 1668 3794 1672
rect 3830 1668 3834 1672
rect 3846 1668 3850 1672
rect 3958 1668 3962 1672
rect 4110 1668 4114 1672
rect 4158 1668 4162 1672
rect 4166 1668 4170 1672
rect 4214 1668 4218 1672
rect 1718 1658 1722 1662
rect 1734 1658 1738 1662
rect 1798 1658 1802 1662
rect 1918 1658 1922 1662
rect 1934 1658 1938 1662
rect 1998 1658 2002 1662
rect 2174 1658 2178 1662
rect 2230 1658 2234 1662
rect 2246 1658 2250 1662
rect 2270 1658 2274 1662
rect 2342 1658 2346 1662
rect 2454 1658 2458 1662
rect 2470 1658 2474 1662
rect 2622 1658 2626 1662
rect 2694 1658 2698 1662
rect 2742 1659 2746 1663
rect 2774 1658 2778 1662
rect 2910 1659 2914 1663
rect 2942 1658 2946 1662
rect 3022 1658 3026 1662
rect 3046 1659 3050 1663
rect 3094 1658 3098 1662
rect 3134 1658 3138 1662
rect 3254 1659 3258 1663
rect 3302 1658 3306 1662
rect 3318 1658 3322 1662
rect 3358 1658 3362 1662
rect 3422 1658 3426 1662
rect 3454 1658 3458 1662
rect 3470 1658 3474 1662
rect 3494 1658 3498 1662
rect 3542 1658 3546 1662
rect 3566 1658 3570 1662
rect 3582 1658 3586 1662
rect 3590 1658 3594 1662
rect 3638 1658 3642 1662
rect 3774 1659 3778 1663
rect 3838 1658 3842 1662
rect 3950 1658 3954 1662
rect 4046 1658 4050 1662
rect 4078 1659 4082 1663
rect 4230 1658 4234 1662
rect 4270 1658 4274 1662
rect 4286 1668 4290 1672
rect 4342 1668 4346 1672
rect 4398 1668 4402 1672
rect 4406 1668 4410 1672
rect 4422 1668 4426 1672
rect 4446 1668 4450 1672
rect 4494 1668 4498 1672
rect 4502 1668 4506 1672
rect 4518 1668 4522 1672
rect 4582 1668 4586 1672
rect 4590 1668 4594 1672
rect 4606 1668 4610 1672
rect 4710 1668 4714 1672
rect 4758 1668 4762 1672
rect 4806 1668 4810 1672
rect 4318 1658 4322 1662
rect 4342 1658 4346 1662
rect 4358 1658 4362 1662
rect 4534 1658 4538 1662
rect 4574 1658 4578 1662
rect 4614 1658 4618 1662
rect 4662 1658 4666 1662
rect 4678 1658 4682 1662
rect 4718 1658 4722 1662
rect 4830 1666 4834 1670
rect 4838 1668 4842 1672
rect 4870 1668 4874 1672
rect 4902 1668 4906 1672
rect 4950 1668 4954 1672
rect 4990 1668 4994 1672
rect 5070 1668 5074 1672
rect 5102 1668 5106 1672
rect 5166 1668 5170 1672
rect 5198 1668 5202 1672
rect 5214 1668 5218 1672
rect 5230 1668 5234 1672
rect 5238 1668 5242 1672
rect 5294 1668 5298 1672
rect 4774 1658 4778 1662
rect 4782 1658 4786 1662
rect 4798 1658 4802 1662
rect 4846 1658 4850 1662
rect 4918 1659 4922 1663
rect 5094 1658 5098 1662
rect 5206 1658 5210 1662
rect 5246 1658 5250 1662
rect 254 1648 258 1652
rect 286 1648 290 1652
rect 398 1648 402 1652
rect 542 1648 546 1652
rect 630 1648 634 1652
rect 646 1648 650 1652
rect 670 1648 674 1652
rect 774 1648 778 1652
rect 830 1648 834 1652
rect 854 1648 858 1652
rect 902 1648 906 1652
rect 966 1648 970 1652
rect 1062 1648 1066 1652
rect 1086 1648 1090 1652
rect 1094 1648 1098 1652
rect 1326 1648 1330 1652
rect 1734 1648 1738 1652
rect 1886 1648 1890 1652
rect 2006 1648 2010 1652
rect 2142 1648 2146 1652
rect 2190 1648 2194 1652
rect 2302 1648 2306 1652
rect 2326 1648 2330 1652
rect 2382 1648 2386 1652
rect 2454 1648 2458 1652
rect 2526 1648 2530 1652
rect 2574 1648 2578 1652
rect 3366 1648 3370 1652
rect 3502 1648 3506 1652
rect 3526 1648 3530 1652
rect 3582 1648 3586 1652
rect 3630 1648 3634 1652
rect 3678 1648 3682 1652
rect 4222 1648 4226 1652
rect 4254 1648 4258 1652
rect 4302 1648 4306 1652
rect 4334 1648 4338 1652
rect 4502 1648 4506 1652
rect 4518 1648 4522 1652
rect 4526 1648 4530 1652
rect 4558 1648 4562 1652
rect 4622 1648 4626 1652
rect 4638 1648 4642 1652
rect 4670 1648 4674 1652
rect 4678 1648 4682 1652
rect 4886 1648 4890 1652
rect 5078 1648 5082 1652
rect 270 1638 274 1642
rect 302 1638 306 1642
rect 974 1638 978 1642
rect 1070 1638 1074 1642
rect 1102 1638 1106 1642
rect 1110 1638 1114 1642
rect 1182 1638 1186 1642
rect 1678 1638 1682 1642
rect 2646 1638 2650 1642
rect 2702 1638 2706 1642
rect 3190 1638 3194 1642
rect 3486 1638 3490 1642
rect 4238 1638 4242 1642
rect 4358 1638 4362 1642
rect 4654 1638 4658 1642
rect 262 1628 266 1632
rect 502 1628 506 1632
rect 1126 1628 1130 1632
rect 3494 1628 3498 1632
rect 3894 1628 3898 1632
rect 334 1618 338 1622
rect 414 1618 418 1622
rect 814 1618 818 1622
rect 966 1618 970 1622
rect 1206 1618 1210 1622
rect 1406 1618 1410 1622
rect 1718 1618 1722 1622
rect 2206 1618 2210 1622
rect 2294 1618 2298 1622
rect 2534 1618 2538 1622
rect 3150 1618 3154 1622
rect 3598 1618 3602 1622
rect 4126 1618 4130 1622
rect 4198 1618 4202 1622
rect 4246 1618 4250 1622
rect 4382 1618 4386 1622
rect 4534 1618 4538 1622
rect 4574 1618 4578 1622
rect 4630 1618 4634 1622
rect 4718 1618 4722 1622
rect 4742 1618 4746 1622
rect 5014 1618 5018 1622
rect 5094 1618 5098 1622
rect 5126 1618 5130 1622
rect 5214 1618 5218 1622
rect 346 1603 350 1607
rect 353 1603 357 1607
rect 1370 1603 1374 1607
rect 1377 1603 1381 1607
rect 2394 1603 2398 1607
rect 2401 1603 2405 1607
rect 3418 1603 3422 1607
rect 3425 1603 3429 1607
rect 4442 1603 4446 1607
rect 4449 1603 4453 1607
rect 326 1588 330 1592
rect 446 1588 450 1592
rect 574 1588 578 1592
rect 630 1588 634 1592
rect 950 1588 954 1592
rect 998 1588 1002 1592
rect 1270 1588 1274 1592
rect 1486 1588 1490 1592
rect 1702 1588 1706 1592
rect 1782 1588 1786 1592
rect 1814 1588 1818 1592
rect 1854 1588 1858 1592
rect 1878 1588 1882 1592
rect 1974 1588 1978 1592
rect 2014 1588 2018 1592
rect 2126 1588 2130 1592
rect 2166 1588 2170 1592
rect 2222 1588 2226 1592
rect 2254 1588 2258 1592
rect 2310 1588 2314 1592
rect 2510 1588 2514 1592
rect 2622 1588 2626 1592
rect 2790 1588 2794 1592
rect 3254 1588 3258 1592
rect 3382 1588 3386 1592
rect 3566 1588 3570 1592
rect 4150 1588 4154 1592
rect 4654 1588 4658 1592
rect 4694 1588 4698 1592
rect 4790 1588 4794 1592
rect 4942 1588 4946 1592
rect 5230 1588 5234 1592
rect 110 1578 114 1582
rect 678 1578 682 1582
rect 814 1578 818 1582
rect 4758 1578 4762 1582
rect 126 1568 130 1572
rect 230 1568 234 1572
rect 822 1568 826 1572
rect 878 1568 882 1572
rect 958 1568 962 1572
rect 982 1568 986 1572
rect 1006 1568 1010 1572
rect 1062 1568 1066 1572
rect 1518 1568 1522 1572
rect 1534 1568 1538 1572
rect 2302 1568 2306 1572
rect 2350 1568 2354 1572
rect 2542 1568 2546 1572
rect 2734 1568 2738 1572
rect 2998 1568 3002 1572
rect 3342 1568 3346 1572
rect 3406 1568 3410 1572
rect 4702 1568 4706 1572
rect 4766 1568 4770 1572
rect 4798 1568 4802 1572
rect 4894 1568 4898 1572
rect 4974 1568 4978 1572
rect 5174 1568 5178 1572
rect 5222 1568 5226 1572
rect 62 1558 66 1562
rect 78 1558 82 1562
rect 182 1558 186 1562
rect 206 1558 210 1562
rect 214 1558 218 1562
rect 310 1558 314 1562
rect 366 1558 370 1562
rect 382 1558 386 1562
rect 38 1548 42 1552
rect 54 1548 58 1552
rect 86 1548 90 1552
rect 126 1548 130 1552
rect 182 1548 186 1552
rect 222 1548 226 1552
rect 302 1548 306 1552
rect 326 1548 330 1552
rect 342 1548 346 1552
rect 382 1548 386 1552
rect 422 1548 426 1552
rect 598 1548 602 1552
rect 654 1558 658 1562
rect 670 1558 674 1562
rect 806 1558 810 1562
rect 846 1558 850 1562
rect 894 1558 898 1562
rect 942 1558 946 1562
rect 990 1558 994 1562
rect 1022 1558 1026 1562
rect 1046 1558 1050 1562
rect 1142 1558 1146 1562
rect 1686 1558 1690 1562
rect 1774 1558 1778 1562
rect 1798 1558 1802 1562
rect 2110 1558 2114 1562
rect 2286 1558 2290 1562
rect 2318 1558 2322 1562
rect 2366 1558 2370 1562
rect 2414 1558 2418 1562
rect 3294 1558 3298 1562
rect 3326 1558 3330 1562
rect 3422 1558 3426 1562
rect 3462 1558 3466 1562
rect 3662 1558 3666 1562
rect 4566 1558 4570 1562
rect 4598 1558 4602 1562
rect 4718 1558 4722 1562
rect 4742 1558 4746 1562
rect 4750 1558 4754 1562
rect 4782 1558 4786 1562
rect 4814 1558 4818 1562
rect 5062 1558 5066 1562
rect 5070 1558 5074 1562
rect 5126 1558 5130 1562
rect 5238 1558 5242 1562
rect 654 1548 658 1552
rect 710 1548 714 1552
rect 726 1548 730 1552
rect 734 1548 738 1552
rect 750 1548 754 1552
rect 814 1548 818 1552
rect 862 1548 866 1552
rect 886 1548 890 1552
rect 902 1548 906 1552
rect 934 1548 938 1552
rect 950 1548 954 1552
rect 982 1548 986 1552
rect 998 1548 1002 1552
rect 1022 1548 1026 1552
rect 1086 1548 1090 1552
rect 1118 1548 1122 1552
rect 1158 1548 1162 1552
rect 1230 1548 1234 1552
rect 1326 1548 1330 1552
rect 6 1538 10 1542
rect 22 1538 26 1542
rect 62 1538 66 1542
rect 118 1538 122 1542
rect 190 1538 194 1542
rect 286 1538 290 1542
rect 342 1538 346 1542
rect 358 1538 362 1542
rect 390 1538 394 1542
rect 430 1538 434 1542
rect 478 1538 482 1542
rect 486 1538 490 1542
rect 534 1538 538 1542
rect 542 1538 546 1542
rect 590 1538 594 1542
rect 638 1538 642 1542
rect 646 1538 650 1542
rect 718 1538 722 1542
rect 790 1538 794 1542
rect 910 1538 914 1542
rect 918 1538 922 1542
rect 926 1538 930 1542
rect 1038 1538 1042 1542
rect 1070 1538 1074 1542
rect 1078 1538 1082 1542
rect 1446 1547 1450 1551
rect 1494 1548 1498 1552
rect 1510 1548 1514 1552
rect 1582 1547 1586 1551
rect 1622 1548 1626 1552
rect 1646 1548 1650 1552
rect 1702 1548 1706 1552
rect 1734 1548 1738 1552
rect 1750 1548 1754 1552
rect 1814 1548 1818 1552
rect 1830 1548 1834 1552
rect 1878 1548 1882 1552
rect 1926 1548 1930 1552
rect 1934 1548 1938 1552
rect 1950 1548 1954 1552
rect 1966 1548 1970 1552
rect 1990 1548 1994 1552
rect 2038 1548 2042 1552
rect 2046 1548 2050 1552
rect 2102 1548 2106 1552
rect 2158 1548 2162 1552
rect 2230 1548 2234 1552
rect 2294 1548 2298 1552
rect 2358 1548 2362 1552
rect 2374 1548 2378 1552
rect 2446 1548 2450 1552
rect 2582 1548 2586 1552
rect 2678 1548 2682 1552
rect 2918 1548 2922 1552
rect 3030 1548 3034 1552
rect 3078 1548 3082 1552
rect 3086 1548 3090 1552
rect 3134 1548 3138 1552
rect 1110 1538 1114 1542
rect 1142 1538 1146 1542
rect 1166 1538 1170 1542
rect 1206 1538 1210 1542
rect 1254 1538 1258 1542
rect 1318 1538 1322 1542
rect 1462 1538 1466 1542
rect 1630 1538 1634 1542
rect 1678 1538 1682 1542
rect 1742 1538 1746 1542
rect 1790 1538 1794 1542
rect 1822 1538 1826 1542
rect 1838 1538 1842 1542
rect 1886 1538 1890 1542
rect 1894 1538 1898 1542
rect 1966 1538 1970 1542
rect 3190 1547 3194 1551
rect 3222 1548 3226 1552
rect 3262 1548 3266 1552
rect 3310 1548 3314 1552
rect 3414 1548 3418 1552
rect 3526 1548 3530 1552
rect 2054 1538 2058 1542
rect 2070 1538 2074 1542
rect 2102 1538 2106 1542
rect 2134 1538 2138 1542
rect 2182 1538 2186 1542
rect 2198 1538 2202 1542
rect 2270 1538 2274 1542
rect 2406 1538 2410 1542
rect 2454 1538 2458 1542
rect 2502 1538 2506 1542
rect 2606 1538 2610 1542
rect 2702 1538 2706 1542
rect 2718 1538 2722 1542
rect 2766 1538 2770 1542
rect 2774 1538 2778 1542
rect 2822 1538 2826 1542
rect 2830 1538 2834 1542
rect 2878 1538 2882 1542
rect 2926 1538 2930 1542
rect 2974 1538 2978 1542
rect 2982 1538 2986 1542
rect 3030 1538 3034 1542
rect 3150 1540 3154 1544
rect 3158 1538 3162 1542
rect 3270 1538 3274 1542
rect 3318 1538 3322 1542
rect 3342 1538 3346 1542
rect 3350 1538 3354 1542
rect 3366 1538 3370 1542
rect 3630 1547 3634 1551
rect 3686 1548 3690 1552
rect 3710 1548 3714 1552
rect 3726 1548 3730 1552
rect 3758 1547 3762 1551
rect 3790 1548 3794 1552
rect 3910 1548 3914 1552
rect 4014 1548 4018 1552
rect 4214 1547 4218 1551
rect 4414 1548 4418 1552
rect 4478 1548 4482 1552
rect 4486 1548 4490 1552
rect 4502 1548 4506 1552
rect 4534 1548 4538 1552
rect 4582 1548 4586 1552
rect 4710 1548 4714 1552
rect 4758 1548 4762 1552
rect 4790 1548 4794 1552
rect 5038 1548 5042 1552
rect 5062 1548 5066 1552
rect 5094 1548 5098 1552
rect 5158 1548 5162 1552
rect 5230 1548 5234 1552
rect 3550 1538 3554 1542
rect 3678 1538 3682 1542
rect 3894 1538 3898 1542
rect 3998 1538 4002 1542
rect 4022 1538 4026 1542
rect 4094 1538 4098 1542
rect 4142 1538 4146 1542
rect 4246 1538 4250 1542
rect 4294 1538 4298 1542
rect 4302 1538 4306 1542
rect 4350 1538 4354 1542
rect 4358 1538 4362 1542
rect 4406 1538 4410 1542
rect 4422 1538 4426 1542
rect 4526 1538 4530 1542
rect 4542 1538 4546 1542
rect 4590 1538 4594 1542
rect 4622 1538 4626 1542
rect 4686 1538 4690 1542
rect 4814 1538 4818 1542
rect 4830 1538 4834 1542
rect 4838 1538 4842 1542
rect 4886 1538 4890 1542
rect 4910 1538 4914 1542
rect 4926 1538 4930 1542
rect 5006 1538 5010 1542
rect 5030 1538 5034 1542
rect 5062 1538 5066 1542
rect 5094 1538 5098 1542
rect 5150 1538 5154 1542
rect 5206 1538 5210 1542
rect 5246 1538 5250 1542
rect 5294 1538 5298 1542
rect 6 1528 10 1532
rect 110 1528 114 1532
rect 158 1528 162 1532
rect 294 1528 298 1532
rect 614 1528 618 1532
rect 686 1528 690 1532
rect 766 1528 770 1532
rect 846 1528 850 1532
rect 982 1528 986 1532
rect 1118 1528 1122 1532
rect 1134 1528 1138 1532
rect 1478 1528 1482 1532
rect 1510 1528 1514 1532
rect 1582 1528 1586 1532
rect 1622 1528 1626 1532
rect 1750 1528 1754 1532
rect 1766 1528 1770 1532
rect 1854 1528 1858 1532
rect 1910 1528 1914 1532
rect 1982 1528 1986 1532
rect 2070 1528 2074 1532
rect 2142 1528 2146 1532
rect 2190 1528 2194 1532
rect 2246 1528 2250 1532
rect 2278 1528 2282 1532
rect 2374 1528 2378 1532
rect 2446 1528 2450 1532
rect 3350 1528 3354 1532
rect 3390 1528 3394 1532
rect 3630 1528 3634 1532
rect 3702 1528 3706 1532
rect 4214 1528 4218 1532
rect 4438 1528 4442 1532
rect 4486 1528 4490 1532
rect 4510 1528 4514 1532
rect 4518 1528 4522 1532
rect 4542 1528 4546 1532
rect 4918 1528 4922 1532
rect 5014 1528 5018 1532
rect 5102 1528 5106 1532
rect 22 1518 26 1522
rect 126 1518 130 1522
rect 206 1518 210 1522
rect 222 1518 226 1522
rect 246 1518 250 1522
rect 494 1518 498 1522
rect 502 1518 506 1522
rect 694 1518 698 1522
rect 782 1518 786 1522
rect 1174 1518 1178 1522
rect 1382 1518 1386 1522
rect 2238 1518 2242 1522
rect 2318 1518 2322 1522
rect 2838 1518 2842 1522
rect 2846 1518 2850 1522
rect 2958 1518 2962 1522
rect 3278 1518 3282 1522
rect 3414 1518 3418 1522
rect 3462 1518 3466 1522
rect 3662 1518 3666 1522
rect 3822 1518 3826 1522
rect 3838 1518 3842 1522
rect 4078 1518 4082 1522
rect 4110 1518 4114 1522
rect 4262 1518 4266 1522
rect 4318 1518 4322 1522
rect 4374 1518 4378 1522
rect 4430 1518 4434 1522
rect 4630 1518 4634 1522
rect 4734 1518 4738 1522
rect 4854 1518 4858 1522
rect 5022 1518 5026 1522
rect 5110 1518 5114 1522
rect 5262 1518 5266 1522
rect 6 1508 10 1512
rect 3918 1508 3922 1512
rect 858 1503 862 1507
rect 865 1503 869 1507
rect 1874 1503 1878 1507
rect 1881 1503 1885 1507
rect 2906 1503 2910 1507
rect 2913 1503 2917 1507
rect 3930 1503 3934 1507
rect 3937 1503 3941 1507
rect 4954 1503 4958 1507
rect 4961 1503 4965 1507
rect 5190 1498 5194 1502
rect 5294 1498 5298 1502
rect 286 1488 290 1492
rect 318 1488 322 1492
rect 462 1488 466 1492
rect 534 1488 538 1492
rect 590 1488 594 1492
rect 718 1488 722 1492
rect 758 1488 762 1492
rect 910 1488 914 1492
rect 1126 1488 1130 1492
rect 1446 1488 1450 1492
rect 1518 1488 1522 1492
rect 1718 1488 1722 1492
rect 1806 1488 1810 1492
rect 1830 1488 1834 1492
rect 1918 1488 1922 1492
rect 1990 1488 1994 1492
rect 2022 1488 2026 1492
rect 2070 1488 2074 1492
rect 2110 1488 2114 1492
rect 2278 1488 2282 1492
rect 2294 1488 2298 1492
rect 2342 1488 2346 1492
rect 2478 1488 2482 1492
rect 2534 1488 2538 1492
rect 2614 1488 2618 1492
rect 2894 1488 2898 1492
rect 3006 1488 3010 1492
rect 3142 1488 3146 1492
rect 3158 1488 3162 1492
rect 3230 1488 3234 1492
rect 3246 1488 3250 1492
rect 3358 1488 3362 1492
rect 3414 1488 3418 1492
rect 3542 1488 3546 1492
rect 3726 1488 3730 1492
rect 3750 1488 3754 1492
rect 3886 1488 3890 1492
rect 3966 1488 3970 1492
rect 4070 1488 4074 1492
rect 4102 1488 4106 1492
rect 4254 1488 4258 1492
rect 4286 1488 4290 1492
rect 4294 1488 4298 1492
rect 4534 1488 4538 1492
rect 4830 1488 4834 1492
rect 4942 1488 4946 1492
rect 5014 1488 5018 1492
rect 5078 1488 5082 1492
rect 5174 1488 5178 1492
rect 5206 1488 5210 1492
rect 6 1478 10 1482
rect 166 1478 170 1482
rect 206 1478 210 1482
rect 310 1478 314 1482
rect 366 1478 370 1482
rect 470 1478 474 1482
rect 478 1478 482 1482
rect 654 1478 658 1482
rect 694 1478 698 1482
rect 734 1478 738 1482
rect 790 1478 794 1482
rect 1158 1478 1162 1482
rect 1278 1478 1282 1482
rect 1286 1478 1290 1482
rect 1302 1478 1306 1482
rect 1526 1478 1530 1482
rect 1686 1478 1690 1482
rect 1710 1478 1714 1482
rect 1782 1478 1786 1482
rect 1814 1478 1818 1482
rect 1870 1478 1874 1482
rect 1894 1478 1898 1482
rect 1910 1478 1914 1482
rect 2030 1478 2034 1482
rect 2102 1478 2106 1482
rect 2182 1478 2186 1482
rect 2214 1478 2218 1482
rect 2486 1478 2490 1482
rect 2670 1478 2674 1482
rect 2710 1478 2714 1482
rect 38 1468 42 1472
rect 70 1468 74 1472
rect 102 1468 106 1472
rect 46 1458 50 1462
rect 94 1458 98 1462
rect 142 1458 146 1462
rect 254 1468 258 1472
rect 302 1468 306 1472
rect 374 1468 378 1472
rect 422 1468 426 1472
rect 550 1468 554 1472
rect 558 1468 562 1472
rect 606 1468 610 1472
rect 686 1468 690 1472
rect 726 1468 730 1472
rect 774 1468 778 1472
rect 878 1468 882 1472
rect 990 1468 994 1472
rect 1110 1468 1114 1472
rect 1206 1468 1210 1472
rect 1222 1468 1226 1472
rect 1238 1468 1242 1472
rect 1334 1468 1338 1472
rect 1342 1468 1346 1472
rect 1390 1468 1394 1472
rect 1398 1468 1402 1472
rect 1462 1468 1466 1472
rect 1470 1468 1474 1472
rect 1510 1468 1514 1472
rect 1542 1468 1546 1472
rect 1582 1468 1586 1472
rect 1726 1468 1730 1472
rect 1742 1468 1746 1472
rect 1758 1468 1762 1472
rect 1774 1468 1778 1472
rect 1822 1468 1826 1472
rect 1838 1468 1842 1472
rect 1862 1468 1866 1472
rect 2926 1478 2930 1482
rect 3014 1478 3018 1482
rect 3182 1478 3186 1482
rect 3198 1478 3202 1482
rect 3350 1478 3354 1482
rect 3422 1478 3426 1482
rect 3518 1478 3522 1482
rect 3542 1478 3546 1482
rect 3574 1478 3578 1482
rect 3606 1478 3610 1482
rect 3630 1478 3634 1482
rect 3646 1478 3650 1482
rect 3790 1478 3794 1482
rect 3950 1478 3954 1482
rect 4006 1478 4010 1482
rect 4094 1478 4098 1482
rect 4358 1478 4362 1482
rect 4374 1478 4378 1482
rect 4414 1478 4418 1482
rect 4510 1478 4514 1482
rect 4542 1478 4546 1482
rect 4574 1478 4578 1482
rect 4582 1478 4586 1482
rect 4750 1478 4754 1482
rect 4814 1478 4818 1482
rect 4854 1478 4858 1482
rect 4894 1478 4898 1482
rect 4926 1478 4930 1482
rect 5054 1478 5058 1482
rect 5086 1478 5090 1482
rect 5142 1478 5146 1482
rect 182 1458 186 1462
rect 206 1458 210 1462
rect 222 1458 226 1462
rect 230 1458 234 1462
rect 334 1458 338 1462
rect 422 1458 426 1462
rect 446 1458 450 1462
rect 454 1458 458 1462
rect 502 1458 506 1462
rect 630 1458 634 1462
rect 646 1458 650 1462
rect 670 1458 674 1462
rect 694 1458 698 1462
rect 734 1458 738 1462
rect 758 1458 762 1462
rect 862 1459 866 1463
rect 974 1459 978 1463
rect 1022 1458 1026 1462
rect 1094 1459 1098 1463
rect 1190 1459 1194 1463
rect 1238 1458 1242 1462
rect 1310 1458 1314 1462
rect 1334 1458 1338 1462
rect 1478 1458 1482 1462
rect 1502 1458 1506 1462
rect 1566 1458 1570 1462
rect 1702 1458 1706 1462
rect 1742 1458 1746 1462
rect 1750 1458 1754 1462
rect 1910 1458 1914 1462
rect 1934 1458 1938 1462
rect 1974 1468 1978 1472
rect 1998 1468 2002 1472
rect 2014 1468 2018 1472
rect 2030 1468 2034 1472
rect 2054 1468 2058 1472
rect 2086 1466 2090 1470
rect 2094 1468 2098 1472
rect 2126 1468 2130 1472
rect 2150 1468 2154 1472
rect 2158 1468 2162 1472
rect 2174 1468 2178 1472
rect 2286 1468 2290 1472
rect 2302 1468 2306 1472
rect 2366 1468 2370 1472
rect 2454 1468 2458 1472
rect 2470 1468 2474 1472
rect 2486 1468 2490 1472
rect 2510 1468 2514 1472
rect 2526 1468 2530 1472
rect 2574 1468 2578 1472
rect 2582 1468 2586 1472
rect 2630 1468 2634 1472
rect 2702 1468 2706 1472
rect 2862 1468 2866 1472
rect 2974 1468 2978 1472
rect 2998 1468 3002 1472
rect 3022 1468 3026 1472
rect 3038 1468 3042 1472
rect 3206 1468 3210 1472
rect 3238 1468 3242 1472
rect 3502 1468 3506 1472
rect 3710 1468 3714 1472
rect 3734 1468 3738 1472
rect 3830 1468 3834 1472
rect 4086 1468 4090 1472
rect 4158 1468 4162 1472
rect 4174 1468 4178 1472
rect 4214 1468 4218 1472
rect 4262 1468 4266 1472
rect 4310 1468 4314 1472
rect 4318 1468 4322 1472
rect 4342 1468 4346 1472
rect 4406 1468 4410 1472
rect 4430 1468 4434 1472
rect 1966 1458 1970 1462
rect 2006 1458 2010 1462
rect 2038 1458 2042 1462
rect 2214 1459 2218 1463
rect 2462 1458 2466 1462
rect 2494 1458 2498 1462
rect 2654 1458 2658 1462
rect 2758 1458 2762 1462
rect 2846 1459 2850 1463
rect 2958 1459 2962 1463
rect 2990 1458 2994 1462
rect 3030 1458 3034 1462
rect 3086 1458 3090 1462
rect 3110 1458 3114 1462
rect 3182 1458 3186 1462
rect 3214 1458 3218 1462
rect 3286 1458 3290 1462
rect 3310 1458 3314 1462
rect 3366 1458 3370 1462
rect 3390 1458 3394 1462
rect 3406 1458 3410 1462
rect 3478 1458 3482 1462
rect 3494 1458 3498 1462
rect 3550 1458 3554 1462
rect 3606 1458 3610 1462
rect 3622 1458 3626 1462
rect 3646 1458 3650 1462
rect 3654 1458 3658 1462
rect 3678 1458 3682 1462
rect 3686 1458 3690 1462
rect 3766 1458 3770 1462
rect 3774 1458 3778 1462
rect 3822 1459 3826 1463
rect 4502 1468 4506 1472
rect 4566 1468 4570 1472
rect 4598 1468 4602 1472
rect 4614 1468 4618 1472
rect 4662 1468 4666 1472
rect 4694 1468 4698 1472
rect 4774 1468 4778 1472
rect 4806 1468 4810 1472
rect 4838 1468 4842 1472
rect 4886 1468 4890 1472
rect 4894 1468 4898 1472
rect 4910 1468 4914 1472
rect 4950 1468 4954 1472
rect 4990 1468 4994 1472
rect 4998 1468 5002 1472
rect 5022 1468 5026 1472
rect 5038 1468 5042 1472
rect 5062 1468 5066 1472
rect 5094 1468 5098 1472
rect 5150 1468 5154 1472
rect 5182 1468 5186 1472
rect 5262 1468 5266 1472
rect 3894 1458 3898 1462
rect 3918 1458 3922 1462
rect 3974 1458 3978 1462
rect 4014 1458 4018 1462
rect 4086 1458 4090 1462
rect 4110 1458 4114 1462
rect 4134 1458 4138 1462
rect 4150 1458 4154 1462
rect 4198 1458 4202 1462
rect 4270 1458 4274 1462
rect 4454 1458 4458 1462
rect 4462 1458 4466 1462
rect 4478 1458 4482 1462
rect 4494 1458 4498 1462
rect 4542 1458 4546 1462
rect 4582 1458 4586 1462
rect 4606 1458 4610 1462
rect 4670 1458 4674 1462
rect 4766 1458 4770 1462
rect 4782 1458 4786 1462
rect 4790 1458 4794 1462
rect 4926 1458 4930 1462
rect 4974 1458 4978 1462
rect 5030 1458 5034 1462
rect 5102 1458 5106 1462
rect 5118 1458 5122 1462
rect 5126 1458 5130 1462
rect 5158 1458 5162 1462
rect 5182 1458 5186 1462
rect 5270 1458 5274 1462
rect 70 1448 74 1452
rect 126 1449 130 1453
rect 198 1448 202 1452
rect 638 1448 642 1452
rect 662 1448 666 1452
rect 758 1448 762 1452
rect 1222 1448 1226 1452
rect 1246 1448 1250 1452
rect 1294 1448 1298 1452
rect 1358 1448 1362 1452
rect 1494 1448 1498 1452
rect 1646 1448 1650 1452
rect 1766 1448 1770 1452
rect 1790 1448 1794 1452
rect 1838 1448 1842 1452
rect 1918 1448 1922 1452
rect 1982 1448 1986 1452
rect 2062 1448 2066 1452
rect 2134 1448 2138 1452
rect 2302 1448 2306 1452
rect 2438 1448 2442 1452
rect 2518 1448 2522 1452
rect 2662 1448 2666 1452
rect 2686 1448 2690 1452
rect 2718 1448 2722 1452
rect 2742 1448 2746 1452
rect 3046 1448 3050 1452
rect 3230 1448 3234 1452
rect 3398 1448 3402 1452
rect 3486 1448 3490 1452
rect 3718 1448 3722 1452
rect 3782 1448 3786 1452
rect 4142 1448 4146 1452
rect 4294 1448 4298 1452
rect 4318 1448 4322 1452
rect 4366 1448 4370 1452
rect 4390 1448 4394 1452
rect 4430 1448 4434 1452
rect 4470 1448 4474 1452
rect 4478 1448 4482 1452
rect 4798 1448 4802 1452
rect 4822 1448 4826 1452
rect 4846 1448 4850 1452
rect 4862 1448 4866 1452
rect 5006 1448 5010 1452
rect 5174 1448 5178 1452
rect 5206 1448 5210 1452
rect 238 1438 242 1442
rect 622 1438 626 1442
rect 694 1438 698 1442
rect 1310 1438 1314 1442
rect 2638 1438 2642 1442
rect 2646 1438 2650 1442
rect 3158 1438 3162 1442
rect 3342 1438 3346 1442
rect 3382 1438 3386 1442
rect 3446 1438 3450 1442
rect 3470 1438 3474 1442
rect 4126 1438 4130 1442
rect 4646 1438 4650 1442
rect 4966 1438 4970 1442
rect 22 1418 26 1422
rect 94 1418 98 1422
rect 230 1418 234 1422
rect 614 1418 618 1422
rect 798 1418 802 1422
rect 1030 1418 1034 1422
rect 1478 1418 1482 1422
rect 2382 1418 2386 1422
rect 2542 1418 2546 1422
rect 2678 1418 2682 1422
rect 2726 1418 2730 1422
rect 3390 1418 3394 1422
rect 3478 1418 3482 1422
rect 4078 1418 4082 1422
rect 4134 1418 4138 1422
rect 4150 1418 4154 1422
rect 4726 1418 4730 1422
rect 5214 1418 5218 1422
rect 346 1403 350 1407
rect 353 1403 357 1407
rect 1370 1403 1374 1407
rect 1377 1403 1381 1407
rect 2394 1403 2398 1407
rect 2401 1403 2405 1407
rect 3418 1403 3422 1407
rect 3425 1403 3429 1407
rect 4442 1403 4446 1407
rect 4449 1403 4453 1407
rect 22 1388 26 1392
rect 70 1388 74 1392
rect 158 1388 162 1392
rect 1182 1388 1186 1392
rect 1206 1388 1210 1392
rect 1646 1388 1650 1392
rect 1758 1388 1762 1392
rect 1798 1388 1802 1392
rect 1926 1388 1930 1392
rect 1950 1388 1954 1392
rect 1982 1388 1986 1392
rect 2022 1388 2026 1392
rect 2174 1388 2178 1392
rect 2222 1388 2226 1392
rect 2278 1388 2282 1392
rect 2302 1388 2306 1392
rect 2334 1388 2338 1392
rect 2534 1388 2538 1392
rect 2790 1388 2794 1392
rect 3182 1388 3186 1392
rect 3310 1388 3314 1392
rect 3534 1388 3538 1392
rect 3558 1388 3562 1392
rect 3654 1388 3658 1392
rect 3846 1388 3850 1392
rect 4046 1388 4050 1392
rect 4142 1388 4146 1392
rect 4150 1388 4154 1392
rect 4358 1388 4362 1392
rect 4470 1388 4474 1392
rect 4558 1388 4562 1392
rect 4822 1388 4826 1392
rect 4846 1388 4850 1392
rect 4998 1388 5002 1392
rect 5054 1388 5058 1392
rect 5110 1388 5114 1392
rect 5246 1388 5250 1392
rect 5278 1388 5282 1392
rect 1006 1378 1010 1382
rect 1830 1378 1834 1382
rect 1910 1378 1914 1382
rect 2070 1378 2074 1382
rect 2238 1378 2242 1382
rect 2678 1378 2682 1382
rect 4502 1378 4506 1382
rect 30 1368 34 1372
rect 38 1368 42 1372
rect 62 1368 66 1372
rect 390 1368 394 1372
rect 430 1368 434 1372
rect 438 1368 442 1372
rect 822 1368 826 1372
rect 838 1368 842 1372
rect 846 1368 850 1372
rect 950 1368 954 1372
rect 974 1368 978 1372
rect 1014 1368 1018 1372
rect 1110 1368 1114 1372
rect 1126 1368 1130 1372
rect 1382 1368 1386 1372
rect 1934 1368 1938 1372
rect 2030 1368 2034 1372
rect 2246 1368 2250 1372
rect 2342 1368 2346 1372
rect 2806 1368 2810 1372
rect 2942 1368 2946 1372
rect 4478 1368 4482 1372
rect 4510 1368 4514 1372
rect 4646 1368 4650 1372
rect 4702 1368 4706 1372
rect 4758 1368 4762 1372
rect 4854 1368 4858 1372
rect 5214 1368 5218 1372
rect 5230 1368 5234 1372
rect 5238 1368 5242 1372
rect 5286 1368 5290 1372
rect 38 1358 42 1362
rect 78 1358 82 1362
rect 254 1358 258 1362
rect 302 1358 306 1362
rect 310 1358 314 1362
rect 414 1358 418 1362
rect 422 1358 426 1362
rect 454 1358 458 1362
rect 462 1358 466 1362
rect 486 1358 490 1362
rect 558 1358 562 1362
rect 598 1358 602 1362
rect 614 1358 618 1362
rect 806 1358 810 1362
rect 870 1358 874 1362
rect 894 1358 898 1362
rect 990 1358 994 1362
rect 998 1358 1002 1362
rect 1030 1358 1034 1362
rect 1054 1358 1058 1362
rect 1070 1358 1074 1362
rect 1150 1358 1154 1362
rect 1918 1358 1922 1362
rect 2046 1358 2050 1362
rect 2110 1358 2114 1362
rect 2190 1358 2194 1362
rect 2262 1358 2266 1362
rect 2286 1358 2290 1362
rect 2318 1358 2322 1362
rect 2838 1358 2842 1362
rect 2854 1358 2858 1362
rect 2862 1358 2866 1362
rect 2902 1358 2906 1362
rect 2926 1358 2930 1362
rect 2982 1358 2986 1362
rect 3062 1358 3066 1362
rect 3646 1358 3650 1362
rect 3750 1358 3754 1362
rect 3806 1358 3810 1362
rect 4182 1358 4186 1362
rect 4222 1358 4226 1362
rect 4294 1358 4298 1362
rect 4494 1358 4498 1362
rect 4550 1358 4554 1362
rect 4590 1358 4594 1362
rect 4838 1358 4842 1362
rect 4870 1358 4874 1362
rect 5006 1358 5010 1362
rect 5014 1358 5018 1362
rect 5062 1358 5066 1362
rect 5182 1358 5186 1362
rect 5238 1358 5242 1362
rect 5270 1358 5274 1362
rect 22 1348 26 1352
rect 70 1348 74 1352
rect 94 1348 98 1352
rect 110 1348 114 1352
rect 134 1348 138 1352
rect 198 1348 202 1352
rect 222 1348 226 1352
rect 286 1348 290 1352
rect 350 1348 354 1352
rect 366 1348 370 1352
rect 382 1348 386 1352
rect 398 1348 402 1352
rect 446 1348 450 1352
rect 462 1348 466 1352
rect 526 1348 530 1352
rect 542 1348 546 1352
rect 574 1348 578 1352
rect 606 1348 610 1352
rect 670 1348 674 1352
rect 846 1348 850 1352
rect 918 1348 922 1352
rect 982 1348 986 1352
rect 1006 1348 1010 1352
rect 1054 1348 1058 1352
rect 1126 1348 1130 1352
rect 1166 1348 1170 1352
rect 1326 1348 1330 1352
rect 1438 1348 1442 1352
rect 1542 1348 1546 1352
rect 1582 1348 1586 1352
rect 102 1338 106 1342
rect 214 1338 218 1342
rect 230 1338 234 1342
rect 270 1338 274 1342
rect 278 1338 282 1342
rect 358 1338 362 1342
rect 478 1338 482 1342
rect 550 1338 554 1342
rect 582 1338 586 1342
rect 630 1338 634 1342
rect 638 1338 642 1342
rect 686 1338 690 1342
rect 694 1338 698 1342
rect 742 1338 746 1342
rect 750 1338 754 1342
rect 822 1338 826 1342
rect 926 1338 930 1342
rect 966 1338 970 1342
rect 1046 1338 1050 1342
rect 1614 1347 1618 1351
rect 1678 1348 1682 1352
rect 1710 1347 1714 1351
rect 1886 1348 1890 1352
rect 1926 1348 1930 1352
rect 2038 1348 2042 1352
rect 2134 1348 2138 1352
rect 2142 1348 2146 1352
rect 2174 1348 2178 1352
rect 2198 1348 2202 1352
rect 2214 1348 2218 1352
rect 2254 1348 2258 1352
rect 2318 1348 2322 1352
rect 2350 1348 2354 1352
rect 2398 1348 2402 1352
rect 2414 1348 2418 1352
rect 2734 1348 2738 1352
rect 2790 1348 2794 1352
rect 2838 1348 2842 1352
rect 2870 1348 2874 1352
rect 3022 1348 3026 1352
rect 3102 1348 3106 1352
rect 3142 1348 3146 1352
rect 3174 1348 3178 1352
rect 3190 1348 3194 1352
rect 1070 1338 1074 1342
rect 1118 1338 1122 1342
rect 1174 1338 1178 1342
rect 1262 1338 1266 1342
rect 1318 1338 1322 1342
rect 1462 1338 1466 1342
rect 1478 1338 1482 1342
rect 1630 1338 1634 1342
rect 1742 1338 1746 1342
rect 1790 1338 1794 1342
rect 1814 1338 1818 1342
rect 1870 1338 1874 1342
rect 1894 1338 1898 1342
rect 1966 1338 1970 1342
rect 2014 1338 2018 1342
rect 2054 1338 2058 1342
rect 2102 1338 2106 1342
rect 2118 1338 2122 1342
rect 2142 1338 2146 1342
rect 2230 1338 2234 1342
rect 2310 1338 2314 1342
rect 2422 1338 2426 1342
rect 2470 1338 2474 1342
rect 2478 1338 2482 1342
rect 2526 1338 2530 1342
rect 2550 1338 2554 1342
rect 2598 1338 2602 1342
rect 2606 1338 2610 1342
rect 2654 1338 2658 1342
rect 2662 1338 2666 1342
rect 2718 1338 2722 1342
rect 2726 1338 2730 1342
rect 2782 1338 2786 1342
rect 2830 1338 2834 1342
rect 2886 1338 2890 1342
rect 2942 1338 2946 1342
rect 2966 1338 2970 1342
rect 2982 1338 2986 1342
rect 2998 1338 3002 1342
rect 3046 1338 3050 1342
rect 3062 1338 3066 1342
rect 3246 1347 3250 1351
rect 3358 1348 3362 1352
rect 3430 1348 3434 1352
rect 3478 1348 3482 1352
rect 3590 1348 3594 1352
rect 3622 1348 3626 1352
rect 3718 1347 3722 1351
rect 3766 1348 3770 1352
rect 3790 1348 3794 1352
rect 3822 1348 3826 1352
rect 3886 1348 3890 1352
rect 3982 1347 3986 1351
rect 4014 1348 4018 1352
rect 4102 1348 4106 1352
rect 4166 1348 4170 1352
rect 4198 1348 4202 1352
rect 4214 1348 4218 1352
rect 4262 1348 4266 1352
rect 4278 1348 4282 1352
rect 4302 1348 4306 1352
rect 4326 1348 4330 1352
rect 4342 1348 4346 1352
rect 4350 1348 4354 1352
rect 4414 1348 4418 1352
rect 4486 1348 4490 1352
rect 4630 1348 4634 1352
rect 4798 1348 4802 1352
rect 4846 1348 4850 1352
rect 4902 1348 4906 1352
rect 5014 1348 5018 1352
rect 5030 1348 5034 1352
rect 5086 1348 5090 1352
rect 5158 1348 5162 1352
rect 5246 1348 5250 1352
rect 5278 1348 5282 1352
rect 3150 1338 3154 1342
rect 3454 1338 3458 1342
rect 3550 1338 3554 1342
rect 3598 1338 3602 1342
rect 3734 1338 3738 1342
rect 3774 1338 3778 1342
rect 3782 1338 3786 1342
rect 3830 1338 3834 1342
rect 3894 1338 3898 1342
rect 4086 1338 4090 1342
rect 4214 1338 4218 1342
rect 4254 1338 4258 1342
rect 4270 1338 4274 1342
rect 4310 1338 4314 1342
rect 4334 1338 4338 1342
rect 4534 1338 4538 1342
rect 4574 1338 4578 1342
rect 4606 1338 4610 1342
rect 4678 1338 4682 1342
rect 4686 1338 4690 1342
rect 4734 1338 4738 1342
rect 4742 1338 4746 1342
rect 4790 1338 4794 1342
rect 4886 1338 4890 1342
rect 4926 1338 4930 1342
rect 4974 1338 4978 1342
rect 5102 1338 5106 1342
rect 5150 1338 5154 1342
rect 5158 1338 5162 1342
rect 5182 1338 5186 1342
rect 5198 1338 5202 1342
rect 38 1328 42 1332
rect 86 1328 90 1332
rect 118 1328 122 1332
rect 134 1328 138 1332
rect 214 1328 218 1332
rect 310 1328 314 1332
rect 374 1328 378 1332
rect 414 1328 418 1332
rect 518 1328 522 1332
rect 886 1328 890 1332
rect 894 1328 898 1332
rect 942 1328 946 1332
rect 950 1328 954 1332
rect 1086 1328 1090 1332
rect 1142 1328 1146 1332
rect 1190 1328 1194 1332
rect 1806 1328 1810 1332
rect 1910 1328 1914 1332
rect 1958 1328 1962 1332
rect 2158 1328 2162 1332
rect 2198 1328 2202 1332
rect 2270 1328 2274 1332
rect 2318 1328 2322 1332
rect 2374 1328 2378 1332
rect 2382 1328 2386 1332
rect 2390 1328 2394 1332
rect 2542 1328 2546 1332
rect 2750 1328 2754 1332
rect 2774 1328 2778 1332
rect 2822 1328 2826 1332
rect 2902 1328 2906 1332
rect 2918 1328 2922 1332
rect 2982 1328 2986 1332
rect 3014 1328 3018 1332
rect 3094 1328 3098 1332
rect 3118 1328 3122 1332
rect 3190 1328 3194 1332
rect 3246 1328 3250 1332
rect 3342 1328 3346 1332
rect 3558 1328 3562 1332
rect 3566 1328 3570 1332
rect 3606 1328 3610 1332
rect 4230 1328 4234 1332
rect 4238 1328 4242 1332
rect 4294 1328 4298 1332
rect 4334 1328 4338 1332
rect 4422 1328 4426 1332
rect 4510 1328 4514 1332
rect 4598 1328 4602 1332
rect 4830 1328 4834 1332
rect 4894 1328 4898 1332
rect 5046 1328 5050 1332
rect 5062 1328 5066 1332
rect 5134 1328 5138 1332
rect 5190 1328 5194 1332
rect 5230 1328 5234 1332
rect 238 1318 242 1322
rect 302 1318 306 1322
rect 494 1318 498 1322
rect 558 1318 562 1322
rect 614 1318 618 1322
rect 710 1318 714 1322
rect 766 1318 770 1322
rect 934 1318 938 1322
rect 1030 1318 1034 1322
rect 1150 1318 1154 1322
rect 1270 1318 1274 1322
rect 1550 1318 1554 1322
rect 2486 1318 2490 1322
rect 2502 1318 2506 1322
rect 2566 1318 2570 1322
rect 2622 1318 2626 1322
rect 2766 1318 2770 1322
rect 3006 1318 3010 1322
rect 3054 1318 3058 1322
rect 3110 1318 3114 1322
rect 3126 1318 3130 1322
rect 3542 1318 3546 1322
rect 3574 1318 3578 1322
rect 3646 1318 3650 1322
rect 4246 1318 4250 1322
rect 4942 1318 4946 1322
rect 5070 1318 5074 1322
rect 5246 1318 5250 1322
rect 1278 1308 1282 1312
rect 2590 1308 2594 1312
rect 858 1303 862 1307
rect 865 1303 869 1307
rect 1874 1303 1878 1307
rect 1881 1303 1885 1307
rect 2906 1303 2910 1307
rect 2913 1303 2917 1307
rect 3930 1303 3934 1307
rect 3937 1303 3941 1307
rect 4954 1303 4958 1307
rect 4961 1303 4965 1307
rect 14 1288 18 1292
rect 38 1288 42 1292
rect 70 1288 74 1292
rect 110 1288 114 1292
rect 190 1288 194 1292
rect 230 1288 234 1292
rect 310 1288 314 1292
rect 390 1288 394 1292
rect 478 1288 482 1292
rect 558 1288 562 1292
rect 638 1288 642 1292
rect 678 1288 682 1292
rect 814 1288 818 1292
rect 1030 1288 1034 1292
rect 1310 1288 1314 1292
rect 1422 1288 1426 1292
rect 1638 1288 1642 1292
rect 1718 1288 1722 1292
rect 1734 1288 1738 1292
rect 1918 1288 1922 1292
rect 1926 1288 1930 1292
rect 1942 1288 1946 1292
rect 2126 1288 2130 1292
rect 2182 1288 2186 1292
rect 2294 1288 2298 1292
rect 2470 1288 2474 1292
rect 2630 1288 2634 1292
rect 2686 1288 2690 1292
rect 2798 1288 2802 1292
rect 3638 1288 3642 1292
rect 3830 1288 3834 1292
rect 3966 1288 3970 1292
rect 4102 1288 4106 1292
rect 4238 1288 4242 1292
rect 4318 1288 4322 1292
rect 4382 1288 4386 1292
rect 4638 1288 4642 1292
rect 4694 1288 4698 1292
rect 4846 1288 4850 1292
rect 4870 1288 4874 1292
rect 4982 1288 4986 1292
rect 5142 1288 5146 1292
rect 5166 1288 5170 1292
rect 5222 1288 5226 1292
rect 5278 1288 5282 1292
rect 94 1278 98 1282
rect 222 1278 226 1282
rect 294 1278 298 1282
rect 446 1278 450 1282
rect 494 1278 498 1282
rect 526 1278 530 1282
rect 758 1278 762 1282
rect 766 1278 770 1282
rect 782 1278 786 1282
rect 830 1278 834 1282
rect 886 1278 890 1282
rect 950 1278 954 1282
rect 982 1278 986 1282
rect 1062 1278 1066 1282
rect 1086 1278 1090 1282
rect 1174 1278 1178 1282
rect 1222 1278 1226 1282
rect 1342 1278 1346 1282
rect 1374 1278 1378 1282
rect 1542 1278 1546 1282
rect 1550 1278 1554 1282
rect 1590 1278 1594 1282
rect 1670 1278 1674 1282
rect 1686 1278 1690 1282
rect 1726 1278 1730 1282
rect 1758 1278 1762 1282
rect 1846 1278 1850 1282
rect 1854 1278 1858 1282
rect 1934 1278 1938 1282
rect 2094 1278 2098 1282
rect 2110 1278 2114 1282
rect 2118 1278 2122 1282
rect 2158 1278 2162 1282
rect 2174 1278 2178 1282
rect 2302 1278 2306 1282
rect 2806 1278 2810 1282
rect 2814 1278 2818 1282
rect 2846 1278 2850 1282
rect 2854 1278 2858 1282
rect 2862 1278 2866 1282
rect 2910 1278 2914 1282
rect 3094 1278 3098 1282
rect 3102 1278 3106 1282
rect 3262 1278 3266 1282
rect 3470 1278 3474 1282
rect 3486 1278 3490 1282
rect 3566 1278 3570 1282
rect 3678 1278 3682 1282
rect 3798 1278 3802 1282
rect 3894 1278 3898 1282
rect 3958 1278 3962 1282
rect 4030 1278 4034 1282
rect 4094 1278 4098 1282
rect 4230 1278 4234 1282
rect 4254 1278 4258 1282
rect 4350 1278 4354 1282
rect 6 1268 10 1272
rect 22 1268 26 1272
rect 54 1268 58 1272
rect 102 1268 106 1272
rect 118 1268 122 1272
rect 134 1268 138 1272
rect 214 1268 218 1272
rect 238 1268 242 1272
rect 318 1268 322 1272
rect 342 1268 346 1272
rect 430 1268 434 1272
rect 454 1268 458 1272
rect 494 1268 498 1272
rect 510 1268 514 1272
rect 542 1268 546 1272
rect 590 1268 594 1272
rect 622 1268 626 1272
rect 670 1268 674 1272
rect 702 1268 706 1272
rect 750 1268 754 1272
rect 790 1268 794 1272
rect 838 1268 842 1272
rect 854 1268 858 1272
rect 878 1268 882 1272
rect 966 1268 970 1272
rect 998 1268 1002 1272
rect 1014 1268 1018 1272
rect 1046 1268 1050 1272
rect 1086 1268 1090 1272
rect 1206 1268 1210 1272
rect 1254 1268 1258 1272
rect 1286 1268 1290 1272
rect 1326 1268 1330 1272
rect 1342 1268 1346 1272
rect 1406 1268 1410 1272
rect 1462 1268 1466 1272
rect 1478 1268 1482 1272
rect 1518 1268 1522 1272
rect 1590 1268 1594 1272
rect 1614 1268 1618 1272
rect 1654 1268 1658 1272
rect 1670 1268 1674 1272
rect 1694 1268 1698 1272
rect 1742 1268 1746 1272
rect 1782 1268 1786 1272
rect 1790 1268 1794 1272
rect 1838 1268 1842 1272
rect 1862 1268 1866 1272
rect 1894 1268 1898 1272
rect 2022 1268 2026 1272
rect 14 1258 18 1262
rect 110 1258 114 1262
rect 142 1258 146 1262
rect 246 1258 250 1262
rect 262 1258 266 1262
rect 326 1258 330 1262
rect 358 1258 362 1262
rect 406 1258 410 1262
rect 422 1258 426 1262
rect 462 1258 466 1262
rect 486 1258 490 1262
rect 526 1258 530 1262
rect 614 1258 618 1262
rect 694 1258 698 1262
rect 726 1258 730 1262
rect 742 1258 746 1262
rect 774 1258 778 1262
rect 798 1258 802 1262
rect 846 1258 850 1262
rect 902 1258 906 1262
rect 942 1258 946 1262
rect 966 1258 970 1262
rect 990 1258 994 1262
rect 1022 1258 1026 1262
rect 1062 1258 1066 1262
rect 1118 1258 1122 1262
rect 1142 1258 1146 1262
rect 1198 1258 1202 1262
rect 1206 1258 1210 1262
rect 1230 1258 1234 1262
rect 1246 1258 1250 1262
rect 1278 1258 1282 1262
rect 1294 1258 1298 1262
rect 1310 1258 1314 1262
rect 1334 1258 1338 1262
rect 1398 1258 1402 1262
rect 1510 1258 1514 1262
rect 1518 1258 1522 1262
rect 1558 1258 1562 1262
rect 1574 1258 1578 1262
rect 1606 1258 1610 1262
rect 1622 1258 1626 1262
rect 1638 1258 1642 1262
rect 1662 1258 1666 1262
rect 1702 1258 1706 1262
rect 1750 1258 1754 1262
rect 1774 1258 1778 1262
rect 1822 1258 1826 1262
rect 1870 1258 1874 1262
rect 1902 1258 1906 1262
rect 2006 1259 2010 1263
rect 2038 1258 2042 1262
rect 2054 1258 2058 1262
rect 2078 1268 2082 1272
rect 2094 1268 2098 1272
rect 2134 1268 2138 1272
rect 2142 1268 2146 1272
rect 2190 1268 2194 1272
rect 2198 1268 2202 1272
rect 2246 1268 2250 1272
rect 2286 1268 2290 1272
rect 2302 1268 2306 1272
rect 2326 1268 2330 1272
rect 2390 1268 2394 1272
rect 2614 1268 2618 1272
rect 2662 1268 2666 1272
rect 2678 1268 2682 1272
rect 2718 1268 2722 1272
rect 2726 1268 2730 1272
rect 2774 1268 2778 1272
rect 2790 1268 2794 1272
rect 2814 1268 2818 1272
rect 2870 1268 2874 1272
rect 2902 1268 2906 1272
rect 2982 1268 2986 1272
rect 3126 1268 3130 1272
rect 3150 1268 3154 1272
rect 3246 1268 3250 1272
rect 3342 1268 3346 1272
rect 3366 1268 3370 1272
rect 3454 1268 3458 1272
rect 3542 1268 3546 1272
rect 3566 1268 3570 1272
rect 3582 1268 3586 1272
rect 3590 1268 3594 1272
rect 3646 1268 3650 1272
rect 3678 1268 3682 1272
rect 3702 1268 3706 1272
rect 3718 1268 3722 1272
rect 4654 1278 4658 1282
rect 4798 1278 4802 1282
rect 5158 1278 5162 1282
rect 4198 1268 4202 1272
rect 4270 1268 4274 1272
rect 4278 1268 4282 1272
rect 4342 1268 4346 1272
rect 4366 1268 4370 1272
rect 4422 1268 4426 1272
rect 4430 1268 4434 1272
rect 4494 1268 4498 1272
rect 4542 1268 4546 1272
rect 4574 1268 4578 1272
rect 4646 1268 4650 1272
rect 2070 1258 2074 1262
rect 2086 1258 2090 1262
rect 2254 1258 2258 1262
rect 2278 1258 2282 1262
rect 2310 1258 2314 1262
rect 2342 1258 2346 1262
rect 2406 1259 2410 1263
rect 2526 1258 2530 1262
rect 2558 1259 2562 1263
rect 2590 1258 2594 1262
rect 2670 1258 2674 1262
rect 2758 1258 2762 1262
rect 2782 1258 2786 1262
rect 2878 1258 2882 1262
rect 2950 1258 2954 1262
rect 2966 1258 2970 1262
rect 2998 1258 3002 1262
rect 3038 1258 3042 1262
rect 3070 1258 3074 1262
rect 3118 1258 3122 1262
rect 3230 1259 3234 1263
rect 3294 1258 3298 1262
rect 3318 1258 3322 1262
rect 3390 1258 3394 1262
rect 3414 1258 3418 1262
rect 3502 1258 3506 1262
rect 3526 1258 3530 1262
rect 3550 1258 3554 1262
rect 3558 1258 3562 1262
rect 3590 1258 3594 1262
rect 3614 1258 3618 1262
rect 3622 1258 3626 1262
rect 3654 1258 3658 1262
rect 3686 1258 3690 1262
rect 3694 1258 3698 1262
rect 3790 1258 3794 1262
rect 3894 1259 3898 1263
rect 4710 1268 4714 1272
rect 4718 1268 4722 1272
rect 4766 1268 4770 1272
rect 4774 1268 4778 1272
rect 4790 1268 4794 1272
rect 4806 1268 4810 1272
rect 4830 1268 4834 1272
rect 4846 1268 4850 1272
rect 4902 1268 4906 1272
rect 4910 1268 4914 1272
rect 4974 1268 4978 1272
rect 5014 1268 5018 1272
rect 5078 1268 5082 1272
rect 5126 1268 5130 1272
rect 5134 1268 5138 1272
rect 5206 1268 5210 1272
rect 5270 1268 5274 1272
rect 5302 1268 5306 1272
rect 3942 1258 3946 1262
rect 3958 1258 3962 1262
rect 4014 1258 4018 1262
rect 4062 1258 4066 1262
rect 4190 1258 4194 1262
rect 4254 1258 4258 1262
rect 4262 1258 4266 1262
rect 4334 1258 4338 1262
rect 4358 1258 4362 1262
rect 4438 1258 4442 1262
rect 4510 1258 4514 1262
rect 4582 1258 4586 1262
rect 4662 1258 4666 1262
rect 4830 1258 4834 1262
rect 5022 1258 5026 1262
rect 5062 1258 5066 1262
rect 5078 1258 5082 1262
rect 5174 1258 5178 1262
rect 5182 1258 5186 1262
rect 5206 1258 5210 1262
rect 5222 1258 5226 1262
rect 5270 1258 5274 1262
rect 30 1248 34 1252
rect 38 1248 42 1252
rect 62 1248 66 1252
rect 78 1248 82 1252
rect 126 1248 130 1252
rect 158 1248 162 1252
rect 254 1248 258 1252
rect 294 1248 298 1252
rect 350 1248 354 1252
rect 398 1248 402 1252
rect 406 1248 410 1252
rect 702 1248 706 1252
rect 734 1248 738 1252
rect 862 1248 866 1252
rect 926 1248 930 1252
rect 998 1248 1002 1252
rect 1030 1248 1034 1252
rect 1054 1248 1058 1252
rect 1126 1248 1130 1252
rect 1134 1248 1138 1252
rect 1222 1248 1226 1252
rect 1310 1248 1314 1252
rect 1478 1248 1482 1252
rect 1534 1248 1538 1252
rect 1550 1248 1554 1252
rect 1598 1248 1602 1252
rect 1638 1248 1642 1252
rect 1758 1248 1762 1252
rect 2038 1248 2042 1252
rect 2334 1248 2338 1252
rect 2702 1248 2706 1252
rect 2734 1248 2738 1252
rect 2750 1248 2754 1252
rect 2758 1248 2762 1252
rect 2886 1248 2890 1252
rect 2958 1248 2962 1252
rect 2966 1248 2970 1252
rect 2982 1248 2986 1252
rect 3022 1248 3026 1252
rect 3046 1248 3050 1252
rect 3158 1248 3162 1252
rect 3534 1248 3538 1252
rect 3614 1248 3618 1252
rect 3710 1248 3714 1252
rect 4150 1248 4154 1252
rect 4318 1248 4322 1252
rect 4790 1248 4794 1252
rect 4846 1248 4850 1252
rect 4998 1248 5002 1252
rect 5070 1248 5074 1252
rect 5150 1248 5154 1252
rect 5182 1248 5186 1252
rect 5214 1248 5218 1252
rect 5246 1248 5250 1252
rect 5262 1248 5266 1252
rect 5278 1248 5282 1252
rect 270 1238 274 1242
rect 342 1238 346 1242
rect 718 1238 722 1242
rect 1070 1238 1074 1242
rect 1142 1238 1146 1242
rect 1150 1238 1154 1242
rect 2174 1238 2178 1242
rect 2214 1238 2218 1242
rect 2454 1238 2458 1242
rect 2942 1238 2946 1242
rect 3006 1238 3010 1242
rect 3030 1238 3034 1242
rect 3062 1238 3066 1242
rect 4750 1238 4754 1242
rect 5054 1238 5058 1242
rect 5230 1238 5234 1242
rect 262 1228 266 1232
rect 1102 1228 1106 1232
rect 1166 1228 1170 1232
rect 3054 1228 3058 1232
rect 5062 1228 5066 1232
rect 438 1218 442 1222
rect 534 1218 538 1222
rect 1142 1218 1146 1222
rect 1198 1218 1202 1222
rect 1294 1218 1298 1222
rect 1470 1218 1474 1222
rect 1494 1218 1498 1222
rect 1926 1218 1930 1222
rect 2166 1218 2170 1222
rect 2478 1218 2482 1222
rect 2918 1218 2922 1222
rect 2998 1218 3002 1222
rect 3478 1218 3482 1222
rect 3502 1218 3506 1222
rect 3638 1218 3642 1222
rect 4118 1218 4122 1222
rect 4302 1218 4306 1222
rect 346 1203 350 1207
rect 353 1203 357 1207
rect 1370 1203 1374 1207
rect 1377 1203 1381 1207
rect 2394 1203 2398 1207
rect 2401 1203 2405 1207
rect 3418 1203 3422 1207
rect 3425 1203 3429 1207
rect 4442 1203 4446 1207
rect 4449 1203 4453 1207
rect 22 1188 26 1192
rect 46 1188 50 1192
rect 118 1188 122 1192
rect 158 1188 162 1192
rect 214 1188 218 1192
rect 310 1188 314 1192
rect 334 1188 338 1192
rect 606 1188 610 1192
rect 710 1188 714 1192
rect 806 1188 810 1192
rect 1758 1188 1762 1192
rect 1782 1188 1786 1192
rect 1838 1188 1842 1192
rect 1854 1188 1858 1192
rect 1910 1188 1914 1192
rect 1958 1188 1962 1192
rect 2134 1188 2138 1192
rect 2286 1188 2290 1192
rect 2366 1188 2370 1192
rect 2462 1188 2466 1192
rect 2494 1188 2498 1192
rect 2518 1188 2522 1192
rect 2638 1188 2642 1192
rect 2710 1188 2714 1192
rect 2750 1188 2754 1192
rect 2902 1188 2906 1192
rect 3006 1188 3010 1192
rect 3102 1188 3106 1192
rect 3334 1188 3338 1192
rect 3934 1188 3938 1192
rect 4190 1188 4194 1192
rect 4254 1188 4258 1192
rect 4846 1188 4850 1192
rect 4886 1188 4890 1192
rect 4934 1188 4938 1192
rect 5014 1188 5018 1192
rect 5102 1188 5106 1192
rect 5142 1188 5146 1192
rect 5206 1188 5210 1192
rect 2414 1178 2418 1182
rect 4502 1178 4506 1182
rect 142 1168 146 1172
rect 150 1168 154 1172
rect 302 1168 306 1172
rect 510 1168 514 1172
rect 758 1168 762 1172
rect 814 1168 818 1172
rect 1270 1168 1274 1172
rect 1598 1168 1602 1172
rect 1614 1168 1618 1172
rect 1830 1168 1834 1172
rect 2486 1168 2490 1172
rect 2742 1168 2746 1172
rect 3630 1168 3634 1172
rect 4238 1168 4242 1172
rect 4806 1168 4810 1172
rect 4894 1168 4898 1172
rect 5094 1168 5098 1172
rect 5246 1168 5250 1172
rect 126 1158 130 1162
rect 134 1158 138 1162
rect 174 1158 178 1162
rect 254 1158 258 1162
rect 318 1158 322 1162
rect 550 1158 554 1162
rect 622 1158 626 1162
rect 654 1158 658 1162
rect 678 1158 682 1162
rect 726 1158 730 1162
rect 742 1158 746 1162
rect 830 1158 834 1162
rect 1094 1158 1098 1162
rect 1398 1158 1402 1162
rect 1454 1158 1458 1162
rect 1630 1158 1634 1162
rect 1670 1158 1674 1162
rect 1798 1158 1802 1162
rect 1846 1158 1850 1162
rect 1886 1158 1890 1162
rect 1902 1158 1906 1162
rect 1926 1158 1930 1162
rect 2070 1158 2074 1162
rect 2262 1158 2266 1162
rect 2342 1158 2346 1162
rect 2470 1158 2474 1162
rect 2558 1158 2562 1162
rect 2614 1158 2618 1162
rect 2686 1158 2690 1162
rect 2694 1158 2698 1162
rect 2726 1158 2730 1162
rect 2950 1158 2954 1162
rect 86 1148 90 1152
rect 118 1148 122 1152
rect 142 1148 146 1152
rect 166 1148 170 1152
rect 238 1148 242 1152
rect 246 1148 250 1152
rect 286 1148 290 1152
rect 310 1148 314 1152
rect 414 1148 418 1152
rect 470 1148 474 1152
rect 566 1148 570 1152
rect 606 1148 610 1152
rect 646 1148 650 1152
rect 710 1148 714 1152
rect 734 1148 738 1152
rect 798 1148 802 1152
rect 822 1148 826 1152
rect 1030 1147 1034 1151
rect 1086 1148 1090 1152
rect 1134 1148 1138 1152
rect 1238 1147 1242 1151
rect 1302 1148 1306 1152
rect 1334 1147 1338 1151
rect 1438 1148 1442 1152
rect 1622 1148 1626 1152
rect 1638 1148 1642 1152
rect 1710 1148 1714 1152
rect 1726 1148 1730 1152
rect 1774 1148 1778 1152
rect 1838 1148 1842 1152
rect 1942 1148 1946 1152
rect 1982 1148 1986 1152
rect 1990 1148 1994 1152
rect 2054 1148 2058 1152
rect 2086 1148 2090 1152
rect 2134 1148 2138 1152
rect 2182 1148 2186 1152
rect 2206 1148 2210 1152
rect 2230 1148 2234 1152
rect 2446 1148 2450 1152
rect 2478 1148 2482 1152
rect 2574 1148 2578 1152
rect 2622 1148 2626 1152
rect 22 1138 26 1142
rect 78 1138 82 1142
rect 230 1138 234 1142
rect 278 1138 282 1142
rect 358 1138 362 1142
rect 406 1138 410 1142
rect 438 1138 442 1142
rect 486 1138 490 1142
rect 494 1138 498 1142
rect 550 1138 554 1142
rect 566 1138 570 1142
rect 598 1138 602 1142
rect 654 1138 658 1142
rect 702 1138 706 1142
rect 774 1138 778 1142
rect 790 1138 794 1142
rect 902 1138 906 1142
rect 910 1138 914 1142
rect 958 1138 962 1142
rect 1022 1138 1026 1142
rect 1078 1138 1082 1142
rect 1110 1138 1114 1142
rect 1158 1140 1162 1144
rect 1166 1138 1170 1142
rect 1406 1138 1410 1142
rect 1422 1138 1426 1142
rect 1446 1138 1450 1142
rect 1462 1138 1466 1142
rect 1510 1138 1514 1142
rect 1518 1138 1522 1142
rect 1566 1138 1570 1142
rect 1582 1138 1586 1142
rect 1646 1138 1650 1142
rect 1670 1138 1674 1142
rect 1686 1138 1690 1142
rect 2686 1148 2690 1152
rect 2710 1148 2714 1152
rect 2734 1148 2738 1152
rect 2782 1148 2786 1152
rect 2822 1148 2826 1152
rect 2942 1148 2946 1152
rect 3062 1148 3066 1152
rect 3134 1148 3138 1152
rect 3142 1148 3146 1152
rect 3198 1148 3202 1152
rect 3294 1148 3298 1152
rect 3326 1148 3330 1152
rect 1798 1138 1802 1142
rect 1814 1138 1818 1142
rect 1870 1138 1874 1142
rect 1918 1138 1922 1142
rect 1934 1138 1938 1142
rect 1950 1138 1954 1142
rect 1974 1138 1978 1142
rect 1990 1138 1994 1142
rect 2038 1138 2042 1142
rect 2046 1138 2050 1142
rect 2094 1138 2098 1142
rect 2102 1138 2106 1142
rect 2126 1138 2130 1142
rect 2142 1138 2146 1142
rect 2174 1138 2178 1142
rect 2246 1138 2250 1142
rect 2270 1138 2274 1142
rect 2326 1138 2330 1142
rect 2398 1138 2402 1142
rect 2438 1138 2442 1142
rect 2454 1138 2458 1142
rect 2502 1138 2506 1142
rect 2590 1138 2594 1142
rect 2638 1138 2642 1142
rect 2654 1138 2658 1142
rect 2670 1138 2674 1142
rect 3398 1147 3402 1151
rect 3438 1148 3442 1152
rect 3462 1148 3466 1152
rect 3526 1158 3530 1162
rect 3598 1158 3602 1162
rect 3750 1158 3754 1162
rect 4006 1158 4010 1162
rect 4030 1158 4034 1162
rect 4046 1158 4050 1162
rect 4166 1158 4170 1162
rect 4222 1158 4226 1162
rect 4262 1158 4266 1162
rect 4374 1158 4378 1162
rect 5110 1158 5114 1162
rect 5150 1158 5154 1162
rect 5190 1158 5194 1162
rect 3550 1148 3554 1152
rect 3694 1147 3698 1151
rect 3774 1148 3778 1152
rect 3862 1147 3866 1151
rect 3950 1148 3954 1152
rect 3982 1148 3986 1152
rect 4054 1148 4058 1152
rect 4102 1148 4106 1152
rect 4110 1148 4114 1152
rect 4134 1148 4138 1152
rect 4214 1148 4218 1152
rect 4230 1148 4234 1152
rect 4342 1148 4346 1152
rect 4438 1148 4442 1152
rect 4678 1148 4682 1152
rect 4742 1147 4746 1151
rect 4886 1148 4890 1152
rect 4902 1148 4906 1152
rect 4990 1148 4994 1152
rect 5078 1148 5082 1152
rect 5102 1148 5106 1152
rect 5118 1148 5122 1152
rect 5166 1148 5170 1152
rect 5190 1148 5194 1152
rect 5206 1148 5210 1152
rect 5238 1148 5242 1152
rect 5302 1148 5306 1152
rect 2718 1138 2722 1142
rect 2758 1138 2762 1142
rect 2774 1138 2778 1142
rect 2838 1138 2842 1142
rect 2846 1138 2850 1142
rect 2894 1138 2898 1142
rect 2934 1138 2938 1142
rect 2966 1138 2970 1142
rect 2974 1138 2978 1142
rect 2990 1138 2994 1142
rect 3046 1138 3050 1142
rect 3086 1138 3090 1142
rect 3390 1138 3394 1142
rect 3470 1138 3474 1142
rect 3478 1138 3482 1142
rect 3542 1138 3546 1142
rect 3558 1138 3562 1142
rect 3582 1138 3586 1142
rect 3606 1138 3610 1142
rect 3710 1138 3714 1142
rect 3726 1138 3730 1142
rect 3774 1138 3778 1142
rect 3830 1138 3834 1142
rect 3846 1138 3850 1142
rect 3870 1138 3874 1142
rect 3958 1138 3962 1142
rect 3990 1138 3994 1142
rect 3998 1138 4002 1142
rect 4030 1138 4034 1142
rect 4046 1138 4050 1142
rect 4134 1138 4138 1142
rect 4182 1138 4186 1142
rect 4206 1138 4210 1142
rect 4230 1138 4234 1142
rect 4294 1138 4298 1142
rect 4446 1138 4450 1142
rect 4558 1138 4562 1142
rect 4566 1138 4570 1142
rect 4614 1138 4618 1142
rect 4814 1138 4818 1142
rect 4942 1138 4946 1142
rect 4982 1138 4986 1142
rect 5030 1138 5034 1142
rect 5078 1138 5082 1142
rect 5126 1138 5130 1142
rect 5214 1138 5218 1142
rect 5262 1138 5266 1142
rect 6 1128 10 1132
rect 86 1128 90 1132
rect 174 1128 178 1132
rect 190 1128 194 1132
rect 262 1128 266 1132
rect 326 1128 330 1132
rect 414 1128 418 1132
rect 430 1128 434 1132
rect 574 1128 578 1132
rect 582 1128 586 1132
rect 694 1128 698 1132
rect 750 1128 754 1132
rect 758 1128 762 1132
rect 1062 1128 1066 1132
rect 1070 1128 1074 1132
rect 1118 1128 1122 1132
rect 1238 1128 1242 1132
rect 1390 1128 1394 1132
rect 1574 1128 1578 1132
rect 1662 1128 1666 1132
rect 1790 1128 1794 1132
rect 1886 1128 1890 1132
rect 1958 1128 1962 1132
rect 2158 1128 2162 1132
rect 2190 1128 2194 1132
rect 2622 1128 2626 1132
rect 2638 1128 2642 1132
rect 2758 1128 2762 1132
rect 2918 1128 2922 1132
rect 2998 1128 3002 1132
rect 3502 1128 3506 1132
rect 3574 1128 3578 1132
rect 3606 1128 3610 1132
rect 3622 1128 3626 1132
rect 3726 1128 3730 1132
rect 3798 1128 3802 1132
rect 3830 1128 3834 1132
rect 3974 1128 3978 1132
rect 4190 1128 4194 1132
rect 4262 1128 4266 1132
rect 4278 1128 4282 1132
rect 4310 1128 4314 1132
rect 4326 1128 4330 1132
rect 4742 1128 4746 1132
rect 4902 1128 4906 1132
rect 4910 1128 4914 1132
rect 4974 1128 4978 1132
rect 5142 1128 5146 1132
rect 5182 1128 5186 1132
rect 5230 1127 5234 1131
rect 5270 1128 5274 1132
rect 22 1118 26 1122
rect 270 1118 274 1122
rect 374 1118 378 1122
rect 550 1118 554 1122
rect 630 1118 634 1122
rect 662 1118 666 1122
rect 870 1118 874 1122
rect 918 1118 922 1122
rect 926 1118 930 1122
rect 966 1118 970 1122
rect 1102 1118 1106 1122
rect 1110 1118 1114 1122
rect 1126 1118 1130 1122
rect 1142 1118 1146 1122
rect 1174 1118 1178 1122
rect 1182 1118 1186 1122
rect 1366 1118 1370 1122
rect 1494 1118 1498 1122
rect 1534 1118 1538 1122
rect 1606 1118 1610 1122
rect 1654 1118 1658 1122
rect 1686 1118 1690 1122
rect 1694 1118 1698 1122
rect 1734 1118 1738 1122
rect 2198 1118 2202 1122
rect 2214 1118 2218 1122
rect 2246 1118 2250 1122
rect 2254 1118 2258 1122
rect 2334 1118 2338 1122
rect 2870 1118 2874 1122
rect 3214 1118 3218 1122
rect 3310 1118 3314 1122
rect 3494 1118 3498 1122
rect 3566 1118 3570 1122
rect 3782 1118 3786 1122
rect 3966 1118 3970 1122
rect 4070 1118 4074 1122
rect 4126 1118 4130 1122
rect 4382 1118 4386 1122
rect 4598 1118 4602 1122
rect 4622 1118 4626 1122
rect 5070 1118 5074 1122
rect 5302 1118 5306 1122
rect 6 1108 10 1112
rect 774 1108 778 1112
rect 1118 1108 1122 1112
rect 1574 1108 1578 1112
rect 2190 1108 2194 1112
rect 3766 1108 3770 1112
rect 5182 1108 5186 1112
rect 5270 1108 5274 1112
rect 858 1103 862 1107
rect 865 1103 869 1107
rect 1874 1103 1878 1107
rect 1881 1103 1885 1107
rect 2906 1103 2910 1107
rect 2913 1103 2917 1107
rect 3930 1103 3934 1107
rect 3937 1103 3941 1107
rect 4954 1103 4958 1107
rect 4961 1103 4965 1107
rect 646 1098 650 1102
rect 718 1098 722 1102
rect 934 1098 938 1102
rect 1518 1098 1522 1102
rect 1598 1098 1602 1102
rect 2302 1098 2306 1102
rect 2822 1098 2826 1102
rect 2846 1098 2850 1102
rect 4918 1098 4922 1102
rect 4990 1098 4994 1102
rect 86 1088 90 1092
rect 182 1088 186 1092
rect 462 1088 466 1092
rect 518 1088 522 1092
rect 654 1088 658 1092
rect 662 1088 666 1092
rect 830 1088 834 1092
rect 846 1088 850 1092
rect 886 1088 890 1092
rect 910 1088 914 1092
rect 1286 1088 1290 1092
rect 1390 1088 1394 1092
rect 1662 1088 1666 1092
rect 1782 1088 1786 1092
rect 1814 1088 1818 1092
rect 1902 1088 1906 1092
rect 2070 1088 2074 1092
rect 2110 1088 2114 1092
rect 2326 1088 2330 1092
rect 2382 1088 2386 1092
rect 2454 1088 2458 1092
rect 2566 1088 2570 1092
rect 2590 1088 2594 1092
rect 2614 1088 2618 1092
rect 2638 1088 2642 1092
rect 2678 1088 2682 1092
rect 2718 1088 2722 1092
rect 2862 1088 2866 1092
rect 2966 1088 2970 1092
rect 3358 1088 3362 1092
rect 3366 1088 3370 1092
rect 3486 1088 3490 1092
rect 3502 1088 3506 1092
rect 3614 1088 3618 1092
rect 3878 1088 3882 1092
rect 4014 1088 4018 1092
rect 4214 1088 4218 1092
rect 4246 1088 4250 1092
rect 4438 1088 4442 1092
rect 4638 1088 4642 1092
rect 4694 1088 4698 1092
rect 4838 1088 4842 1092
rect 4870 1088 4874 1092
rect 4886 1088 4890 1092
rect 4894 1088 4898 1092
rect 4950 1088 4954 1092
rect 4982 1088 4986 1092
rect 5142 1088 5146 1092
rect 5158 1088 5162 1092
rect 5166 1088 5170 1092
rect 5222 1088 5226 1092
rect 14 1079 18 1083
rect 30 1078 34 1082
rect 142 1078 146 1082
rect 166 1078 170 1082
rect 390 1078 394 1082
rect 526 1078 530 1082
rect 646 1078 650 1082
rect 710 1078 714 1082
rect 718 1078 722 1082
rect 934 1078 938 1082
rect 990 1078 994 1082
rect 1070 1078 1074 1082
rect 1126 1078 1130 1082
rect 1134 1078 1138 1082
rect 1198 1078 1202 1082
rect 1238 1078 1242 1082
rect 1278 1078 1282 1082
rect 1326 1078 1330 1082
rect 1550 1078 1554 1082
rect 1598 1078 1602 1082
rect 1622 1078 1626 1082
rect 1630 1078 1634 1082
rect 1878 1078 1882 1082
rect 1942 1078 1946 1082
rect 1974 1078 1978 1082
rect 2134 1078 2138 1082
rect 2190 1078 2194 1082
rect 2302 1078 2306 1082
rect 2350 1078 2354 1082
rect 2542 1078 2546 1082
rect 2574 1078 2578 1082
rect 2606 1078 2610 1082
rect 2742 1078 2746 1082
rect 2894 1078 2898 1082
rect 3070 1079 3074 1083
rect 3494 1078 3498 1082
rect 3622 1078 3626 1082
rect 3686 1078 3690 1082
rect 3742 1078 3746 1082
rect 4022 1078 4026 1082
rect 4094 1078 4098 1082
rect 4238 1078 4242 1082
rect 4310 1078 4314 1082
rect 4366 1078 4370 1082
rect 4462 1079 4466 1083
rect 4478 1078 4482 1082
rect 4494 1078 4498 1082
rect 4502 1078 4506 1082
rect 4526 1078 4530 1082
rect 4542 1078 4546 1082
rect 4550 1078 4554 1082
rect 4742 1078 4746 1082
rect 4918 1078 4922 1082
rect 4990 1078 4994 1082
rect 5174 1078 5178 1082
rect 5198 1078 5202 1082
rect 5278 1079 5282 1083
rect 126 1068 130 1072
rect 150 1068 154 1072
rect 214 1068 218 1072
rect 222 1068 226 1072
rect 270 1068 274 1072
rect 366 1068 370 1072
rect 6 1058 10 1062
rect 38 1058 42 1062
rect 62 1058 66 1062
rect 118 1058 122 1062
rect 150 1058 154 1062
rect 278 1058 282 1062
rect 302 1058 306 1062
rect 374 1058 378 1062
rect 406 1068 410 1072
rect 470 1068 474 1072
rect 510 1068 514 1072
rect 582 1068 586 1072
rect 622 1068 626 1072
rect 638 1068 642 1072
rect 662 1068 666 1072
rect 702 1068 706 1072
rect 734 1068 738 1072
rect 774 1068 778 1072
rect 822 1068 826 1072
rect 854 1068 858 1072
rect 878 1068 882 1072
rect 934 1068 938 1072
rect 942 1068 946 1072
rect 1110 1068 1114 1072
rect 1118 1068 1122 1072
rect 1142 1068 1146 1072
rect 1182 1068 1186 1072
rect 1262 1068 1266 1072
rect 1334 1068 1338 1072
rect 1398 1068 1402 1072
rect 1438 1068 1442 1072
rect 1526 1068 1530 1072
rect 1550 1068 1554 1072
rect 1566 1068 1570 1072
rect 1742 1068 1746 1072
rect 1758 1068 1762 1072
rect 1806 1068 1810 1072
rect 1838 1068 1842 1072
rect 1846 1068 1850 1072
rect 1926 1068 1930 1072
rect 2078 1068 2082 1072
rect 2126 1068 2130 1072
rect 2142 1068 2146 1072
rect 2174 1068 2178 1072
rect 2198 1068 2202 1072
rect 2294 1068 2298 1072
rect 2310 1068 2314 1072
rect 2366 1068 2370 1072
rect 414 1058 418 1062
rect 446 1058 450 1062
rect 478 1058 482 1062
rect 502 1058 506 1062
rect 542 1058 546 1062
rect 566 1058 570 1062
rect 606 1058 610 1062
rect 638 1058 642 1062
rect 678 1058 682 1062
rect 734 1058 738 1062
rect 758 1058 762 1062
rect 846 1058 850 1062
rect 966 1058 970 1062
rect 1014 1058 1018 1062
rect 1046 1058 1050 1062
rect 1094 1058 1098 1062
rect 1102 1058 1106 1062
rect 1150 1058 1154 1062
rect 1206 1058 1210 1062
rect 1222 1058 1226 1062
rect 1270 1058 1274 1062
rect 1302 1058 1306 1062
rect 1310 1058 1314 1062
rect 1326 1058 1330 1062
rect 1342 1058 1346 1062
rect 1422 1058 1426 1062
rect 1446 1058 1450 1062
rect 1478 1058 1482 1062
rect 1510 1058 1514 1062
rect 1550 1058 1554 1062
rect 1558 1058 1562 1062
rect 1590 1058 1594 1062
rect 1614 1058 1618 1062
rect 1654 1058 1658 1062
rect 1726 1059 1730 1063
rect 1830 1058 1834 1062
rect 1966 1058 1970 1062
rect 2014 1058 2018 1062
rect 2038 1058 2042 1062
rect 2206 1058 2210 1062
rect 2238 1058 2242 1062
rect 2254 1058 2258 1062
rect 2350 1058 2354 1062
rect 2438 1068 2442 1072
rect 2486 1068 2490 1072
rect 2598 1068 2602 1072
rect 2694 1066 2698 1070
rect 2702 1068 2706 1072
rect 2726 1068 2730 1072
rect 2854 1068 2858 1072
rect 2886 1068 2890 1072
rect 2950 1066 2954 1070
rect 2958 1068 2962 1072
rect 3046 1068 3050 1072
rect 3086 1068 3090 1072
rect 3150 1068 3154 1072
rect 3158 1068 3162 1072
rect 3206 1068 3210 1072
rect 3230 1068 3234 1072
rect 3294 1068 3298 1072
rect 3334 1068 3338 1072
rect 3446 1068 3450 1072
rect 3582 1068 3586 1072
rect 3606 1068 3610 1072
rect 3662 1068 3666 1072
rect 3694 1068 3698 1072
rect 3910 1068 3914 1072
rect 3982 1068 3986 1072
rect 4006 1068 4010 1072
rect 4238 1068 4242 1072
rect 4342 1068 4346 1072
rect 4358 1068 4362 1072
rect 4406 1068 4410 1072
rect 4414 1068 4418 1072
rect 4494 1068 4498 1072
rect 4526 1068 4530 1072
rect 4598 1068 4602 1072
rect 4606 1068 4610 1072
rect 4654 1068 4658 1072
rect 4662 1068 4666 1072
rect 4710 1068 4714 1072
rect 4862 1068 4866 1072
rect 4870 1068 4874 1072
rect 4918 1068 4922 1072
rect 4926 1068 4930 1072
rect 4990 1068 4994 1072
rect 5046 1068 5050 1072
rect 5166 1068 5170 1072
rect 5190 1068 5194 1072
rect 5262 1068 5266 1072
rect 2478 1058 2482 1062
rect 2510 1058 2514 1062
rect 2526 1058 2530 1062
rect 2550 1058 2554 1062
rect 2622 1058 2626 1062
rect 2662 1058 2666 1062
rect 2742 1058 2746 1062
rect 2782 1058 2786 1062
rect 2814 1058 2818 1062
rect 2830 1058 2834 1062
rect 2846 1058 2850 1062
rect 2878 1058 2882 1062
rect 2910 1058 2914 1062
rect 2926 1058 2930 1062
rect 3022 1058 3026 1062
rect 3062 1058 3066 1062
rect 3166 1058 3170 1062
rect 3198 1058 3202 1062
rect 3262 1059 3266 1063
rect 3342 1058 3346 1062
rect 3430 1059 3434 1063
rect 3478 1058 3482 1062
rect 3558 1058 3562 1062
rect 3622 1058 3626 1062
rect 3702 1058 3706 1062
rect 3734 1058 3738 1062
rect 3758 1058 3762 1062
rect 3766 1058 3770 1062
rect 3822 1058 3826 1062
rect 3846 1058 3850 1062
rect 3966 1058 3970 1062
rect 4086 1058 4090 1062
rect 4150 1059 4154 1063
rect 4222 1058 4226 1062
rect 4294 1058 4298 1062
rect 4382 1058 4386 1062
rect 4398 1058 4402 1062
rect 4454 1058 4458 1062
rect 4518 1058 4522 1062
rect 4598 1058 4602 1062
rect 4742 1059 4746 1063
rect 4774 1058 4778 1062
rect 4934 1058 4938 1062
rect 4974 1058 4978 1062
rect 4998 1058 5002 1062
rect 5078 1059 5082 1063
rect 5110 1058 5114 1062
rect 5198 1058 5202 1062
rect 5254 1058 5258 1062
rect 5286 1058 5290 1062
rect 70 1048 74 1052
rect 78 1048 82 1052
rect 102 1048 106 1052
rect 174 1048 178 1052
rect 198 1048 202 1052
rect 430 1048 434 1052
rect 494 1048 498 1052
rect 534 1048 538 1052
rect 566 1048 570 1052
rect 582 1048 586 1052
rect 622 1048 626 1052
rect 694 1048 698 1052
rect 726 1048 730 1052
rect 742 1048 746 1052
rect 830 1048 834 1052
rect 1022 1048 1026 1052
rect 1094 1048 1098 1052
rect 1166 1048 1170 1052
rect 1214 1048 1218 1052
rect 1358 1048 1362 1052
rect 1430 1048 1434 1052
rect 1462 1048 1466 1052
rect 1470 1048 1474 1052
rect 1502 1048 1506 1052
rect 1846 1048 1850 1052
rect 1902 1048 1906 1052
rect 1942 1048 1946 1052
rect 2166 1048 2170 1052
rect 2326 1048 2330 1052
rect 2358 1048 2362 1052
rect 2462 1048 2466 1052
rect 2494 1048 2498 1052
rect 2582 1048 2586 1052
rect 2670 1048 2674 1052
rect 2710 1048 2714 1052
rect 2734 1048 2738 1052
rect 2766 1048 2770 1052
rect 2790 1048 2794 1052
rect 2798 1048 2802 1052
rect 2830 1048 2834 1052
rect 2862 1048 2866 1052
rect 3182 1048 3186 1052
rect 3902 1048 3906 1052
rect 3934 1048 3938 1052
rect 4358 1048 4362 1052
rect 4382 1048 4386 1052
rect 4430 1048 4434 1052
rect 4574 1048 4578 1052
rect 4886 1048 4890 1052
rect 5150 1048 5154 1052
rect 54 1038 58 1042
rect 238 1038 242 1042
rect 550 1038 554 1042
rect 958 1038 962 1042
rect 1006 1038 1010 1042
rect 1014 1038 1018 1042
rect 1038 1038 1042 1042
rect 1414 1038 1418 1042
rect 1470 1038 1474 1042
rect 1486 1038 1490 1042
rect 2262 1038 2266 1042
rect 2278 1038 2282 1042
rect 2342 1038 2346 1042
rect 2654 1038 2658 1042
rect 2750 1038 2754 1042
rect 2774 1038 2778 1042
rect 2806 1038 2810 1042
rect 3222 1038 3226 1042
rect 4030 1038 4034 1042
rect 4398 1038 4402 1042
rect 62 1028 66 1032
rect 542 1028 546 1032
rect 1046 1028 1050 1032
rect 2662 1028 2666 1032
rect 478 1018 482 1022
rect 678 1018 682 1022
rect 790 1018 794 1022
rect 990 1018 994 1022
rect 1230 1018 1234 1022
rect 1246 1018 1250 1022
rect 1446 1018 1450 1022
rect 2230 1018 2234 1022
rect 2270 1018 2274 1022
rect 2510 1018 2514 1022
rect 3326 1018 3330 1022
rect 3670 1018 3674 1022
rect 3726 1018 3730 1022
rect 3990 1018 3994 1022
rect 5222 1018 5226 1022
rect 346 1003 350 1007
rect 353 1003 357 1007
rect 1370 1003 1374 1007
rect 1377 1003 1381 1007
rect 2394 1003 2398 1007
rect 2401 1003 2405 1007
rect 3418 1003 3422 1007
rect 3425 1003 3429 1007
rect 4442 1003 4446 1007
rect 4449 1003 4453 1007
rect 150 988 154 992
rect 286 988 290 992
rect 382 988 386 992
rect 438 988 442 992
rect 1494 988 1498 992
rect 1534 988 1538 992
rect 1590 988 1594 992
rect 1710 988 1714 992
rect 2102 988 2106 992
rect 2358 988 2362 992
rect 2374 988 2378 992
rect 2742 988 2746 992
rect 2854 988 2858 992
rect 2862 988 2866 992
rect 3142 988 3146 992
rect 3310 988 3314 992
rect 3478 988 3482 992
rect 3574 988 3578 992
rect 3646 988 3650 992
rect 3854 988 3858 992
rect 3886 988 3890 992
rect 3982 988 3986 992
rect 4182 988 4186 992
rect 4286 988 4290 992
rect 4318 988 4322 992
rect 4334 988 4338 992
rect 4422 988 4426 992
rect 4526 988 4530 992
rect 4566 988 4570 992
rect 4582 988 4586 992
rect 4670 988 4674 992
rect 4830 988 4834 992
rect 4854 988 4858 992
rect 4910 988 4914 992
rect 5022 988 5026 992
rect 846 978 850 982
rect 974 978 978 982
rect 3118 978 3122 982
rect 3694 978 3698 982
rect 238 968 242 972
rect 366 968 370 972
rect 462 968 466 972
rect 502 968 506 972
rect 526 968 530 972
rect 614 968 618 972
rect 630 968 634 972
rect 654 968 658 972
rect 942 968 946 972
rect 966 968 970 972
rect 990 968 994 972
rect 1030 968 1034 972
rect 1206 968 1210 972
rect 1310 968 1314 972
rect 1430 968 1434 972
rect 1542 968 1546 972
rect 1718 968 1722 972
rect 1758 968 1762 972
rect 2350 968 2354 972
rect 2382 968 2386 972
rect 2878 968 2882 972
rect 3374 968 3378 972
rect 3486 968 3490 972
rect 3638 968 3642 972
rect 3670 968 3674 972
rect 3862 968 3866 972
rect 3990 968 3994 972
rect 4310 968 4314 972
rect 4534 968 4538 972
rect 4598 968 4602 972
rect 4750 968 4754 972
rect 4862 968 4866 972
rect 5102 968 5106 972
rect 134 958 138 962
rect 22 948 26 952
rect 46 948 50 952
rect 70 948 74 952
rect 78 948 82 952
rect 174 958 178 962
rect 214 958 218 962
rect 390 958 394 962
rect 422 958 426 962
rect 478 958 482 962
rect 542 958 546 962
rect 582 958 586 962
rect 638 958 642 962
rect 670 958 674 962
rect 678 958 682 962
rect 830 958 834 962
rect 982 958 986 962
rect 990 958 994 962
rect 1014 958 1018 962
rect 1046 958 1050 962
rect 1094 958 1098 962
rect 1230 958 1234 962
rect 1302 958 1306 962
rect 1446 958 1450 962
rect 1454 958 1458 962
rect 1526 958 1530 962
rect 1694 958 1698 962
rect 1702 958 1706 962
rect 1750 958 1754 962
rect 1846 958 1850 962
rect 2118 958 2122 962
rect 2366 958 2370 962
rect 2414 958 2418 962
rect 2438 958 2442 962
rect 2526 958 2530 962
rect 2558 958 2562 962
rect 2990 958 2994 962
rect 166 948 170 952
rect 198 948 202 952
rect 222 948 226 952
rect 278 948 282 952
rect 366 948 370 952
rect 406 948 410 952
rect 438 948 442 952
rect 470 948 474 952
rect 534 948 538 952
rect 574 948 578 952
rect 662 948 666 952
rect 678 948 682 952
rect 710 948 714 952
rect 726 948 730 952
rect 766 948 770 952
rect 158 938 162 942
rect 190 938 194 942
rect 222 938 226 942
rect 270 938 274 942
rect 414 938 418 942
rect 446 938 450 942
rect 494 938 498 942
rect 566 938 570 942
rect 622 938 626 942
rect 638 938 642 942
rect 798 947 802 951
rect 886 948 890 952
rect 902 948 906 952
rect 942 948 946 952
rect 974 948 978 952
rect 998 948 1002 952
rect 1038 948 1042 952
rect 1054 948 1058 952
rect 1110 948 1114 952
rect 1246 948 1250 952
rect 710 938 714 942
rect 854 938 858 942
rect 1374 947 1378 951
rect 1414 948 1418 952
rect 1438 948 1442 952
rect 1494 948 1498 952
rect 1550 948 1554 952
rect 1566 948 1570 952
rect 1622 948 1626 952
rect 1630 948 1634 952
rect 1694 948 1698 952
rect 1710 948 1714 952
rect 1782 948 1786 952
rect 1934 948 1938 952
rect 934 938 938 942
rect 1078 938 1082 942
rect 1094 938 1098 942
rect 1134 938 1138 942
rect 1174 938 1178 942
rect 1222 938 1226 942
rect 1246 938 1250 942
rect 1262 938 1266 942
rect 1286 938 1290 942
rect 1390 938 1394 942
rect 1470 938 1474 942
rect 1510 938 1514 942
rect 1582 938 1586 942
rect 1670 938 1674 942
rect 1734 938 1738 942
rect 1758 938 1762 942
rect 1774 938 1778 942
rect 1790 938 1794 942
rect 1838 938 1842 942
rect 1862 938 1866 942
rect 1886 938 1890 942
rect 2022 947 2026 951
rect 2054 948 2058 952
rect 2102 948 2106 952
rect 2118 948 2122 952
rect 2142 948 2146 952
rect 2190 948 2194 952
rect 2214 948 2218 952
rect 2270 948 2274 952
rect 2358 948 2362 952
rect 2390 948 2394 952
rect 2430 948 2434 952
rect 2494 948 2498 952
rect 2534 948 2538 952
rect 2598 948 2602 952
rect 2646 948 2650 952
rect 14 927 18 931
rect 38 927 42 931
rect 62 927 66 931
rect 110 928 114 932
rect 278 928 282 932
rect 302 928 306 932
rect 334 928 338 932
rect 390 928 394 932
rect 502 928 506 932
rect 550 928 554 932
rect 726 928 730 932
rect 918 928 922 932
rect 1038 928 1042 932
rect 1134 928 1138 932
rect 1150 928 1154 932
rect 1166 928 1170 932
rect 1278 928 1282 932
rect 1478 928 1482 932
rect 1566 928 1570 932
rect 1614 928 1618 932
rect 1662 928 1666 932
rect 2054 938 2058 942
rect 2094 938 2098 942
rect 2134 938 2138 942
rect 2334 938 2338 942
rect 2678 947 2682 951
rect 2798 948 2802 952
rect 2822 948 2826 952
rect 2958 947 2962 951
rect 3054 947 3058 951
rect 3102 948 3106 952
rect 3126 948 3130 952
rect 3150 948 3154 952
rect 3182 958 3186 962
rect 3350 958 3354 962
rect 3430 958 3434 962
rect 3502 958 3506 962
rect 3542 958 3546 962
rect 3198 948 3202 952
rect 3222 948 3226 952
rect 3246 948 3250 952
rect 3374 948 3378 952
rect 3390 948 3394 952
rect 3470 948 3474 952
rect 3494 948 3498 952
rect 3534 948 3538 952
rect 3542 948 3546 952
rect 3614 958 3618 962
rect 3622 958 3626 962
rect 3758 958 3762 962
rect 3838 958 3842 962
rect 3846 958 3850 962
rect 3934 958 3938 962
rect 3974 958 3978 962
rect 4022 958 4026 962
rect 4438 958 4442 962
rect 4494 958 4498 962
rect 4558 958 4562 962
rect 4574 958 4578 962
rect 4614 958 4618 962
rect 4654 958 4658 962
rect 4734 958 4738 962
rect 4790 958 4794 962
rect 4878 958 4882 962
rect 4950 958 4954 962
rect 5046 958 5050 962
rect 5262 958 5266 962
rect 3590 948 3594 952
rect 3630 948 3634 952
rect 3678 948 3682 952
rect 3726 948 3730 952
rect 3782 948 3786 952
rect 3790 948 3794 952
rect 3806 948 3810 952
rect 3854 948 3858 952
rect 3902 948 3906 952
rect 3966 948 3970 952
rect 3982 948 3986 952
rect 4046 948 4050 952
rect 4118 948 4122 952
rect 4150 948 4154 952
rect 4174 948 4178 952
rect 4222 948 4226 952
rect 4302 948 4306 952
rect 4342 948 4346 952
rect 4374 948 4378 952
rect 4462 948 4466 952
rect 4478 948 4482 952
rect 4494 948 4498 952
rect 4510 948 4514 952
rect 4542 948 4546 952
rect 4646 948 4650 952
rect 4670 948 4674 952
rect 4686 948 4690 952
rect 4726 948 4730 952
rect 4774 948 4778 952
rect 4870 948 4874 952
rect 4990 948 4994 952
rect 5174 948 5178 952
rect 5198 948 5202 952
rect 5238 948 5242 952
rect 5286 948 5290 952
rect 2462 938 2466 942
rect 2486 938 2490 942
rect 2526 938 2530 942
rect 2574 938 2578 942
rect 2606 938 2610 942
rect 2710 938 2714 942
rect 2758 938 2762 942
rect 2774 938 2778 942
rect 2974 938 2978 942
rect 3046 938 3050 942
rect 3086 938 3090 942
rect 3158 938 3162 942
rect 3206 938 3210 942
rect 3254 938 3258 942
rect 3294 938 3298 942
rect 3334 938 3338 942
rect 3414 938 3418 942
rect 3534 938 3538 942
rect 3598 938 3602 942
rect 3614 938 3618 942
rect 3718 938 3722 942
rect 3814 938 3818 942
rect 3822 938 3826 942
rect 3894 938 3898 942
rect 3958 938 3962 942
rect 4006 938 4010 942
rect 4030 938 4034 942
rect 4062 938 4066 942
rect 4086 938 4090 942
rect 4126 938 4130 942
rect 4142 938 4146 942
rect 4174 938 4178 942
rect 4214 938 4218 942
rect 4270 938 4274 942
rect 4374 938 4378 942
rect 4382 938 4386 942
rect 4486 938 4490 942
rect 4518 938 4522 942
rect 4558 938 4562 942
rect 4598 938 4602 942
rect 4614 938 4618 942
rect 4638 938 4642 942
rect 4678 938 4682 942
rect 4694 938 4698 942
rect 4766 938 4770 942
rect 4846 938 4850 942
rect 4886 938 4890 942
rect 4934 938 4938 942
rect 4974 938 4978 942
rect 5038 938 5042 942
rect 5062 938 5066 942
rect 5070 938 5074 942
rect 5126 938 5130 942
rect 2022 928 2026 932
rect 2070 928 2074 932
rect 2078 928 2082 932
rect 2150 928 2154 932
rect 2214 928 2218 932
rect 2262 928 2266 932
rect 2430 928 2434 932
rect 2478 928 2482 932
rect 2494 928 2498 932
rect 2550 928 2554 932
rect 2870 928 2874 932
rect 3086 928 3090 932
rect 3110 928 3114 932
rect 3134 928 3138 932
rect 3222 928 3226 932
rect 3270 928 3274 932
rect 3294 928 3298 932
rect 3326 928 3330 932
rect 3422 928 3426 932
rect 3510 928 3514 932
rect 3654 928 3658 932
rect 3710 928 3714 932
rect 3878 928 3882 932
rect 4054 928 4058 932
rect 4134 928 4138 932
rect 4174 928 4178 932
rect 4198 928 4202 932
rect 4206 928 4210 932
rect 4262 928 4266 932
rect 4326 928 4330 932
rect 4366 928 4370 932
rect 4398 928 4402 932
rect 5262 938 5266 942
rect 5278 938 5282 942
rect 4438 928 4442 932
rect 4702 928 4706 932
rect 4710 928 4714 932
rect 4726 928 4730 932
rect 4958 928 4962 932
rect 534 918 538 922
rect 558 918 562 922
rect 710 918 714 922
rect 734 918 738 922
rect 1094 918 1098 922
rect 1238 918 1242 922
rect 1270 918 1274 922
rect 1302 918 1306 922
rect 1454 918 1458 922
rect 1638 918 1642 922
rect 1822 918 1826 922
rect 1918 918 1922 922
rect 2422 918 2426 922
rect 2558 918 2562 922
rect 2574 918 2578 922
rect 2582 918 2586 922
rect 2614 918 2618 922
rect 2622 918 2626 922
rect 2854 918 2858 922
rect 3174 918 3178 922
rect 3230 918 3234 922
rect 3462 918 3466 922
rect 3518 918 3522 922
rect 3838 918 3842 922
rect 3886 918 3890 922
rect 3950 918 3954 922
rect 4126 918 4130 922
rect 4246 918 4250 922
rect 1662 908 1666 912
rect 1734 908 1738 912
rect 2238 908 2242 912
rect 2550 908 2554 912
rect 5150 908 5154 912
rect 858 903 862 907
rect 865 903 869 907
rect 1874 903 1878 907
rect 1881 903 1885 907
rect 2906 903 2910 907
rect 2913 903 2917 907
rect 3930 903 3934 907
rect 3937 903 3941 907
rect 4954 903 4958 907
rect 4961 903 4965 907
rect 702 898 706 902
rect 2206 898 2210 902
rect 2502 898 2506 902
rect 3782 898 3786 902
rect 198 888 202 892
rect 390 888 394 892
rect 446 888 450 892
rect 510 888 514 892
rect 614 888 618 892
rect 686 888 690 892
rect 710 888 714 892
rect 726 888 730 892
rect 830 888 834 892
rect 838 888 842 892
rect 942 888 946 892
rect 1102 888 1106 892
rect 1150 888 1154 892
rect 1486 888 1490 892
rect 1534 888 1538 892
rect 1550 888 1554 892
rect 1590 888 1594 892
rect 1614 888 1618 892
rect 1686 888 1690 892
rect 1726 888 1730 892
rect 1886 888 1890 892
rect 1958 888 1962 892
rect 2054 888 2058 892
rect 2094 888 2098 892
rect 2134 888 2138 892
rect 2166 888 2170 892
rect 2230 888 2234 892
rect 2262 888 2266 892
rect 2302 888 2306 892
rect 2486 888 2490 892
rect 2646 888 2650 892
rect 2830 888 2834 892
rect 2966 888 2970 892
rect 2998 888 3002 892
rect 3022 888 3026 892
rect 3150 888 3154 892
rect 3350 888 3354 892
rect 3470 888 3474 892
rect 3518 888 3522 892
rect 3670 888 3674 892
rect 3726 888 3730 892
rect 3774 888 3778 892
rect 4110 888 4114 892
rect 4126 888 4130 892
rect 4222 888 4226 892
rect 4326 888 4330 892
rect 4366 888 4370 892
rect 4630 888 4634 892
rect 4670 888 4674 892
rect 4734 888 4738 892
rect 4742 888 4746 892
rect 4798 888 4802 892
rect 4822 888 4826 892
rect 4878 888 4882 892
rect 4974 888 4978 892
rect 5006 888 5010 892
rect 5110 888 5114 892
rect 5142 888 5146 892
rect 5190 888 5194 892
rect 5198 888 5202 892
rect 5270 888 5274 892
rect 5286 888 5290 892
rect 14 879 18 883
rect 38 879 42 883
rect 62 879 66 883
rect 454 878 458 882
rect 534 878 538 882
rect 550 878 554 882
rect 558 878 562 882
rect 646 878 650 882
rect 702 878 706 882
rect 886 878 890 882
rect 910 878 914 882
rect 990 878 994 882
rect 1134 878 1138 882
rect 1142 878 1146 882
rect 1174 878 1178 882
rect 1230 878 1234 882
rect 2006 878 2010 882
rect 2174 878 2178 882
rect 2206 878 2210 882
rect 2294 878 2298 882
rect 2494 878 2498 882
rect 2502 878 2506 882
rect 2550 878 2554 882
rect 2574 878 2578 882
rect 2582 878 2586 882
rect 2974 878 2978 882
rect 3006 878 3010 882
rect 3054 878 3058 882
rect 3078 878 3082 882
rect 3342 878 3346 882
rect 3406 878 3410 882
rect 3438 878 3442 882
rect 3462 878 3466 882
rect 3486 878 3490 882
rect 3510 878 3514 882
rect 3582 878 3586 882
rect 3622 878 3626 882
rect 3718 878 3722 882
rect 3742 878 3746 882
rect 4038 878 4042 882
rect 4046 878 4050 882
rect 4086 878 4090 882
rect 4118 878 4122 882
rect 4350 879 4354 883
rect 4486 878 4490 882
rect 4542 878 4546 882
rect 4678 878 4682 882
rect 4790 878 4794 882
rect 4814 878 4818 882
rect 4862 878 4866 882
rect 5030 878 5034 882
rect 5246 879 5250 883
rect 5262 878 5266 882
rect 278 868 282 872
rect 294 868 298 872
rect 358 868 362 872
rect 366 868 370 872
rect 382 868 386 872
rect 446 868 450 872
rect 486 868 490 872
rect 502 868 506 872
rect 534 868 538 872
rect 550 868 554 872
rect 606 868 610 872
rect 686 868 690 872
rect 734 868 738 872
rect 766 868 770 872
rect 862 868 866 872
rect 918 868 922 872
rect 966 868 970 872
rect 974 868 978 872
rect 990 868 994 872
rect 1062 868 1066 872
rect 1078 868 1082 872
rect 1086 868 1090 872
rect 1102 868 1106 872
rect 1158 868 1162 872
rect 1166 868 1170 872
rect 1198 868 1202 872
rect 1206 868 1210 872
rect 22 858 26 862
rect 46 858 50 862
rect 70 858 74 862
rect 126 859 130 863
rect 158 858 162 862
rect 262 859 266 863
rect 438 858 442 862
rect 494 858 498 862
rect 582 858 586 862
rect 654 858 658 862
rect 686 858 690 862
rect 726 858 730 862
rect 774 858 778 862
rect 854 858 858 862
rect 886 858 890 862
rect 942 858 946 862
rect 1006 858 1010 862
rect 1046 858 1050 862
rect 1110 858 1114 862
rect 1166 858 1170 862
rect 1214 858 1218 862
rect 1254 858 1258 862
rect 1270 868 1274 872
rect 1278 868 1282 872
rect 1318 868 1322 872
rect 1350 868 1354 872
rect 1414 868 1418 872
rect 1422 868 1426 872
rect 1454 868 1458 872
rect 1502 868 1506 872
rect 1534 868 1538 872
rect 1550 868 1554 872
rect 1606 868 1610 872
rect 1638 868 1642 872
rect 1646 868 1650 872
rect 1694 868 1698 872
rect 1294 858 1298 862
rect 1326 858 1330 862
rect 1430 858 1434 862
rect 1454 858 1458 862
rect 1510 858 1514 862
rect 1630 858 1634 862
rect 1766 868 1770 872
rect 1902 868 1906 872
rect 1918 868 1922 872
rect 1974 868 1978 872
rect 1982 868 1986 872
rect 2014 868 2018 872
rect 2038 868 2042 872
rect 2054 868 2058 872
rect 2110 868 2114 872
rect 2158 868 2162 872
rect 2174 868 2178 872
rect 2214 868 2218 872
rect 2222 868 2226 872
rect 2230 868 2234 872
rect 2238 868 2242 872
rect 2270 868 2274 872
rect 2286 868 2290 872
rect 2310 868 2314 872
rect 2318 868 2322 872
rect 2358 868 2362 872
rect 2502 868 2506 872
rect 2542 868 2546 872
rect 2566 868 2570 872
rect 2590 868 2594 872
rect 2638 868 2642 872
rect 2726 868 2730 872
rect 2742 868 2746 872
rect 2790 868 2794 872
rect 2822 868 2826 872
rect 2910 868 2914 872
rect 2942 868 2946 872
rect 3030 868 3034 872
rect 3102 868 3106 872
rect 3118 868 3122 872
rect 3126 868 3130 872
rect 3134 868 3138 872
rect 3214 868 3218 872
rect 3286 868 3290 872
rect 3302 868 3306 872
rect 3334 868 3338 872
rect 3390 868 3394 872
rect 3422 868 3426 872
rect 3438 868 3442 872
rect 3478 868 3482 872
rect 3630 868 3634 872
rect 3694 868 3698 872
rect 3774 868 3778 872
rect 3846 868 3850 872
rect 3870 868 3874 872
rect 3878 868 3882 872
rect 4030 868 4034 872
rect 4046 868 4050 872
rect 4182 868 4186 872
rect 4334 868 4338 872
rect 1790 858 1794 862
rect 2038 858 2042 862
rect 2134 858 2138 862
rect 2150 858 2154 862
rect 2246 858 2250 862
rect 2366 858 2370 862
rect 2382 858 2386 862
rect 2414 858 2418 862
rect 2446 858 2450 862
rect 2470 858 2474 862
rect 2518 858 2522 862
rect 2526 858 2530 862
rect 2558 858 2562 862
rect 2710 859 2714 863
rect 2790 858 2794 862
rect 2814 858 2818 862
rect 2894 859 2898 863
rect 2950 858 2954 862
rect 2990 858 2994 862
rect 3038 858 3042 862
rect 3054 858 3058 862
rect 3094 858 3098 862
rect 3206 858 3210 862
rect 3262 858 3266 862
rect 3302 858 3306 862
rect 3326 858 3330 862
rect 3382 858 3386 862
rect 3454 858 3458 862
rect 3478 858 3482 862
rect 3566 858 3570 862
rect 3638 858 3642 862
rect 3670 858 3674 862
rect 3694 858 3698 862
rect 3782 858 3786 862
rect 3838 858 3842 862
rect 3854 858 3858 862
rect 3886 858 3890 862
rect 3910 858 3914 862
rect 3966 858 3970 862
rect 3990 859 3994 863
rect 4022 858 4026 862
rect 4070 858 4074 862
rect 4094 858 4098 862
rect 4174 858 4178 862
rect 4254 858 4258 862
rect 4278 858 4282 862
rect 4358 858 4362 862
rect 4414 868 4418 872
rect 4462 868 4466 872
rect 4478 868 4482 872
rect 4486 868 4490 872
rect 4526 868 4530 872
rect 4646 868 4650 872
rect 4662 868 4666 872
rect 4702 868 4706 872
rect 4710 868 4714 872
rect 4398 858 4402 862
rect 4422 858 4426 862
rect 4718 866 4722 870
rect 4750 868 4754 872
rect 4766 868 4770 872
rect 4782 868 4786 872
rect 4870 868 4874 872
rect 4894 868 4898 872
rect 4926 868 4930 872
rect 4990 868 4994 872
rect 5014 868 5018 872
rect 5054 868 5058 872
rect 5174 868 5178 872
rect 5182 868 5186 872
rect 5230 868 5234 872
rect 5278 868 5282 872
rect 4518 858 4522 862
rect 4534 858 4538 862
rect 4574 858 4578 862
rect 4614 858 4618 862
rect 4646 858 4650 862
rect 4758 858 4762 862
rect 4838 858 4842 862
rect 4846 858 4850 862
rect 4902 858 4906 862
rect 4934 858 4938 862
rect 5030 858 5034 862
rect 5254 858 5258 862
rect 5286 858 5290 862
rect 398 848 402 852
rect 470 848 474 852
rect 590 848 594 852
rect 614 848 618 852
rect 710 848 714 852
rect 942 848 946 852
rect 998 848 1002 852
rect 1062 848 1066 852
rect 1078 848 1082 852
rect 1102 848 1106 852
rect 1134 848 1138 852
rect 1230 848 1234 852
rect 1238 848 1242 852
rect 1286 848 1290 852
rect 1342 848 1346 852
rect 1382 848 1386 852
rect 1446 848 1450 852
rect 1550 848 1554 852
rect 1982 848 1986 852
rect 2054 848 2058 852
rect 2142 848 2146 852
rect 2214 848 2218 852
rect 2286 848 2290 852
rect 2326 848 2330 852
rect 2406 848 2410 852
rect 2438 848 2442 852
rect 3046 848 3050 852
rect 3078 848 3082 852
rect 3110 848 3114 852
rect 3150 848 3154 852
rect 3254 848 3258 852
rect 3366 848 3370 852
rect 3678 848 3682 852
rect 3854 848 3858 852
rect 4078 848 4082 852
rect 4318 848 4322 852
rect 4366 848 4370 852
rect 4390 848 4394 852
rect 4478 848 4482 852
rect 4622 848 4626 852
rect 4630 848 4634 852
rect 4686 848 4690 852
rect 4886 848 4890 852
rect 4902 848 4906 852
rect 4918 848 4922 852
rect 4950 848 4954 852
rect 4998 848 5002 852
rect 5014 848 5018 852
rect 686 838 690 842
rect 1014 838 1018 842
rect 1022 838 1026 842
rect 1038 838 1042 842
rect 1302 838 1306 842
rect 1830 838 1834 842
rect 2134 838 2138 842
rect 2422 838 2426 842
rect 2454 838 2458 842
rect 3062 838 3066 842
rect 3158 838 3162 842
rect 3270 838 3274 842
rect 3926 838 3930 842
rect 4062 838 4066 842
rect 4406 838 4410 842
rect 4582 838 4586 842
rect 4606 838 4610 842
rect 5038 838 5042 842
rect 1046 828 1050 832
rect 1326 828 1330 832
rect 2414 828 2418 832
rect 190 818 194 822
rect 1254 818 1258 822
rect 1310 818 1314 822
rect 2622 818 2626 822
rect 2774 818 2778 822
rect 3278 818 3282 822
rect 3702 818 3706 822
rect 3822 818 3826 822
rect 4558 818 4562 822
rect 4574 818 4578 822
rect 4598 818 4602 822
rect 5110 818 5114 822
rect 4030 808 4034 812
rect 4078 808 4082 812
rect 346 803 350 807
rect 353 803 357 807
rect 1370 803 1374 807
rect 1377 803 1381 807
rect 2394 803 2398 807
rect 2401 803 2405 807
rect 3418 803 3422 807
rect 3425 803 3429 807
rect 4442 803 4446 807
rect 4449 803 4453 807
rect 638 788 642 792
rect 1094 788 1098 792
rect 1142 788 1146 792
rect 1166 788 1170 792
rect 1430 788 1434 792
rect 1630 788 1634 792
rect 1742 788 1746 792
rect 1846 788 1850 792
rect 1870 788 1874 792
rect 2094 788 2098 792
rect 2166 788 2170 792
rect 2270 788 2274 792
rect 2286 788 2290 792
rect 2358 788 2362 792
rect 2798 788 2802 792
rect 3294 788 3298 792
rect 3614 788 3618 792
rect 3726 788 3730 792
rect 3966 788 3970 792
rect 4294 788 4298 792
rect 4366 788 4370 792
rect 4430 788 4434 792
rect 4566 788 4570 792
rect 4606 788 4610 792
rect 4694 788 4698 792
rect 4766 788 4770 792
rect 4814 788 4818 792
rect 4830 788 4834 792
rect 4982 788 4986 792
rect 5030 788 5034 792
rect 5126 788 5130 792
rect 5262 788 5266 792
rect 302 778 306 782
rect 1958 778 1962 782
rect 2494 778 2498 782
rect 4318 778 4322 782
rect 4670 778 4674 782
rect 342 768 346 772
rect 446 768 450 772
rect 470 768 474 772
rect 494 768 498 772
rect 694 768 698 772
rect 1118 768 1122 772
rect 1150 768 1154 772
rect 1174 768 1178 772
rect 1470 768 1474 772
rect 1510 768 1514 772
rect 1542 768 1546 772
rect 1790 768 1794 772
rect 2142 768 2146 772
rect 2294 768 2298 772
rect 3558 768 3562 772
rect 3694 768 3698 772
rect 3734 768 3738 772
rect 3814 768 3818 772
rect 4286 768 4290 772
rect 4310 768 4314 772
rect 4422 768 4426 772
rect 4558 768 4562 772
rect 4598 768 4602 772
rect 4614 768 4618 772
rect 4662 768 4666 772
rect 4686 768 4690 772
rect 4950 768 4954 772
rect 4990 768 4994 772
rect 5022 768 5026 772
rect 5126 768 5130 772
rect 5134 768 5138 772
rect 5150 768 5154 772
rect 5166 768 5170 772
rect 30 747 34 751
rect 62 748 66 752
rect 110 748 114 752
rect 134 748 138 752
rect 150 748 154 752
rect 174 748 178 752
rect 190 748 194 752
rect 246 758 250 762
rect 326 758 330 762
rect 390 758 394 762
rect 510 758 514 762
rect 550 758 554 762
rect 598 758 602 762
rect 926 758 930 762
rect 1054 758 1058 762
rect 1118 758 1122 762
rect 1190 758 1194 762
rect 1310 758 1314 762
rect 1342 758 1346 762
rect 1414 758 1418 762
rect 1486 758 1490 762
rect 1518 758 1522 762
rect 1526 758 1530 762
rect 1574 758 1578 762
rect 1902 758 1906 762
rect 1950 758 1954 762
rect 2086 758 2090 762
rect 2182 758 2186 762
rect 2254 758 2258 762
rect 2278 758 2282 762
rect 2430 758 2434 762
rect 2478 758 2482 762
rect 2510 758 2514 762
rect 2614 758 2618 762
rect 2694 758 2698 762
rect 3038 758 3042 762
rect 3118 758 3122 762
rect 3310 758 3314 762
rect 3350 758 3354 762
rect 3454 758 3458 762
rect 3502 758 3506 762
rect 3686 758 3690 762
rect 3710 758 3714 762
rect 3718 758 3722 762
rect 4054 758 4058 762
rect 4102 758 4106 762
rect 4270 758 4274 762
rect 4382 758 4386 762
rect 4398 758 4402 762
rect 4438 758 4442 762
rect 4494 758 4498 762
rect 4510 758 4514 762
rect 4542 758 4546 762
rect 4574 758 4578 762
rect 4582 758 4586 762
rect 4646 758 4650 762
rect 4782 758 4786 762
rect 4974 758 4978 762
rect 5006 758 5010 762
rect 5110 758 5114 762
rect 214 748 218 752
rect 270 748 274 752
rect 334 748 338 752
rect 414 748 418 752
rect 46 738 50 742
rect 102 738 106 742
rect 158 738 162 742
rect 182 738 186 742
rect 206 738 210 742
rect 222 738 226 742
rect 262 738 266 742
rect 502 748 506 752
rect 518 748 522 752
rect 582 748 586 752
rect 710 748 714 752
rect 766 748 770 752
rect 318 738 322 742
rect 374 738 378 742
rect 438 738 442 742
rect 454 738 458 742
rect 502 738 506 742
rect 526 738 530 742
rect 566 738 570 742
rect 798 747 802 751
rect 830 748 834 752
rect 1006 748 1010 752
rect 1054 748 1058 752
rect 1062 748 1066 752
rect 1094 748 1098 752
rect 1142 748 1146 752
rect 1174 748 1178 752
rect 1182 748 1186 752
rect 1230 748 1234 752
rect 1262 747 1266 751
rect 1350 748 1354 752
rect 1438 748 1442 752
rect 1454 748 1458 752
rect 1478 748 1482 752
rect 1542 748 1546 752
rect 1598 748 1602 752
rect 1694 748 1698 752
rect 1718 748 1722 752
rect 2006 748 2010 752
rect 2038 747 2042 751
rect 2238 748 2242 752
rect 2286 748 2290 752
rect 2310 748 2314 752
rect 2358 748 2362 752
rect 2422 748 2426 752
rect 2470 748 2474 752
rect 2534 748 2538 752
rect 2630 748 2634 752
rect 2710 748 2714 752
rect 2894 748 2898 752
rect 590 738 594 742
rect 654 738 658 742
rect 662 738 666 742
rect 814 738 818 742
rect 870 738 874 742
rect 918 738 922 742
rect 942 738 946 742
rect 950 738 954 742
rect 1030 738 1034 742
rect 1086 738 1090 742
rect 1294 738 1298 742
rect 1310 738 1314 742
rect 1326 738 1330 742
rect 1358 738 1362 742
rect 1366 738 1370 742
rect 1374 738 1378 742
rect 1438 738 1442 742
rect 1478 738 1482 742
rect 1550 738 1554 742
rect 1558 738 1562 742
rect 1590 738 1594 742
rect 1598 738 1602 742
rect 1654 738 1658 742
rect 1662 738 1666 742
rect 1710 738 1714 742
rect 1758 738 1762 742
rect 1806 738 1810 742
rect 1814 738 1818 742
rect 1862 738 1866 742
rect 1934 738 1938 742
rect 2070 738 2074 742
rect 2086 738 2090 742
rect 2110 738 2114 742
rect 2158 738 2162 742
rect 2214 738 2218 742
rect 2238 738 2242 742
rect 2254 738 2258 742
rect 2366 738 2370 742
rect 2454 738 2458 742
rect 2462 738 2466 742
rect 2502 738 2506 742
rect 2550 738 2554 742
rect 2934 747 2938 751
rect 2966 748 2970 752
rect 3054 748 3058 752
rect 3134 748 3138 752
rect 3174 748 3178 752
rect 3182 748 3186 752
rect 3190 748 3194 752
rect 2638 738 2642 742
rect 2718 738 2722 742
rect 2726 738 2730 742
rect 2774 738 2778 742
rect 2782 738 2786 742
rect 2830 738 2834 742
rect 2838 738 2842 742
rect 2886 738 2890 742
rect 3054 738 3058 742
rect 3230 747 3234 751
rect 3262 748 3266 752
rect 3326 748 3330 752
rect 3374 748 3378 752
rect 3422 748 3426 752
rect 3462 748 3466 752
rect 3526 748 3530 752
rect 3630 748 3634 752
rect 3726 748 3730 752
rect 3830 748 3834 752
rect 3870 748 3874 752
rect 3910 748 3914 752
rect 4150 748 4154 752
rect 4198 747 4202 751
rect 4278 748 4282 752
rect 4318 748 4322 752
rect 4382 748 4386 752
rect 4398 748 4402 752
rect 4430 748 4434 752
rect 4470 748 4474 752
rect 4478 748 4482 752
rect 4494 748 4498 752
rect 4526 748 4530 752
rect 4534 748 4538 752
rect 4566 748 4570 752
rect 4590 748 4594 752
rect 4638 748 4642 752
rect 4654 748 4658 752
rect 4694 748 4698 752
rect 4726 748 4730 752
rect 4742 748 4746 752
rect 4790 748 4794 752
rect 4854 748 4858 752
rect 4886 748 4890 752
rect 4934 748 4938 752
rect 4982 748 4986 752
rect 5014 748 5018 752
rect 5038 748 5042 752
rect 5078 748 5082 752
rect 5118 748 5122 752
rect 5126 748 5130 752
rect 5182 748 5186 752
rect 5206 748 5210 752
rect 3110 738 3114 742
rect 3126 738 3130 742
rect 3150 738 3154 742
rect 3166 738 3170 742
rect 3214 738 3218 742
rect 3318 738 3322 742
rect 3382 738 3386 742
rect 3390 738 3394 742
rect 3406 738 3410 742
rect 3430 738 3434 742
rect 3470 738 3474 742
rect 3526 738 3530 742
rect 3574 738 3578 742
rect 3582 738 3586 742
rect 3654 738 3658 742
rect 3750 738 3754 742
rect 3806 738 3810 742
rect 3862 738 3866 742
rect 3894 738 3898 742
rect 4022 738 4026 742
rect 4030 738 4034 742
rect 4078 738 4082 742
rect 4086 738 4090 742
rect 4126 738 4130 742
rect 4134 738 4138 742
rect 4182 738 4186 742
rect 4374 738 4378 742
rect 4406 738 4410 742
rect 4478 738 4482 742
rect 4518 738 4522 742
rect 4630 738 4634 742
rect 4750 738 4754 742
rect 4798 738 4802 742
rect 4910 738 4914 742
rect 4950 738 4954 742
rect 5094 738 5098 742
rect 5110 738 5114 742
rect 5246 738 5250 742
rect 5302 738 5306 742
rect 174 728 178 732
rect 238 728 242 732
rect 334 728 338 732
rect 382 728 386 732
rect 398 728 402 732
rect 438 728 442 732
rect 478 728 482 732
rect 542 728 546 732
rect 550 728 554 732
rect 1022 728 1026 732
rect 1118 728 1122 732
rect 1182 728 1186 732
rect 1318 728 1322 732
rect 1374 728 1378 732
rect 1406 728 1410 732
rect 1454 728 1458 732
rect 1494 728 1498 732
rect 1510 728 1514 732
rect 1582 728 1586 732
rect 1750 728 1754 732
rect 1886 728 1890 732
rect 1910 728 1914 732
rect 1926 728 1930 732
rect 2038 728 2042 732
rect 2102 728 2106 732
rect 2174 728 2178 732
rect 2190 728 2194 732
rect 2206 728 2210 732
rect 2262 728 2266 732
rect 2310 728 2314 732
rect 2326 728 2330 732
rect 2374 728 2378 732
rect 2422 728 2426 732
rect 2430 728 2434 732
rect 2446 728 2450 732
rect 2646 728 2650 732
rect 2662 728 2666 732
rect 2670 728 2674 732
rect 3150 728 3154 732
rect 3198 728 3202 732
rect 3406 728 3410 732
rect 3454 728 3458 732
rect 3486 728 3490 732
rect 3662 728 3666 732
rect 3918 728 3922 732
rect 4134 728 4138 732
rect 4342 728 4346 732
rect 4446 728 4450 732
rect 4462 728 4466 732
rect 4614 728 4618 732
rect 4710 728 4714 732
rect 4814 728 4818 732
rect 4870 728 4874 732
rect 4902 728 4906 732
rect 4950 728 4954 732
rect 5054 728 5058 732
rect 94 718 98 722
rect 126 718 130 722
rect 230 718 234 722
rect 446 718 450 722
rect 534 718 538 722
rect 902 718 906 722
rect 934 718 938 722
rect 1574 718 1578 722
rect 2590 718 2594 722
rect 2758 718 2762 722
rect 3094 718 3098 722
rect 3158 718 3162 722
rect 3366 718 3370 722
rect 3478 718 3482 722
rect 3758 718 3762 722
rect 3774 718 3778 722
rect 3886 718 3890 722
rect 3894 718 3898 722
rect 3926 718 3930 722
rect 4086 718 4090 722
rect 4102 718 4106 722
rect 4110 718 4114 722
rect 4166 718 4170 722
rect 5046 718 5050 722
rect 5062 718 5066 722
rect 5094 718 5098 722
rect 614 708 618 712
rect 4134 708 4138 712
rect 4646 708 4650 712
rect 4710 708 4714 712
rect 4814 708 4818 712
rect 4902 708 4906 712
rect 5054 708 5058 712
rect 858 703 862 707
rect 865 703 869 707
rect 1874 703 1878 707
rect 1881 703 1885 707
rect 2906 703 2910 707
rect 2913 703 2917 707
rect 3930 703 3934 707
rect 3937 703 3941 707
rect 4954 703 4958 707
rect 4961 703 4965 707
rect 102 698 106 702
rect 238 698 242 702
rect 1654 698 1658 702
rect 3870 698 3874 702
rect 4254 698 4258 702
rect 4702 698 4706 702
rect 4758 698 4762 702
rect 4854 698 4858 702
rect 142 688 146 692
rect 214 688 218 692
rect 278 688 282 692
rect 358 688 362 692
rect 398 688 402 692
rect 454 688 458 692
rect 486 688 490 692
rect 630 688 634 692
rect 790 688 794 692
rect 934 688 938 692
rect 942 688 946 692
rect 1142 688 1146 692
rect 1166 688 1170 692
rect 1190 688 1194 692
rect 1206 688 1210 692
rect 1254 688 1258 692
rect 1470 688 1474 692
rect 1686 688 1690 692
rect 1710 688 1714 692
rect 1758 688 1762 692
rect 1854 688 1858 692
rect 1926 688 1930 692
rect 1966 688 1970 692
rect 2110 688 2114 692
rect 2150 688 2154 692
rect 2278 688 2282 692
rect 2318 688 2322 692
rect 2462 688 2466 692
rect 2590 688 2594 692
rect 2670 688 2674 692
rect 2726 688 2730 692
rect 2766 688 2770 692
rect 2814 688 2818 692
rect 2830 688 2834 692
rect 2854 688 2858 692
rect 2934 688 2938 692
rect 3054 688 3058 692
rect 3126 688 3130 692
rect 3310 688 3314 692
rect 3326 688 3330 692
rect 3430 688 3434 692
rect 3446 688 3450 692
rect 3654 688 3658 692
rect 3806 688 3810 692
rect 4070 688 4074 692
rect 4302 688 4306 692
rect 4318 688 4322 692
rect 4342 688 4346 692
rect 4382 688 4386 692
rect 4398 688 4402 692
rect 4470 688 4474 692
rect 4566 688 4570 692
rect 4614 688 4618 692
rect 4654 688 4658 692
rect 4670 688 4674 692
rect 4678 688 4682 692
rect 4734 688 4738 692
rect 4798 688 4802 692
rect 4846 688 4850 692
rect 4902 688 4906 692
rect 4926 688 4930 692
rect 4974 688 4978 692
rect 4990 688 4994 692
rect 5198 688 5202 692
rect 14 679 18 683
rect 62 679 66 683
rect 86 679 90 683
rect 150 678 154 682
rect 238 678 242 682
rect 270 678 274 682
rect 446 678 450 682
rect 478 678 482 682
rect 870 678 874 682
rect 1022 678 1026 682
rect 1110 678 1114 682
rect 1134 678 1138 682
rect 1158 678 1162 682
rect 1974 678 1978 682
rect 2286 678 2290 682
rect 2430 678 2434 682
rect 2486 678 2490 682
rect 2614 678 2618 682
rect 2646 678 2650 682
rect 3670 679 3674 683
rect 3782 678 3786 682
rect 3798 678 3802 682
rect 3870 678 3874 682
rect 3990 678 3994 682
rect 4062 678 4066 682
rect 4158 678 4162 682
rect 4254 678 4258 682
rect 4366 678 4370 682
rect 4702 678 4706 682
rect 4742 678 4746 682
rect 4758 678 4762 682
rect 4854 678 4858 682
rect 4942 678 4946 682
rect 5038 678 5042 682
rect 5086 678 5090 682
rect 5094 678 5098 682
rect 5166 678 5170 682
rect 158 668 162 672
rect 166 668 170 672
rect 190 668 194 672
rect 206 668 210 672
rect 214 668 218 672
rect 230 668 234 672
rect 286 668 290 672
rect 478 668 482 672
rect 494 668 498 672
rect 526 668 530 672
rect 558 668 562 672
rect 590 668 594 672
rect 598 668 602 672
rect 654 668 658 672
rect 702 668 706 672
rect 710 668 714 672
rect 782 668 786 672
rect 846 668 850 672
rect 886 668 890 672
rect 902 668 906 672
rect 958 668 962 672
rect 990 668 994 672
rect 1030 668 1034 672
rect 1046 668 1050 672
rect 1078 668 1082 672
rect 1198 668 1202 672
rect 1230 668 1234 672
rect 1238 668 1242 672
rect 1262 668 1266 672
rect 1310 668 1314 672
rect 1318 668 1322 672
rect 1366 668 1370 672
rect 1390 668 1394 672
rect 1438 668 1442 672
rect 1446 668 1450 672
rect 1494 668 1498 672
rect 1502 668 1506 672
rect 1566 668 1570 672
rect 1622 668 1626 672
rect 1670 668 1674 672
rect 1718 668 1722 672
rect 1726 668 1730 672
rect 1774 668 1778 672
rect 22 658 26 662
rect 54 658 58 662
rect 78 658 82 662
rect 134 658 138 662
rect 190 658 194 662
rect 214 658 218 662
rect 294 658 298 662
rect 310 658 314 662
rect 358 658 362 662
rect 390 658 394 662
rect 430 658 434 662
rect 470 658 474 662
rect 502 658 506 662
rect 534 658 538 662
rect 550 658 554 662
rect 814 658 818 662
rect 838 658 842 662
rect 854 658 858 662
rect 870 658 874 662
rect 918 658 922 662
rect 982 658 986 662
rect 1006 658 1010 662
rect 1054 658 1058 662
rect 1094 658 1098 662
rect 1118 658 1122 662
rect 1126 658 1130 662
rect 1150 658 1154 662
rect 1174 658 1178 662
rect 1222 658 1226 662
rect 1278 658 1282 662
rect 1422 658 1426 662
rect 1638 659 1642 663
rect 1774 658 1778 662
rect 1830 668 1834 672
rect 1838 668 1842 672
rect 1894 668 1898 672
rect 1910 668 1914 672
rect 1958 668 1962 672
rect 2038 668 2042 672
rect 2062 668 2066 672
rect 2078 668 2082 672
rect 2126 668 2130 672
rect 2134 668 2138 672
rect 2182 668 2186 672
rect 2198 668 2202 672
rect 2294 668 2298 672
rect 2350 668 2354 672
rect 2366 668 2370 672
rect 2438 668 2442 672
rect 2518 668 2522 672
rect 2606 668 2610 672
rect 2630 668 2634 672
rect 2654 668 2658 672
rect 2710 668 2714 672
rect 2726 668 2730 672
rect 2758 668 2762 672
rect 2782 668 2786 672
rect 2790 668 2794 672
rect 1798 658 1802 662
rect 2030 658 2034 662
rect 2222 658 2226 662
rect 2334 658 2338 662
rect 2390 658 2394 662
rect 2446 658 2450 662
rect 2470 658 2474 662
rect 2486 658 2490 662
rect 2510 658 2514 662
rect 2550 658 2554 662
rect 2566 658 2570 662
rect 2798 666 2802 670
rect 2822 668 2826 672
rect 2862 668 2866 672
rect 2910 668 2914 672
rect 2998 668 3002 672
rect 2686 658 2690 662
rect 2734 658 2738 662
rect 2822 658 2826 662
rect 2870 658 2874 662
rect 2886 658 2890 662
rect 2966 658 2970 662
rect 3038 668 3042 672
rect 3086 668 3090 672
rect 3094 668 3098 672
rect 3142 668 3146 672
rect 3214 668 3218 672
rect 3230 668 3234 672
rect 3334 668 3338 672
rect 3350 668 3354 672
rect 3742 668 3746 672
rect 3774 668 3778 672
rect 3878 668 3882 672
rect 3910 668 3914 672
rect 3974 668 3978 672
rect 3998 668 4002 672
rect 4078 668 4082 672
rect 4166 668 4170 672
rect 4198 668 4202 672
rect 4230 668 4234 672
rect 4262 668 4266 672
rect 4310 668 4314 672
rect 4334 668 4338 672
rect 4358 668 4362 672
rect 4422 668 4426 672
rect 4430 668 4434 672
rect 4446 668 4450 672
rect 4454 666 4458 670
rect 4486 668 4490 672
rect 4574 668 4578 672
rect 4622 668 4626 672
rect 4670 668 4674 672
rect 4694 668 4698 672
rect 4710 668 4714 672
rect 4766 668 4770 672
rect 4814 668 4818 672
rect 4862 668 4866 672
rect 4902 668 4906 672
rect 4918 668 4922 672
rect 5030 668 5034 672
rect 5054 668 5058 672
rect 5070 668 5074 672
rect 3014 658 3018 662
rect 3030 658 3034 662
rect 3158 658 3162 662
rect 3254 658 3258 662
rect 3366 659 3370 663
rect 3390 658 3394 662
rect 3486 658 3490 662
rect 3510 658 3514 662
rect 3574 659 3578 663
rect 3678 658 3682 662
rect 3702 658 3706 662
rect 3718 658 3722 662
rect 3734 658 3738 662
rect 3766 658 3770 662
rect 3782 658 3786 662
rect 3822 658 3826 662
rect 3830 658 3834 662
rect 3846 658 3850 662
rect 3918 658 3922 662
rect 3942 658 3946 662
rect 3966 658 3970 662
rect 3974 658 3978 662
rect 4006 658 4010 662
rect 4046 658 4050 662
rect 4086 658 4090 662
rect 4102 658 4106 662
rect 4142 658 4146 662
rect 4190 658 4194 662
rect 4222 658 4226 662
rect 4238 658 4242 662
rect 4254 658 4258 662
rect 4390 658 4394 662
rect 4414 658 4418 662
rect 4502 659 4506 663
rect 4622 658 4626 662
rect 4646 658 4650 662
rect 4718 658 4722 662
rect 4742 658 4746 662
rect 4830 658 4834 662
rect 4910 658 4914 662
rect 4974 658 4978 662
rect 5022 658 5026 662
rect 5158 658 5162 662
rect 5230 658 5234 662
rect 5254 658 5258 662
rect 230 648 234 652
rect 262 648 266 652
rect 302 648 306 652
rect 342 648 346 652
rect 358 648 362 652
rect 406 648 410 652
rect 414 648 418 652
rect 430 648 434 652
rect 510 648 514 652
rect 534 648 538 652
rect 550 648 554 652
rect 590 648 594 652
rect 798 648 802 652
rect 806 648 810 652
rect 902 648 906 652
rect 942 648 946 652
rect 966 648 970 652
rect 1022 648 1026 652
rect 1070 648 1074 652
rect 1102 648 1106 652
rect 1182 648 1186 652
rect 1254 648 1258 652
rect 2342 648 2346 652
rect 2350 648 2354 652
rect 2366 648 2370 652
rect 2430 648 2434 652
rect 2494 648 2498 652
rect 2550 648 2554 652
rect 2582 648 2586 652
rect 2670 648 2674 652
rect 2678 648 2682 652
rect 2710 648 2714 652
rect 2726 648 2730 652
rect 2766 648 2770 652
rect 2838 648 2842 652
rect 2878 648 2882 652
rect 2950 648 2954 652
rect 2982 648 2986 652
rect 3030 648 3034 652
rect 3318 648 3322 652
rect 3710 648 3714 652
rect 3718 648 3722 652
rect 3750 648 3754 652
rect 3798 648 3802 652
rect 3838 648 3842 652
rect 3950 648 3954 652
rect 4022 648 4026 652
rect 4054 648 4058 652
rect 4094 648 4098 652
rect 4174 648 4178 652
rect 4206 648 4210 652
rect 4318 648 4322 652
rect 4654 648 4658 652
rect 4878 648 4882 652
rect 4886 648 4890 652
rect 4982 648 4986 652
rect 318 638 322 642
rect 390 638 394 642
rect 982 638 986 642
rect 2310 638 2314 642
rect 2326 638 2330 642
rect 2382 638 2386 642
rect 2390 638 2394 642
rect 2510 638 2514 642
rect 2566 638 2570 642
rect 2694 638 2698 642
rect 2886 638 2890 642
rect 2894 638 2898 642
rect 2942 638 2946 642
rect 3694 638 3698 642
rect 3854 638 3858 642
rect 3894 638 3898 642
rect 3910 638 3914 642
rect 4006 638 4010 642
rect 4038 638 4042 642
rect 4110 638 4114 642
rect 4134 638 4138 642
rect 4294 638 4298 642
rect 4966 638 4970 642
rect 5102 638 5106 642
rect 2574 628 2578 632
rect 2646 628 2650 632
rect 3830 628 3834 632
rect 4222 628 4226 632
rect 678 618 682 622
rect 766 618 770 622
rect 830 618 834 622
rect 1350 618 1354 622
rect 1574 618 1578 622
rect 1982 618 1986 622
rect 3686 618 3690 622
rect 3766 618 3770 622
rect 3846 618 3850 622
rect 4030 618 4034 622
rect 4102 618 4106 622
rect 4142 618 4146 622
rect 4190 618 4194 622
rect 4462 608 4466 612
rect 346 603 350 607
rect 353 603 357 607
rect 1370 603 1374 607
rect 1377 603 1381 607
rect 2394 603 2398 607
rect 2401 603 2405 607
rect 3418 603 3422 607
rect 3425 603 3429 607
rect 4442 603 4446 607
rect 4449 603 4453 607
rect 222 588 226 592
rect 270 588 274 592
rect 414 588 418 592
rect 438 588 442 592
rect 486 588 490 592
rect 518 588 522 592
rect 598 588 602 592
rect 646 588 650 592
rect 798 588 802 592
rect 902 588 906 592
rect 1038 588 1042 592
rect 1102 588 1106 592
rect 1126 588 1130 592
rect 1446 588 1450 592
rect 1478 588 1482 592
rect 1606 588 1610 592
rect 1662 588 1666 592
rect 1726 588 1730 592
rect 1990 588 1994 592
rect 2006 588 2010 592
rect 2118 588 2122 592
rect 2462 588 2466 592
rect 2534 588 2538 592
rect 2654 588 2658 592
rect 2742 588 2746 592
rect 2758 588 2762 592
rect 2814 588 2818 592
rect 3030 588 3034 592
rect 3094 588 3098 592
rect 3374 588 3378 592
rect 3678 588 3682 592
rect 3694 588 3698 592
rect 3886 588 3890 592
rect 3894 588 3898 592
rect 5270 588 5274 592
rect 3750 578 3754 582
rect 3846 578 3850 582
rect 3854 578 3858 582
rect 5046 578 5050 582
rect 214 568 218 572
rect 486 568 490 572
rect 526 568 530 572
rect 566 568 570 572
rect 638 568 642 572
rect 774 568 778 572
rect 822 568 826 572
rect 1094 568 1098 572
rect 1894 568 1898 572
rect 1926 568 1930 572
rect 2358 568 2362 572
rect 2430 568 2434 572
rect 2518 568 2522 572
rect 2542 568 2546 572
rect 2606 568 2610 572
rect 2614 568 2618 572
rect 2646 568 2650 572
rect 2990 568 2994 572
rect 3038 568 3042 572
rect 3102 568 3106 572
rect 3238 568 3242 572
rect 3318 568 3322 572
rect 3510 568 3514 572
rect 3670 568 3674 572
rect 3726 568 3730 572
rect 3750 568 3754 572
rect 3758 568 3762 572
rect 3902 568 3906 572
rect 3926 568 3930 572
rect 4374 568 4378 572
rect 4422 568 4426 572
rect 4550 568 4554 572
rect 4854 568 4858 572
rect 5078 568 5082 572
rect 5278 568 5282 572
rect 182 558 186 562
rect 198 558 202 562
rect 398 558 402 562
rect 510 558 514 562
rect 654 558 658 562
rect 742 558 746 562
rect 750 558 754 562
rect 766 558 770 562
rect 910 558 914 562
rect 934 558 938 562
rect 1078 558 1082 562
rect 1470 558 1474 562
rect 1702 558 1706 562
rect 1854 558 1858 562
rect 2374 558 2378 562
rect 2446 558 2450 562
rect 2558 558 2562 562
rect 2598 558 2602 562
rect 2630 558 2634 562
rect 2830 558 2834 562
rect 2854 558 2858 562
rect 3022 558 3026 562
rect 3054 558 3058 562
rect 3086 558 3090 562
rect 3174 558 3178 562
rect 3262 558 3266 562
rect 3278 558 3282 562
rect 3582 558 3586 562
rect 3638 558 3642 562
rect 3702 558 3706 562
rect 3718 558 3722 562
rect 3742 558 3746 562
rect 3774 558 3778 562
rect 3830 558 3834 562
rect 3910 558 3914 562
rect 4518 558 4522 562
rect 4534 558 4538 562
rect 4566 558 4570 562
rect 4870 558 4874 562
rect 4878 558 4882 562
rect 5022 558 5026 562
rect 5174 558 5178 562
rect 5294 558 5298 562
rect 22 548 26 552
rect 62 548 66 552
rect 142 548 146 552
rect 198 548 202 552
rect 222 548 226 552
rect 238 548 242 552
rect 270 548 274 552
rect 318 548 322 552
rect 414 548 418 552
rect 494 548 498 552
rect 518 548 522 552
rect 542 548 546 552
rect 646 548 650 552
rect 678 548 682 552
rect 686 548 690 552
rect 710 548 714 552
rect 782 548 786 552
rect 862 548 866 552
rect 990 548 994 552
rect 1086 548 1090 552
rect 1198 548 1202 552
rect 38 538 42 542
rect 158 538 162 542
rect 182 538 186 542
rect 1230 547 1234 551
rect 1334 548 1338 552
rect 1550 548 1554 552
rect 1798 548 1802 552
rect 1838 548 1842 552
rect 1862 548 1866 552
rect 1878 548 1882 552
rect 1918 548 1922 552
rect 1950 548 1954 552
rect 2062 548 2066 552
rect 278 538 282 542
rect 294 538 298 542
rect 430 538 434 542
rect 550 538 554 542
rect 574 538 578 542
rect 622 538 626 542
rect 694 538 698 542
rect 718 538 722 542
rect 766 538 770 542
rect 870 538 874 542
rect 910 538 914 542
rect 966 538 970 542
rect 1030 538 1034 542
rect 1110 538 1114 542
rect 1158 538 1162 542
rect 1262 538 1266 542
rect 1310 538 1314 542
rect 1342 538 1346 542
rect 1406 538 1410 542
rect 1414 538 1418 542
rect 1462 538 1466 542
rect 1486 538 1490 542
rect 1494 538 1498 542
rect 1574 538 1578 542
rect 1622 538 1626 542
rect 1678 538 1682 542
rect 1686 538 1690 542
rect 2086 547 2090 551
rect 2174 548 2178 552
rect 2230 548 2234 552
rect 2286 548 2290 552
rect 2310 548 2314 552
rect 2430 548 2434 552
rect 2462 548 2466 552
rect 2510 548 2514 552
rect 2526 548 2530 552
rect 2550 548 2554 552
rect 2566 548 2570 552
rect 2606 548 2610 552
rect 2622 548 2626 552
rect 2638 548 2642 552
rect 2694 548 2698 552
rect 2718 548 2722 552
rect 2734 548 2738 552
rect 2782 548 2786 552
rect 2814 548 2818 552
rect 2894 548 2898 552
rect 2942 548 2946 552
rect 2958 548 2962 552
rect 2974 548 2978 552
rect 3006 548 3010 552
rect 3046 548 3050 552
rect 3094 548 3098 552
rect 3166 548 3170 552
rect 3198 548 3202 552
rect 3398 548 3402 552
rect 3566 548 3570 552
rect 3630 548 3634 552
rect 3678 548 3682 552
rect 3718 548 3722 552
rect 3750 548 3754 552
rect 3774 548 3778 552
rect 3798 548 3802 552
rect 3902 548 3906 552
rect 3934 548 3938 552
rect 3982 548 3986 552
rect 4022 548 4026 552
rect 4030 548 4034 552
rect 4078 548 4082 552
rect 4086 548 4090 552
rect 4110 548 4114 552
rect 1830 538 1834 542
rect 1846 538 1850 542
rect 1926 538 1930 542
rect 1974 538 1978 542
rect 1982 538 1986 542
rect 2166 538 2170 542
rect 2238 538 2242 542
rect 2286 538 2290 542
rect 2318 538 2322 542
rect 2334 538 2338 542
rect 2358 538 2362 542
rect 2414 538 2418 542
rect 2454 538 2458 542
rect 2574 538 2578 542
rect 2662 538 2666 542
rect 2710 538 2714 542
rect 2718 538 2722 542
rect 2806 538 2810 542
rect 2838 538 2842 542
rect 2958 538 2962 542
rect 3014 538 3018 542
rect 3062 538 3066 542
rect 3078 538 3082 542
rect 3118 538 3122 542
rect 3166 538 3170 542
rect 3198 538 3202 542
rect 3206 538 3210 542
rect 3262 538 3266 542
rect 3334 538 3338 542
rect 3342 538 3346 542
rect 3390 538 3394 542
rect 3438 538 3442 542
rect 3486 538 3490 542
rect 3494 538 3498 542
rect 3542 538 3546 542
rect 3582 538 3586 542
rect 3606 538 3610 542
rect 3638 538 3642 542
rect 3654 538 3658 542
rect 3790 538 3794 542
rect 3806 538 3810 542
rect 3830 538 3834 542
rect 3846 538 3850 542
rect 3870 538 3874 542
rect 3926 538 3930 542
rect 3950 538 3954 542
rect 4158 548 4162 552
rect 4198 548 4202 552
rect 4262 548 4266 552
rect 4270 548 4274 552
rect 4302 548 4306 552
rect 4318 548 4322 552
rect 4358 548 4362 552
rect 4390 548 4394 552
rect 4518 548 4522 552
rect 4558 548 4562 552
rect 4070 538 4074 542
rect 4134 538 4138 542
rect 4150 538 4154 542
rect 4206 538 4210 542
rect 4270 538 4274 542
rect 4326 538 4330 542
rect 4334 538 4338 542
rect 4382 538 4386 542
rect 4414 538 4418 542
rect 4462 538 4466 542
rect 4494 538 4498 542
rect 4518 538 4522 542
rect 4630 548 4634 552
rect 4670 548 4674 552
rect 4702 548 4706 552
rect 4726 548 4730 552
rect 4750 548 4754 552
rect 4790 548 4794 552
rect 4838 548 4842 552
rect 4862 548 4866 552
rect 4894 548 4898 552
rect 5014 548 5018 552
rect 5038 548 5042 552
rect 5046 548 5050 552
rect 5110 548 5114 552
rect 4590 538 4594 542
rect 4638 538 4642 542
rect 5142 547 5146 551
rect 5206 548 5210 552
rect 5238 547 5242 551
rect 5286 548 5290 552
rect 4734 538 4738 542
rect 4742 538 4746 542
rect 4830 538 4834 542
rect 4878 538 4882 542
rect 4894 538 4898 542
rect 4902 538 4906 542
rect 4950 538 4954 542
rect 5054 540 5058 544
rect 14 527 18 531
rect 150 528 154 532
rect 238 528 242 532
rect 462 528 466 532
rect 566 528 570 532
rect 710 528 714 532
rect 718 528 722 532
rect 750 528 754 532
rect 806 528 810 532
rect 838 528 842 532
rect 878 528 882 532
rect 894 528 898 532
rect 958 528 962 532
rect 982 528 986 532
rect 1014 528 1018 532
rect 1070 528 1074 532
rect 1814 528 1818 532
rect 1862 528 1866 532
rect 1942 528 1946 532
rect 1958 527 1962 531
rect 1998 528 2002 532
rect 2014 528 2018 532
rect 2398 528 2402 532
rect 2486 528 2490 532
rect 2590 528 2594 532
rect 2750 528 2754 532
rect 2798 528 2802 532
rect 2926 528 2930 532
rect 2942 528 2946 532
rect 3174 528 3178 532
rect 3406 527 3410 531
rect 3590 528 3594 532
rect 3606 528 3610 532
rect 3702 528 3706 532
rect 3822 528 3826 532
rect 3878 528 3882 532
rect 3958 528 3962 532
rect 3966 528 3970 532
rect 3998 528 4002 532
rect 4006 528 4010 532
rect 4046 528 4050 532
rect 4054 528 4058 532
rect 4094 527 4098 531
rect 4134 528 4138 532
rect 4174 528 4178 532
rect 4222 528 4226 532
rect 4278 528 4282 532
rect 4294 528 4298 532
rect 4486 528 4490 532
rect 4590 528 4594 532
rect 4598 528 4602 532
rect 4606 528 4610 532
rect 4654 528 4658 532
rect 4774 528 4778 532
rect 4814 528 4818 532
rect 5022 528 5026 532
rect 118 518 122 522
rect 182 518 186 522
rect 246 518 250 522
rect 454 518 458 522
rect 614 518 618 522
rect 1166 518 1170 522
rect 1294 518 1298 522
rect 1358 518 1362 522
rect 1526 518 1530 522
rect 1694 518 1698 522
rect 1790 518 1794 522
rect 2022 518 2026 522
rect 2270 518 2274 522
rect 2278 518 2282 522
rect 2374 518 2378 522
rect 2718 518 2722 522
rect 2838 518 2842 522
rect 2854 518 2858 522
rect 2870 518 2874 522
rect 2958 518 2962 522
rect 3158 518 3162 522
rect 3230 518 3234 522
rect 3454 518 3458 522
rect 3614 518 3618 522
rect 3638 518 3642 522
rect 3718 518 3722 522
rect 3814 518 3818 522
rect 4038 518 4042 522
rect 4246 518 4250 522
rect 4342 518 4346 522
rect 4446 518 4450 522
rect 4518 518 4522 522
rect 4558 518 4562 522
rect 4614 518 4618 522
rect 4662 518 4666 522
rect 4766 518 4770 522
rect 4782 518 4786 522
rect 4790 518 4794 522
rect 4798 518 4802 522
rect 4822 518 4826 522
rect 4862 518 4866 522
rect 4894 518 4898 522
rect 5030 518 5034 522
rect 5038 518 5042 522
rect 5070 518 5074 522
rect 134 508 138 512
rect 150 508 154 512
rect 1614 508 1618 512
rect 1862 508 1866 512
rect 2942 508 2946 512
rect 4294 508 4298 512
rect 4486 508 4490 512
rect 4590 508 4594 512
rect 4774 508 4778 512
rect 4910 508 4914 512
rect 858 503 862 507
rect 865 503 869 507
rect 1874 503 1878 507
rect 1881 503 1885 507
rect 2906 503 2910 507
rect 2913 503 2917 507
rect 3930 503 3934 507
rect 3937 503 3941 507
rect 4954 503 4958 507
rect 4961 503 4965 507
rect 142 498 146 502
rect 238 498 242 502
rect 422 498 426 502
rect 462 498 466 502
rect 1926 498 1930 502
rect 2230 498 2234 502
rect 2630 498 2634 502
rect 2958 498 2962 502
rect 3222 498 3226 502
rect 4198 498 4202 502
rect 4390 498 4394 502
rect 4534 498 4538 502
rect 4734 498 4738 502
rect 5046 498 5050 502
rect 110 488 114 492
rect 158 488 162 492
rect 294 488 298 492
rect 358 488 362 492
rect 414 488 418 492
rect 430 488 434 492
rect 486 488 490 492
rect 494 488 498 492
rect 510 488 514 492
rect 606 488 610 492
rect 630 488 634 492
rect 662 488 666 492
rect 702 488 706 492
rect 790 488 794 492
rect 846 488 850 492
rect 966 488 970 492
rect 1222 488 1226 492
rect 1318 488 1322 492
rect 1406 488 1410 492
rect 1542 488 1546 492
rect 1590 488 1594 492
rect 1622 488 1626 492
rect 1774 488 1778 492
rect 1870 488 1874 492
rect 2006 488 2010 492
rect 2054 488 2058 492
rect 2102 488 2106 492
rect 2278 488 2282 492
rect 2526 488 2530 492
rect 2614 488 2618 492
rect 2622 488 2626 492
rect 2670 488 2674 492
rect 2710 488 2714 492
rect 2790 488 2794 492
rect 2862 488 2866 492
rect 2878 488 2882 492
rect 2926 488 2930 492
rect 3166 488 3170 492
rect 3390 488 3394 492
rect 3774 488 3778 492
rect 3966 488 3970 492
rect 3998 488 4002 492
rect 4222 488 4226 492
rect 4846 488 4850 492
rect 14 479 18 483
rect 62 479 66 483
rect 238 478 242 482
rect 246 478 250 482
rect 422 478 426 482
rect 462 478 466 482
rect 670 478 674 482
rect 758 478 762 482
rect 822 478 826 482
rect 870 478 874 482
rect 1006 478 1010 482
rect 1270 478 1274 482
rect 1566 478 1570 482
rect 1734 478 1738 482
rect 1926 478 1930 482
rect 2630 478 2634 482
rect 2662 478 2666 482
rect 2718 478 2722 482
rect 2758 478 2762 482
rect 2774 478 2778 482
rect 2782 478 2786 482
rect 2918 478 2922 482
rect 2958 478 2962 482
rect 3470 478 3474 482
rect 3694 478 3698 482
rect 3726 478 3730 482
rect 3758 478 3762 482
rect 3766 478 3770 482
rect 3990 478 3994 482
rect 4054 478 4058 482
rect 4110 478 4114 482
rect 4198 478 4202 482
rect 4238 479 4242 483
rect 4478 478 4482 482
rect 4694 478 4698 482
rect 4734 478 4738 482
rect 4798 478 4802 482
rect 4870 478 4874 482
rect 4902 478 4906 482
rect 4982 478 4986 482
rect 5070 478 5074 482
rect 5278 478 5282 482
rect 78 468 82 472
rect 134 468 138 472
rect 182 468 186 472
rect 190 468 194 472
rect 198 466 202 470
rect 270 468 274 472
rect 350 468 354 472
rect 398 468 402 472
rect 462 468 466 472
rect 470 468 474 472
rect 510 468 514 472
rect 526 468 530 472
rect 646 468 650 472
rect 710 468 714 472
rect 766 468 770 472
rect 798 468 802 472
rect 926 468 930 472
rect 942 468 946 472
rect 998 468 1002 472
rect 1078 468 1082 472
rect 1190 468 1194 472
rect 1206 468 1210 472
rect 1262 468 1266 472
rect 1350 468 1354 472
rect 1374 468 1378 472
rect 1422 468 1426 472
rect 1438 468 1442 472
rect 1558 468 1562 472
rect 1598 468 1602 472
rect 1718 468 1722 472
rect 1742 468 1746 472
rect 1822 468 1826 472
rect 1862 468 1866 472
rect 1918 468 1922 472
rect 1934 468 1938 472
rect 2006 468 2010 472
rect 2014 468 2018 472
rect 2062 468 2066 472
rect 2070 468 2074 472
rect 2166 468 2170 472
rect 2206 468 2210 472
rect 2222 468 2226 472
rect 2270 468 2274 472
rect 2278 468 2282 472
rect 2350 468 2354 472
rect 2446 468 2450 472
rect 2542 468 2546 472
rect 2630 468 2634 472
rect 2678 468 2682 472
rect 2702 468 2706 472
rect 2734 468 2738 472
rect 2750 468 2754 472
rect 2774 468 2778 472
rect 2798 468 2802 472
rect 2814 468 2818 472
rect 2846 468 2850 472
rect 2950 468 2954 472
rect 3102 468 3106 472
rect 3174 468 3178 472
rect 3238 468 3242 472
rect 3246 468 3250 472
rect 3294 468 3298 472
rect 3310 468 3314 472
rect 3414 468 3418 472
rect 3462 468 3466 472
rect 3502 468 3506 472
rect 3558 468 3562 472
rect 3566 468 3570 472
rect 3574 468 3578 472
rect 3590 468 3594 472
rect 3654 468 3658 472
rect 3662 468 3666 472
rect 3750 468 3754 472
rect 3782 468 3786 472
rect 3798 468 3802 472
rect 3846 468 3850 472
rect 3886 468 3890 472
rect 3918 468 3922 472
rect 3934 468 3938 472
rect 4006 468 4010 472
rect 4022 468 4026 472
rect 4046 468 4050 472
rect 4102 468 4106 472
rect 4126 468 4130 472
rect 4190 468 4194 472
rect 4206 468 4210 472
rect 4222 468 4226 472
rect 4302 468 4306 472
rect 4358 468 4362 472
rect 4382 468 4386 472
rect 4438 468 4442 472
rect 4446 468 4450 472
rect 4518 468 4522 472
rect 4534 468 4538 472
rect 4598 468 4602 472
rect 4662 468 4666 472
rect 4678 468 4682 472
rect 4710 468 4714 472
rect 4766 468 4770 472
rect 4782 468 4786 472
rect 4806 468 4810 472
rect 4854 468 4858 472
rect 4886 468 4890 472
rect 4910 468 4914 472
rect 4998 468 5002 472
rect 5046 468 5050 472
rect 5054 468 5058 472
rect 5094 468 5098 472
rect 5118 468 5122 472
rect 5174 468 5178 472
rect 22 458 26 462
rect 54 458 58 462
rect 214 458 218 462
rect 222 458 226 462
rect 270 458 274 462
rect 310 458 314 462
rect 406 458 410 462
rect 446 458 450 462
rect 550 458 554 462
rect 630 458 634 462
rect 646 458 650 462
rect 686 458 690 462
rect 718 458 722 462
rect 734 458 738 462
rect 742 458 746 462
rect 774 458 778 462
rect 806 458 810 462
rect 838 458 842 462
rect 862 458 866 462
rect 902 458 906 462
rect 958 458 962 462
rect 1046 458 1050 462
rect 1070 458 1074 462
rect 1142 458 1146 462
rect 1174 459 1178 463
rect 1222 458 1226 462
rect 1454 459 1458 463
rect 1542 458 1546 462
rect 1654 458 1658 462
rect 1694 458 1698 462
rect 1710 458 1714 462
rect 1726 458 1730 462
rect 1846 458 1850 462
rect 1886 458 1890 462
rect 1974 458 1978 462
rect 1982 458 1986 462
rect 2006 458 2010 462
rect 2182 458 2186 462
rect 2422 458 2426 462
rect 2462 459 2466 463
rect 2558 459 2562 463
rect 2686 458 2690 462
rect 2694 458 2698 462
rect 2726 458 2730 462
rect 2758 458 2762 462
rect 2806 458 2810 462
rect 2822 458 2826 462
rect 2830 458 2834 462
rect 2870 458 2874 462
rect 2878 458 2882 462
rect 3022 458 3026 462
rect 3094 458 3098 462
rect 3334 458 3338 462
rect 3446 458 3450 462
rect 3486 458 3490 462
rect 3510 458 3514 462
rect 3534 458 3538 462
rect 3614 458 3618 462
rect 3646 458 3650 462
rect 3670 458 3674 462
rect 3686 458 3690 462
rect 3726 458 3730 462
rect 3790 458 3794 462
rect 3878 458 3882 462
rect 3910 458 3914 462
rect 3974 458 3978 462
rect 4014 458 4018 462
rect 4054 458 4058 462
rect 4070 458 4074 462
rect 4078 458 4082 462
rect 4094 458 4098 462
rect 4134 458 4138 462
rect 4150 458 4154 462
rect 4222 458 4226 462
rect 4246 458 4250 462
rect 4270 458 4274 462
rect 4278 458 4282 462
rect 4454 458 4458 462
rect 4502 458 4506 462
rect 4558 458 4562 462
rect 4582 458 4586 462
rect 4590 458 4594 462
rect 4614 458 4618 462
rect 4646 458 4650 462
rect 4654 458 4658 462
rect 4670 458 4674 462
rect 4686 458 4690 462
rect 4718 458 4722 462
rect 4790 458 4794 462
rect 4862 458 4866 462
rect 4894 458 4898 462
rect 4950 458 4954 462
rect 5006 458 5010 462
rect 5030 458 5034 462
rect 5086 458 5090 462
rect 5142 458 5146 462
rect 5214 458 5218 462
rect 5246 459 5250 463
rect 382 448 386 452
rect 494 448 498 452
rect 630 448 634 452
rect 678 448 682 452
rect 790 448 794 452
rect 822 448 826 452
rect 830 448 834 452
rect 942 448 946 452
rect 950 448 954 452
rect 1222 448 1226 452
rect 1246 448 1250 452
rect 1294 448 1298 452
rect 1542 448 1546 452
rect 1702 448 1706 452
rect 1798 448 1802 452
rect 1854 448 1858 452
rect 1886 448 1890 452
rect 1894 448 1898 452
rect 1990 448 1994 452
rect 2030 448 2034 452
rect 2838 448 2842 452
rect 2862 448 2866 452
rect 3470 448 3474 452
rect 3526 448 3530 452
rect 3534 448 3538 452
rect 3574 448 3578 452
rect 3590 448 3594 452
rect 3630 448 3634 452
rect 3694 448 3698 452
rect 3854 448 3858 452
rect 3910 448 3914 452
rect 3934 448 3938 452
rect 3958 448 3962 452
rect 4062 448 4066 452
rect 4078 448 4082 452
rect 4142 448 4146 452
rect 4206 448 4210 452
rect 4374 448 4378 452
rect 4518 448 4522 452
rect 4566 448 4570 452
rect 4574 448 4578 452
rect 4606 448 4610 452
rect 4638 448 4642 452
rect 4742 448 4746 452
rect 4958 448 4962 452
rect 5038 448 5042 452
rect 5062 448 5066 452
rect 5070 448 5074 452
rect 5126 448 5130 452
rect 5174 448 5178 452
rect 622 438 626 442
rect 638 438 642 442
rect 686 438 690 442
rect 846 438 850 442
rect 910 438 914 442
rect 966 438 970 442
rect 1014 438 1018 442
rect 1702 438 1706 442
rect 1838 438 1842 442
rect 1950 438 1954 442
rect 1966 438 1970 442
rect 2142 438 2146 442
rect 2886 438 2890 442
rect 2934 438 2938 442
rect 2982 438 2986 442
rect 3134 438 3138 442
rect 3510 438 3514 442
rect 3614 438 3618 442
rect 3710 438 3714 442
rect 3870 438 3874 442
rect 3974 438 3978 442
rect 4150 438 4154 442
rect 4158 438 4162 442
rect 4174 438 4178 442
rect 4494 438 4498 442
rect 4550 438 4554 442
rect 4622 438 4626 442
rect 4718 438 4722 442
rect 4758 438 4762 442
rect 4926 438 4930 442
rect 4942 438 4946 442
rect 5022 438 5026 442
rect 5150 438 5154 442
rect 4934 428 4938 432
rect 5046 428 5050 432
rect 902 418 906 422
rect 982 418 986 422
rect 1110 418 1114 422
rect 1678 418 1682 422
rect 1830 418 1834 422
rect 1958 418 1962 422
rect 2254 418 2258 422
rect 2654 418 2658 422
rect 2878 418 2882 422
rect 2966 418 2970 422
rect 3262 418 3266 422
rect 3606 418 3610 422
rect 3646 418 3650 422
rect 3822 418 3826 422
rect 4326 418 4330 422
rect 4406 418 4410 422
rect 4478 418 4482 422
rect 4502 418 4506 422
rect 4558 418 4562 422
rect 4614 418 4618 422
rect 4702 418 4706 422
rect 4870 418 4874 422
rect 4966 418 4970 422
rect 5014 418 5018 422
rect 5142 418 5146 422
rect 5286 418 5290 422
rect 346 403 350 407
rect 353 403 357 407
rect 1370 403 1374 407
rect 1377 403 1381 407
rect 2394 403 2398 407
rect 2401 403 2405 407
rect 3418 403 3422 407
rect 3425 403 3429 407
rect 4442 403 4446 407
rect 4449 403 4453 407
rect 4910 398 4914 402
rect 174 388 178 392
rect 606 388 610 392
rect 654 388 658 392
rect 686 388 690 392
rect 950 388 954 392
rect 1022 388 1026 392
rect 1174 388 1178 392
rect 1214 388 1218 392
rect 1406 388 1410 392
rect 1462 388 1466 392
rect 1702 388 1706 392
rect 1822 388 1826 392
rect 1894 388 1898 392
rect 1918 388 1922 392
rect 1974 388 1978 392
rect 2542 388 2546 392
rect 2574 388 2578 392
rect 2598 388 2602 392
rect 2662 388 2666 392
rect 2694 388 2698 392
rect 2766 388 2770 392
rect 2806 388 2810 392
rect 2854 388 2858 392
rect 3510 388 3514 392
rect 3790 388 3794 392
rect 4390 388 4394 392
rect 4750 388 4754 392
rect 5054 388 5058 392
rect 5150 388 5154 392
rect 5310 388 5314 392
rect 1502 378 1506 382
rect 2438 378 2442 382
rect 3886 378 3890 382
rect 4430 378 4434 382
rect 342 368 346 372
rect 398 368 402 372
rect 566 368 570 372
rect 598 368 602 372
rect 1550 368 1554 372
rect 1742 368 1746 372
rect 1846 368 1850 372
rect 1926 368 1930 372
rect 1966 368 1970 372
rect 2086 368 2090 372
rect 2182 368 2186 372
rect 2238 368 2242 372
rect 2270 368 2274 372
rect 2654 368 2658 372
rect 2678 368 2682 372
rect 2726 368 2730 372
rect 2742 368 2746 372
rect 2750 368 2754 372
rect 2814 368 2818 372
rect 2830 368 2834 372
rect 3646 368 3650 372
rect 3798 368 3802 372
rect 3822 368 3826 372
rect 3902 368 3906 372
rect 4086 368 4090 372
rect 4174 368 4178 372
rect 4262 368 4266 372
rect 4318 368 4322 372
rect 4494 368 4498 372
rect 4678 368 4682 372
rect 4894 368 4898 372
rect 4910 368 4914 372
rect 4942 368 4946 372
rect 5046 368 5050 372
rect 214 358 218 362
rect 582 358 586 362
rect 670 358 674 362
rect 774 358 778 362
rect 1270 358 1274 362
rect 1510 358 1514 362
rect 1518 358 1522 362
rect 1574 358 1578 362
rect 1582 358 1586 362
rect 1726 358 1730 362
rect 1830 358 1834 362
rect 1862 358 1866 362
rect 1910 358 1914 362
rect 1950 358 1954 362
rect 2102 358 2106 362
rect 2182 358 2186 362
rect 2222 358 2226 362
rect 2558 358 2562 362
rect 2630 358 2634 362
rect 2638 358 2642 362
rect 2670 358 2674 362
rect 2758 358 2762 362
rect 2798 358 2802 362
rect 2830 358 2834 362
rect 3430 358 3434 362
rect 3558 358 3562 362
rect 3582 358 3586 362
rect 3630 358 3634 362
rect 3782 358 3786 362
rect 3846 358 3850 362
rect 3870 358 3874 362
rect 3926 358 3930 362
rect 4006 358 4010 362
rect 4478 358 4482 362
rect 4510 358 4514 362
rect 4542 358 4546 362
rect 4582 358 4586 362
rect 4614 358 4618 362
rect 4806 358 4810 362
rect 4862 358 4866 362
rect 4926 358 4930 362
rect 4958 358 4962 362
rect 5030 358 5034 362
rect 22 348 26 352
rect 62 348 66 352
rect 246 348 250 352
rect 254 348 258 352
rect 502 347 506 351
rect 606 348 610 352
rect 654 348 658 352
rect 686 348 690 352
rect 702 348 706 352
rect 710 348 714 352
rect 726 348 730 352
rect 830 348 834 352
rect 838 348 842 352
rect 854 348 858 352
rect 886 348 890 352
rect 926 348 930 352
rect 1078 348 1082 352
rect 1102 348 1106 352
rect 1294 348 1298 352
rect 1366 348 1370 352
rect 1430 348 1434 352
rect 1526 348 1530 352
rect 1542 348 1546 352
rect 1566 348 1570 352
rect 1678 348 1682 352
rect 1702 348 1706 352
rect 1750 348 1754 352
rect 1758 348 1762 352
rect 1782 348 1786 352
rect 1790 348 1794 352
rect 1846 348 1850 352
rect 1894 348 1898 352
rect 1934 348 1938 352
rect 1958 348 1962 352
rect 2038 348 2042 352
rect 2086 348 2090 352
rect 2110 348 2114 352
rect 2214 348 2218 352
rect 2230 348 2234 352
rect 2302 348 2306 352
rect 2366 348 2370 352
rect 2406 348 2410 352
rect 2486 348 2490 352
rect 2534 348 2538 352
rect 2542 348 2546 352
rect 2574 348 2578 352
rect 2646 348 2650 352
rect 2678 348 2682 352
rect 2686 348 2690 352
rect 2750 348 2754 352
rect 2790 348 2794 352
rect 2806 348 2810 352
rect 2838 348 2842 352
rect 2934 348 2938 352
rect 38 338 42 342
rect 134 338 138 342
rect 142 338 146 342
rect 190 338 194 342
rect 198 338 202 342
rect 238 338 242 342
rect 294 340 298 344
rect 302 338 306 342
rect 310 338 314 342
rect 358 338 362 342
rect 430 338 434 342
rect 518 338 522 342
rect 542 338 546 342
rect 566 338 570 342
rect 582 338 586 342
rect 662 338 666 342
rect 694 338 698 342
rect 742 340 746 344
rect 750 338 754 342
rect 758 338 762 342
rect 798 338 802 342
rect 862 338 866 342
rect 934 338 938 342
rect 982 338 986 342
rect 990 338 994 342
rect 1038 338 1042 342
rect 1142 338 1146 342
rect 1190 338 1194 342
rect 1198 338 1202 342
rect 1254 338 1258 342
rect 1318 338 1322 342
rect 1342 338 1346 342
rect 1358 338 1362 342
rect 1430 338 1434 342
rect 1486 338 1490 342
rect 1494 338 1498 342
rect 1542 338 1546 342
rect 1582 338 1586 342
rect 1598 338 1602 342
rect 1622 338 1626 342
rect 1654 338 1658 342
rect 1662 338 1666 342
rect 1678 338 1682 342
rect 1750 338 1754 342
rect 1814 338 1818 342
rect 1830 338 1834 342
rect 1838 338 1842 342
rect 1886 338 1890 342
rect 2062 338 2066 342
rect 2078 338 2082 342
rect 2118 338 2122 342
rect 2206 338 2210 342
rect 2230 338 2234 342
rect 2334 338 2338 342
rect 2350 338 2354 342
rect 2398 338 2402 342
rect 2998 347 3002 351
rect 3086 348 3090 352
rect 3182 347 3186 351
rect 3326 348 3330 352
rect 3398 348 3402 352
rect 3462 348 3466 352
rect 3486 348 3490 352
rect 3502 348 3506 352
rect 3550 348 3554 352
rect 3646 348 3650 352
rect 3790 348 3794 352
rect 3830 348 3834 352
rect 3870 348 3874 352
rect 3910 348 3914 352
rect 3974 348 3978 352
rect 4022 348 4026 352
rect 4054 348 4058 352
rect 4062 348 4066 352
rect 4078 348 4082 352
rect 4246 348 4250 352
rect 4486 348 4490 352
rect 4510 348 4514 352
rect 4526 348 4530 352
rect 4542 348 4546 352
rect 4598 348 4602 352
rect 4638 348 4642 352
rect 2470 338 2474 342
rect 2478 338 2482 342
rect 2510 338 2514 342
rect 2534 338 2538 342
rect 2566 338 2570 342
rect 2614 338 2618 342
rect 2630 338 2634 342
rect 2710 338 2714 342
rect 2782 338 2786 342
rect 2982 338 2986 342
rect 3094 338 3098 342
rect 3102 338 3106 342
rect 3150 338 3154 342
rect 3166 338 3170 342
rect 3254 338 3258 342
rect 3302 338 3306 342
rect 3334 338 3338 342
rect 3342 338 3346 342
rect 3390 338 3394 342
rect 3454 338 3458 342
rect 3542 338 3546 342
rect 3614 338 3618 342
rect 3670 338 3674 342
rect 3718 338 3722 342
rect 3726 338 3730 342
rect 3774 338 3778 342
rect 3814 338 3818 342
rect 3862 338 3866 342
rect 3982 338 3986 342
rect 3998 338 4002 342
rect 4030 338 4034 342
rect 4086 338 4090 342
rect 4110 338 4114 342
rect 4166 338 4170 342
rect 4214 338 4218 342
rect 4222 338 4226 342
rect 4270 338 4274 342
rect 4278 338 4282 342
rect 4326 338 4330 342
rect 4334 338 4338 342
rect 4382 338 4386 342
rect 4398 338 4402 342
rect 4406 338 4410 342
rect 4454 338 4458 342
rect 4534 338 4538 342
rect 4686 348 4690 352
rect 4694 348 4698 352
rect 4790 348 4794 352
rect 4902 348 4906 352
rect 4918 348 4922 352
rect 4934 348 4938 352
rect 4950 348 4954 352
rect 4974 348 4978 352
rect 5014 348 5018 352
rect 5054 348 5058 352
rect 5102 348 5106 352
rect 5118 348 5122 352
rect 5126 348 5130 352
rect 5214 348 5218 352
rect 5230 348 5234 352
rect 5270 348 5274 352
rect 4558 338 4562 342
rect 4566 338 4570 342
rect 4662 338 4666 342
rect 4686 338 4690 342
rect 4726 338 4730 342
rect 4774 338 4778 342
rect 4782 338 4786 342
rect 4798 338 4802 342
rect 4830 340 4834 344
rect 4838 338 4842 342
rect 4846 338 4850 342
rect 4878 338 4882 342
rect 4990 338 4994 342
rect 5014 338 5018 342
rect 5110 338 5114 342
rect 5142 338 5146 342
rect 5174 338 5178 342
rect 5270 338 5274 342
rect 14 327 18 331
rect 222 328 226 332
rect 270 328 274 332
rect 534 328 538 332
rect 630 328 634 332
rect 718 328 722 332
rect 814 328 818 332
rect 1278 328 1282 332
rect 1334 328 1338 332
rect 1342 328 1346 332
rect 1382 328 1386 332
rect 1414 328 1418 332
rect 1606 328 1610 332
rect 1638 328 1642 332
rect 1694 328 1698 332
rect 1718 328 1722 332
rect 1758 328 1762 332
rect 1806 328 1810 332
rect 2126 328 2130 332
rect 2190 328 2194 332
rect 2510 328 2514 332
rect 2518 328 2522 332
rect 2606 328 2610 332
rect 2702 328 2706 332
rect 2766 328 2770 332
rect 3406 327 3410 331
rect 3462 328 3466 332
rect 3478 328 3482 332
rect 3526 328 3530 332
rect 3566 328 3570 332
rect 3606 328 3610 332
rect 3990 328 3994 332
rect 4038 328 4042 332
rect 4102 328 4106 332
rect 4510 328 4514 332
rect 4574 328 4578 332
rect 4622 328 4626 332
rect 4670 328 4674 332
rect 4718 328 4722 332
rect 4870 328 4874 332
rect 5006 328 5010 332
rect 5078 328 5082 332
rect 5134 328 5138 332
rect 5294 328 5298 332
rect 230 318 234 322
rect 262 318 266 322
rect 278 318 282 322
rect 438 318 442 322
rect 766 318 770 322
rect 782 318 786 322
rect 822 318 826 322
rect 1046 318 1050 322
rect 1614 318 1618 322
rect 1982 318 1986 322
rect 2126 318 2130 322
rect 2254 318 2258 322
rect 2462 318 2466 322
rect 2870 318 2874 322
rect 3062 318 3066 322
rect 3070 318 3074 322
rect 3126 318 3130 322
rect 3246 318 3250 322
rect 3262 318 3266 322
rect 3270 318 3274 322
rect 3310 318 3314 322
rect 3358 318 3362 322
rect 3438 318 3442 322
rect 3534 318 3538 322
rect 3646 318 3650 322
rect 3686 318 3690 322
rect 3742 318 3746 322
rect 3846 318 3850 322
rect 3982 318 3986 322
rect 4134 318 4138 322
rect 4182 318 4186 322
rect 4230 318 4234 322
rect 4294 318 4298 322
rect 4358 318 4362 322
rect 4614 318 4618 322
rect 4710 318 4714 322
rect 4814 318 4818 322
rect 4862 318 4866 322
rect 4998 318 5002 322
rect 5014 318 5018 322
rect 5086 318 5090 322
rect 5118 318 5122 322
rect 270 308 274 312
rect 1534 308 1538 312
rect 1950 308 1954 312
rect 1990 308 1994 312
rect 2430 308 2434 312
rect 2510 308 2514 312
rect 2614 308 2618 312
rect 2702 308 2706 312
rect 3782 308 3786 312
rect 3838 308 3842 312
rect 4038 308 4042 312
rect 4870 308 4874 312
rect 5134 308 5138 312
rect 858 303 862 307
rect 865 303 869 307
rect 1874 303 1878 307
rect 1881 303 1885 307
rect 2906 303 2910 307
rect 2913 303 2917 307
rect 3930 303 3934 307
rect 3937 303 3941 307
rect 4954 303 4958 307
rect 4961 303 4965 307
rect 294 298 298 302
rect 406 298 410 302
rect 422 298 426 302
rect 1782 298 1786 302
rect 1958 298 1962 302
rect 2062 298 2066 302
rect 2478 298 2482 302
rect 2862 298 2866 302
rect 3046 298 3050 302
rect 3150 298 3154 302
rect 4086 298 4090 302
rect 4182 298 4186 302
rect 4878 298 4882 302
rect 78 288 82 292
rect 446 288 450 292
rect 598 288 602 292
rect 870 288 874 292
rect 878 288 882 292
rect 982 288 986 292
rect 1102 288 1106 292
rect 1174 288 1178 292
rect 1198 288 1202 292
rect 1254 288 1258 292
rect 1302 288 1306 292
rect 1422 288 1426 292
rect 1438 288 1442 292
rect 1470 288 1474 292
rect 1518 288 1522 292
rect 1622 288 1626 292
rect 1734 288 1738 292
rect 1822 288 1826 292
rect 2014 288 2018 292
rect 2022 288 2026 292
rect 2038 288 2042 292
rect 2054 288 2058 292
rect 2214 288 2218 292
rect 2310 288 2314 292
rect 2422 288 2426 292
rect 2454 288 2458 292
rect 2526 288 2530 292
rect 2574 288 2578 292
rect 2662 288 2666 292
rect 2670 288 2674 292
rect 2734 288 2738 292
rect 2742 288 2746 292
rect 2814 288 2818 292
rect 3094 288 3098 292
rect 3118 288 3122 292
rect 3542 288 3546 292
rect 3726 288 3730 292
rect 3766 288 3770 292
rect 4006 288 4010 292
rect 4102 288 4106 292
rect 4134 288 4138 292
rect 4206 288 4210 292
rect 4246 288 4250 292
rect 4342 288 4346 292
rect 4798 288 4802 292
rect 4886 288 4890 292
rect 4990 288 4994 292
rect 5030 288 5034 292
rect 5182 288 5186 292
rect 5190 288 5194 292
rect 5294 288 5298 292
rect 238 278 242 282
rect 286 278 290 282
rect 318 278 322 282
rect 422 278 426 282
rect 726 278 730 282
rect 766 278 770 282
rect 1014 278 1018 282
rect 1078 278 1082 282
rect 1206 278 1210 282
rect 1382 278 1386 282
rect 1430 278 1434 282
rect 1598 278 1602 282
rect 1630 278 1634 282
rect 1742 278 1746 282
rect 1782 278 1786 282
rect 1870 279 1874 283
rect 1958 278 1962 282
rect 2062 278 2066 282
rect 2342 278 2346 282
rect 2478 278 2482 282
rect 2534 278 2538 282
rect 2582 278 2586 282
rect 2590 278 2594 282
rect 2782 278 2786 282
rect 2862 278 2866 282
rect 2870 278 2874 282
rect 3046 278 3050 282
rect 3070 278 3074 282
rect 3150 278 3154 282
rect 3246 278 3250 282
rect 3294 278 3298 282
rect 3486 278 3490 282
rect 3518 278 3522 282
rect 3582 278 3586 282
rect 3662 278 3666 282
rect 3774 278 3778 282
rect 4182 278 4186 282
rect 4294 278 4298 282
rect 4398 278 4402 282
rect 4574 279 4578 283
rect 4838 278 4842 282
rect 4870 278 4874 282
rect 4878 278 4882 282
rect 4958 278 4962 282
rect 4982 278 4986 282
rect 5134 278 5138 282
rect 5262 279 5266 283
rect 62 268 66 272
rect 222 268 226 272
rect 270 268 274 272
rect 294 268 298 272
rect 358 268 362 272
rect 414 268 418 272
rect 422 268 426 272
rect 478 268 482 272
rect 518 268 522 272
rect 582 268 586 272
rect 630 268 634 272
rect 710 268 714 272
rect 806 268 810 272
rect 862 268 866 272
rect 910 268 914 272
rect 22 258 26 262
rect 46 258 50 262
rect 102 258 106 262
rect 126 258 130 262
rect 166 258 170 262
rect 214 258 218 262
rect 230 258 234 262
rect 262 258 266 262
rect 270 258 274 262
rect 294 258 298 262
rect 342 258 346 262
rect 374 258 378 262
rect 526 258 530 262
rect 654 258 658 262
rect 686 258 690 262
rect 702 258 706 262
rect 750 258 754 262
rect 822 258 826 262
rect 926 258 930 262
rect 950 258 954 262
rect 966 258 970 262
rect 1014 268 1018 272
rect 1038 268 1042 272
rect 1086 268 1090 272
rect 1134 268 1138 272
rect 1142 268 1146 272
rect 1190 268 1194 272
rect 1238 268 1242 272
rect 1278 268 1282 272
rect 1310 268 1314 272
rect 1318 268 1322 272
rect 1326 268 1330 272
rect 1350 268 1354 272
rect 1358 268 1362 272
rect 1398 268 1402 272
rect 1446 268 1450 272
rect 1478 268 1482 272
rect 1486 268 1490 272
rect 1534 268 1538 272
rect 1550 268 1554 272
rect 1582 268 1586 272
rect 1598 268 1602 272
rect 1678 268 1682 272
rect 1710 268 1714 272
rect 1726 268 1730 272
rect 1742 268 1746 272
rect 1774 268 1778 272
rect 1822 268 1826 272
rect 1854 268 1858 272
rect 1902 268 1906 272
rect 1950 268 1954 272
rect 1958 268 1962 272
rect 1982 268 1986 272
rect 1990 268 1994 272
rect 2022 268 2026 272
rect 2118 268 2122 272
rect 2230 268 2234 272
rect 2430 268 2434 272
rect 2486 268 2490 272
rect 2526 268 2530 272
rect 2550 268 2554 272
rect 2646 268 2650 272
rect 2654 268 2658 272
rect 2702 268 2706 272
rect 2726 268 2730 272
rect 2742 268 2746 272
rect 2798 268 2802 272
rect 2814 268 2818 272
rect 2830 268 2834 272
rect 2854 268 2858 272
rect 2974 268 2978 272
rect 3006 268 3010 272
rect 3038 268 3042 272
rect 3086 268 3090 272
rect 3118 268 3122 272
rect 3142 268 3146 272
rect 3150 268 3154 272
rect 3206 268 3210 272
rect 3254 268 3258 272
rect 3294 268 3298 272
rect 3318 268 3322 272
rect 3470 268 3474 272
rect 3494 268 3498 272
rect 3510 268 3514 272
rect 3526 268 3530 272
rect 3574 268 3578 272
rect 3598 268 3602 272
rect 3630 268 3634 272
rect 3646 268 3650 272
rect 3670 268 3674 272
rect 3718 268 3722 272
rect 3758 268 3762 272
rect 3782 268 3786 272
rect 3830 268 3834 272
rect 3838 268 3842 272
rect 3886 268 3890 272
rect 3998 268 4002 272
rect 4102 268 4106 272
rect 4174 268 4178 272
rect 4182 268 4186 272
rect 4246 268 4250 272
rect 4302 268 4306 272
rect 4374 268 4378 272
rect 4462 268 4466 272
rect 4494 268 4498 272
rect 4590 268 4594 272
rect 4638 268 4642 272
rect 4646 268 4650 272
rect 4702 268 4706 272
rect 4750 268 4754 272
rect 4758 268 4762 272
rect 4790 268 4794 272
rect 4894 268 4898 272
rect 4910 268 4914 272
rect 4926 268 4930 272
rect 4950 268 4954 272
rect 4998 268 5002 272
rect 5062 268 5066 272
rect 5102 268 5106 272
rect 5126 268 5130 272
rect 5158 268 5162 272
rect 5166 268 5170 272
rect 5214 268 5218 272
rect 998 258 1002 262
rect 1022 258 1026 262
rect 1030 258 1034 262
rect 1046 258 1050 262
rect 1054 258 1058 262
rect 1086 258 1090 262
rect 1238 258 1242 262
rect 1262 258 1266 262
rect 1286 258 1290 262
rect 1406 258 1410 262
rect 1454 258 1458 262
rect 1558 258 1562 262
rect 1574 258 1578 262
rect 1606 258 1610 262
rect 1654 258 1658 262
rect 1686 258 1690 262
rect 1702 258 1706 262
rect 1718 258 1722 262
rect 1766 258 1770 262
rect 1822 258 1826 262
rect 1830 258 1834 262
rect 1846 258 1850 262
rect 1878 258 1882 262
rect 1950 258 1954 262
rect 1998 258 2002 262
rect 2046 258 2050 262
rect 2150 259 2154 263
rect 2182 258 2186 262
rect 2254 258 2258 262
rect 2270 258 2274 262
rect 2350 258 2354 262
rect 2438 258 2442 262
rect 2462 258 2466 262
rect 2518 258 2522 262
rect 2766 258 2770 262
rect 2806 258 2810 262
rect 5238 266 5242 270
rect 5246 268 5250 272
rect 2902 258 2906 262
rect 2950 258 2954 262
rect 2998 258 3002 262
rect 3030 258 3034 262
rect 3062 258 3066 262
rect 3078 258 3082 262
rect 3094 258 3098 262
rect 3158 258 3162 262
rect 3230 258 3234 262
rect 3262 258 3266 262
rect 3310 258 3314 262
rect 3318 258 3322 262
rect 3358 258 3362 262
rect 3390 258 3394 262
rect 3438 258 3442 262
rect 3462 258 3466 262
rect 54 248 58 252
rect 78 248 82 252
rect 110 248 114 252
rect 118 248 122 252
rect 150 248 154 252
rect 246 248 250 252
rect 310 248 314 252
rect 350 248 354 252
rect 662 248 666 252
rect 694 248 698 252
rect 798 248 802 252
rect 838 248 842 252
rect 918 248 922 252
rect 950 248 954 252
rect 1270 248 1274 252
rect 1302 248 1306 252
rect 1326 248 1330 252
rect 1398 248 1402 252
rect 1462 248 1466 252
rect 1566 248 1570 252
rect 1750 248 1754 252
rect 1806 248 1810 252
rect 2038 248 2042 252
rect 2726 248 2730 252
rect 2774 248 2778 252
rect 2830 248 2834 252
rect 2910 248 2914 252
rect 3014 248 3018 252
rect 3102 248 3106 252
rect 3118 248 3122 252
rect 3238 248 3242 252
rect 3326 248 3330 252
rect 3342 248 3346 252
rect 3350 248 3354 252
rect 3382 248 3386 252
rect 3430 248 3434 252
rect 3622 248 3626 252
rect 3646 258 3650 262
rect 3750 258 3754 262
rect 3814 258 3818 262
rect 3862 258 3866 262
rect 3910 258 3914 262
rect 3942 258 3946 262
rect 4038 258 4042 262
rect 4054 258 4058 262
rect 4102 258 4106 262
rect 4134 258 4138 262
rect 4326 258 4330 262
rect 4430 258 4434 262
rect 4550 258 4554 262
rect 4582 258 4586 262
rect 4662 258 4666 262
rect 4686 258 4690 262
rect 4710 258 4714 262
rect 4718 258 4722 262
rect 4726 258 4730 262
rect 4766 258 4770 262
rect 4806 258 4810 262
rect 4830 258 4834 262
rect 4902 258 4906 262
rect 5006 258 5010 262
rect 5030 258 5034 262
rect 5046 258 5050 262
rect 5078 258 5082 262
rect 5102 258 5106 262
rect 5118 258 5122 262
rect 5150 258 5154 262
rect 5182 258 5186 262
rect 5206 258 5210 262
rect 5222 258 5226 262
rect 5270 258 5274 262
rect 5286 258 5290 262
rect 5294 258 5298 262
rect 3726 248 3730 252
rect 4118 248 4122 252
rect 4134 248 4138 252
rect 4246 248 4250 252
rect 4270 248 4274 252
rect 4662 248 4666 252
rect 4694 248 4698 252
rect 4726 248 4730 252
rect 4734 248 4738 252
rect 4782 248 4786 252
rect 4830 248 4834 252
rect 4910 248 4914 252
rect 5038 248 5042 252
rect 5046 248 5050 252
rect 5078 248 5082 252
rect 5102 248 5106 252
rect 5134 248 5138 252
rect 5302 248 5306 252
rect 38 238 42 242
rect 118 238 122 242
rect 134 238 138 242
rect 358 238 362 242
rect 382 238 386 242
rect 398 238 402 242
rect 646 238 650 242
rect 654 238 658 242
rect 678 238 682 242
rect 742 238 746 242
rect 934 238 938 242
rect 1230 238 1234 242
rect 1254 238 1258 242
rect 1550 238 1554 242
rect 1646 238 1650 242
rect 2294 238 2298 242
rect 2758 238 2762 242
rect 2894 238 2898 242
rect 2942 238 2946 242
rect 3222 238 3226 242
rect 3310 238 3314 242
rect 3366 238 3370 242
rect 3398 238 3402 242
rect 3446 238 3450 242
rect 4142 238 4146 242
rect 4158 238 4162 242
rect 4398 238 4402 242
rect 4614 238 4618 242
rect 4678 238 4682 242
rect 4854 238 4858 242
rect 4926 238 4930 242
rect 5022 238 5026 242
rect 5030 238 5034 242
rect 5086 238 5090 242
rect 5286 238 5290 242
rect 1654 228 1658 232
rect 3390 228 3394 232
rect 3438 228 3442 232
rect 5014 228 5018 232
rect 46 218 50 222
rect 86 218 90 222
rect 142 218 146 222
rect 166 218 170 222
rect 190 218 194 222
rect 318 218 322 222
rect 390 218 394 222
rect 574 218 578 222
rect 654 218 658 222
rect 726 218 730 222
rect 750 218 754 222
rect 822 218 826 222
rect 926 218 930 222
rect 1598 218 1602 222
rect 2086 218 2090 222
rect 2630 218 2634 222
rect 2710 218 2714 222
rect 2750 218 2754 222
rect 2782 218 2786 222
rect 2878 218 2882 222
rect 2902 218 2906 222
rect 2950 218 2954 222
rect 2998 218 3002 222
rect 3030 218 3034 222
rect 3230 218 3234 222
rect 3278 218 3282 222
rect 3358 218 3362 222
rect 3486 218 3490 222
rect 3686 218 3690 222
rect 4686 218 4690 222
rect 4766 218 4770 222
rect 4462 208 4466 212
rect 4542 208 4546 212
rect 4598 208 4602 212
rect 346 203 350 207
rect 353 203 357 207
rect 1370 203 1374 207
rect 1377 203 1381 207
rect 2394 203 2398 207
rect 2401 203 2405 207
rect 3418 203 3422 207
rect 3425 203 3429 207
rect 4442 203 4446 207
rect 4449 203 4453 207
rect 102 188 106 192
rect 150 188 154 192
rect 214 188 218 192
rect 270 188 274 192
rect 622 188 626 192
rect 726 188 730 192
rect 1094 188 1098 192
rect 1126 188 1130 192
rect 1150 188 1154 192
rect 1398 188 1402 192
rect 1478 188 1482 192
rect 1526 188 1530 192
rect 1582 188 1586 192
rect 1654 188 1658 192
rect 1678 188 1682 192
rect 1710 188 1714 192
rect 1774 188 1778 192
rect 1830 188 1834 192
rect 1926 188 1930 192
rect 1974 188 1978 192
rect 2078 188 2082 192
rect 2350 188 2354 192
rect 2614 188 2618 192
rect 3758 188 3762 192
rect 3782 188 3786 192
rect 4166 188 4170 192
rect 4342 188 4346 192
rect 4502 188 4506 192
rect 5070 188 5074 192
rect 5102 188 5106 192
rect 5134 188 5138 192
rect 1622 178 1626 182
rect 3950 178 3954 182
rect 4878 178 4882 182
rect 78 168 82 172
rect 94 168 98 172
rect 454 168 458 172
rect 542 168 546 172
rect 574 168 578 172
rect 638 168 642 172
rect 814 168 818 172
rect 1038 168 1042 172
rect 1102 168 1106 172
rect 1134 168 1138 172
rect 1534 168 1538 172
rect 1542 168 1546 172
rect 1598 168 1602 172
rect 1630 168 1634 172
rect 1662 168 1666 172
rect 1686 168 1690 172
rect 1718 168 1722 172
rect 1870 168 1874 172
rect 2558 168 2562 172
rect 2742 168 2746 172
rect 2862 168 2866 172
rect 3190 168 3194 172
rect 3574 168 3578 172
rect 3638 168 3642 172
rect 3742 168 3746 172
rect 3790 168 3794 172
rect 3814 168 3818 172
rect 4422 168 4426 172
rect 4702 168 4706 172
rect 4758 168 4762 172
rect 4854 168 4858 172
rect 5062 168 5066 172
rect 5078 168 5082 172
rect 5110 168 5114 172
rect 5294 168 5298 172
rect 230 158 234 162
rect 6 148 10 152
rect 30 148 34 152
rect 94 148 98 152
rect 118 148 122 152
rect 182 148 186 152
rect 334 158 338 162
rect 438 158 442 162
rect 558 158 562 162
rect 566 158 570 162
rect 590 158 594 162
rect 646 158 650 162
rect 702 158 706 162
rect 798 158 802 162
rect 830 158 834 162
rect 902 158 906 162
rect 1054 158 1058 162
rect 1078 158 1082 162
rect 1086 158 1090 162
rect 1118 158 1122 162
rect 1174 158 1178 162
rect 1190 158 1194 162
rect 1390 158 1394 162
rect 1446 158 1450 162
rect 1550 158 1554 162
rect 1558 158 1562 162
rect 1606 158 1610 162
rect 1614 158 1618 162
rect 1646 158 1650 162
rect 1702 158 1706 162
rect 1790 158 1794 162
rect 2038 158 2042 162
rect 2118 158 2122 162
rect 2174 158 2178 162
rect 2654 158 2658 162
rect 2734 158 2738 162
rect 366 148 370 152
rect 382 148 386 152
rect 398 148 402 152
rect 406 148 410 152
rect 446 148 450 152
rect 494 148 498 152
rect 526 148 530 152
rect 550 148 554 152
rect 582 148 586 152
rect 598 148 602 152
rect 662 148 666 152
rect 702 148 706 152
rect 806 148 810 152
rect 902 148 906 152
rect 958 148 962 152
rect 1030 148 1034 152
rect 1046 148 1050 152
rect 1094 148 1098 152
rect 1126 148 1130 152
rect 1150 148 1154 152
rect 62 138 66 142
rect 158 138 162 142
rect 166 138 170 142
rect 246 138 250 142
rect 254 138 258 142
rect 310 138 314 142
rect 334 138 338 142
rect 374 138 378 142
rect 486 138 490 142
rect 518 138 522 142
rect 526 138 530 142
rect 606 138 610 142
rect 646 138 650 142
rect 670 138 674 142
rect 710 138 714 142
rect 782 140 786 144
rect 790 138 794 142
rect 846 138 850 142
rect 854 138 858 142
rect 886 138 890 142
rect 918 138 922 142
rect 926 138 930 142
rect 942 138 946 142
rect 1022 138 1026 142
rect 1294 147 1298 151
rect 1326 148 1330 152
rect 1350 148 1354 152
rect 1470 148 1474 152
rect 1518 148 1522 152
rect 1542 148 1546 152
rect 1598 148 1602 152
rect 1622 148 1626 152
rect 1654 148 1658 152
rect 1694 148 1698 152
rect 1726 148 1730 152
rect 1774 148 1778 152
rect 1838 148 1842 152
rect 1862 148 1866 152
rect 2014 148 2018 152
rect 2190 148 2194 152
rect 2270 148 2274 152
rect 2326 148 2330 152
rect 2398 148 2402 152
rect 2678 148 2682 152
rect 2726 148 2730 152
rect 2766 158 2770 162
rect 2798 158 2802 162
rect 2814 158 2818 162
rect 2870 158 2874 162
rect 2966 158 2970 162
rect 3022 158 3026 162
rect 3142 158 3146 162
rect 3278 158 3282 162
rect 3310 158 3314 162
rect 3326 158 3330 162
rect 3366 158 3370 162
rect 3454 158 3458 162
rect 3566 158 3570 162
rect 3590 158 3594 162
rect 3598 158 3602 162
rect 3622 158 3626 162
rect 3654 158 3658 162
rect 3694 158 3698 162
rect 3710 158 3714 162
rect 3774 158 3778 162
rect 3830 158 3834 162
rect 4774 158 4778 162
rect 4806 158 4810 162
rect 4838 158 4842 162
rect 4870 158 4874 162
rect 4918 158 4922 162
rect 4950 158 4954 162
rect 4990 158 4994 162
rect 5094 158 5098 162
rect 5142 158 5146 162
rect 5150 158 5154 162
rect 5270 158 5274 162
rect 2782 148 2786 152
rect 2814 148 2818 152
rect 2846 148 2850 152
rect 2862 148 2866 152
rect 2886 148 2890 152
rect 2926 148 2930 152
rect 2958 148 2962 152
rect 3022 148 3026 152
rect 3078 148 3082 152
rect 3134 148 3138 152
rect 3158 148 3162 152
rect 3174 148 3178 152
rect 3230 148 3234 152
rect 3254 148 3258 152
rect 3302 148 3306 152
rect 3350 148 3354 152
rect 3438 148 3442 152
rect 3486 148 3490 152
rect 3582 148 3586 152
rect 3630 148 3634 152
rect 3654 148 3658 152
rect 3694 148 3698 152
rect 3710 148 3714 152
rect 3734 148 3738 152
rect 3782 148 3786 152
rect 3822 148 3826 152
rect 3886 148 3890 152
rect 1174 138 1178 142
rect 1190 138 1194 142
rect 1214 138 1218 142
rect 1294 138 1298 142
rect 1406 138 1410 142
rect 1414 138 1418 142
rect 1438 138 1442 142
rect 1462 138 1466 142
rect 1510 138 1514 142
rect 1558 138 1562 142
rect 1574 138 1578 142
rect 1742 138 1746 142
rect 1782 138 1786 142
rect 1798 138 1802 142
rect 1814 138 1818 142
rect 1870 138 1874 142
rect 1910 138 1914 142
rect 1942 138 1946 142
rect 1958 138 1962 142
rect 2006 138 2010 142
rect 2054 138 2058 142
rect 2062 138 2066 142
rect 2110 138 2114 142
rect 2134 138 2138 142
rect 2142 138 2146 142
rect 2158 138 2162 142
rect 2174 138 2178 142
rect 2294 138 2298 142
rect 2334 138 2338 142
rect 2382 138 2386 142
rect 2430 138 2434 142
rect 2478 138 2482 142
rect 2486 138 2490 142
rect 2534 138 2538 142
rect 2542 138 2546 142
rect 2590 138 2594 142
rect 2686 138 2690 142
rect 2718 138 2722 142
rect 2742 138 2746 142
rect 2790 138 2794 142
rect 2822 138 2826 142
rect 2894 138 2898 142
rect 2934 138 2938 142
rect 2950 138 2954 142
rect 2982 138 2986 142
rect 3006 138 3010 142
rect 3014 138 3018 142
rect 3046 138 3050 142
rect 3070 138 3074 142
rect 3110 138 3114 142
rect 3222 138 3226 142
rect 3230 138 3234 142
rect 3310 138 3314 142
rect 3326 138 3330 142
rect 3358 138 3362 142
rect 3382 138 3386 142
rect 3406 138 3410 142
rect 3438 138 3442 142
rect 3478 138 3482 142
rect 3526 138 3530 142
rect 3614 138 3618 142
rect 3638 138 3642 142
rect 3902 147 3906 151
rect 3990 148 3994 152
rect 4046 148 4050 152
rect 4094 147 4098 151
rect 4198 148 4202 152
rect 4230 147 4234 151
rect 4334 148 4338 152
rect 3686 138 3690 142
rect 3766 138 3770 142
rect 3918 138 3922 142
rect 14 127 18 131
rect 54 128 58 132
rect 118 128 122 132
rect 126 128 130 132
rect 174 128 178 132
rect 382 128 386 132
rect 430 128 434 132
rect 470 128 474 132
rect 478 128 482 132
rect 502 128 506 132
rect 630 128 634 132
rect 870 128 874 132
rect 926 128 930 132
rect 958 128 962 132
rect 990 128 994 132
rect 1022 128 1026 132
rect 1070 128 1074 132
rect 1166 128 1170 132
rect 1222 128 1226 132
rect 1438 128 1442 132
rect 1494 128 1498 132
rect 1822 128 1826 132
rect 1918 128 1922 132
rect 1950 128 1954 132
rect 2038 128 2042 132
rect 2174 128 2178 132
rect 2702 128 2706 132
rect 2750 128 2754 132
rect 2830 128 2834 132
rect 2838 128 2842 132
rect 2870 128 2874 132
rect 2918 128 2922 132
rect 2990 128 2994 132
rect 3062 128 3066 132
rect 3118 128 3122 132
rect 4102 138 4106 142
rect 4262 138 4266 142
rect 4310 138 4314 142
rect 4358 138 4362 142
rect 4406 138 4410 142
rect 4414 138 4418 142
rect 4462 138 4466 142
rect 4646 148 4650 152
rect 4654 148 4658 152
rect 4678 148 4682 152
rect 4702 148 4706 152
rect 4726 148 4730 152
rect 4782 148 4786 152
rect 4798 148 4802 152
rect 4862 148 4866 152
rect 4894 148 4898 152
rect 5030 148 5034 152
rect 5086 148 5090 152
rect 5118 148 5122 152
rect 5206 148 5210 152
rect 4534 138 4538 142
rect 4542 138 4546 142
rect 4590 138 4594 142
rect 4598 138 4602 142
rect 5238 147 5242 151
rect 4686 138 4690 142
rect 4734 138 4738 142
rect 4790 138 4794 142
rect 4798 138 4802 142
rect 4918 138 4922 142
rect 4934 138 4938 142
rect 4974 138 4978 142
rect 5006 138 5010 142
rect 5046 138 5050 142
rect 5070 138 5074 142
rect 5166 138 5170 142
rect 5286 138 5290 142
rect 3246 128 3250 132
rect 3254 128 3258 132
rect 3374 128 3378 132
rect 3390 128 3394 132
rect 3398 128 3402 132
rect 3462 128 3466 132
rect 3470 128 3474 132
rect 3494 128 3498 132
rect 3526 128 3530 132
rect 3534 128 3538 132
rect 3558 128 3562 132
rect 3718 128 3722 132
rect 3742 128 3746 132
rect 3982 128 3986 132
rect 4014 128 4018 132
rect 4054 127 4058 131
rect 4350 128 4354 132
rect 4702 128 4706 132
rect 4718 128 4722 132
rect 4742 128 4746 132
rect 4758 128 4762 132
rect 4838 128 4842 132
rect 4886 128 4890 132
rect 4982 128 4986 132
rect 4998 128 5002 132
rect 5038 128 5042 132
rect 5142 128 5146 132
rect 5174 128 5178 132
rect 5238 128 5242 132
rect 238 118 242 122
rect 422 118 426 122
rect 462 118 466 122
rect 510 118 514 122
rect 766 118 770 122
rect 822 118 826 122
rect 830 118 834 122
rect 902 118 906 122
rect 966 118 970 122
rect 1230 118 1234 122
rect 1446 118 1450 122
rect 1846 118 1850 122
rect 1998 118 2002 122
rect 2118 118 2122 122
rect 2446 118 2450 122
rect 2502 118 2506 122
rect 2662 118 2666 122
rect 2694 118 2698 122
rect 2974 118 2978 122
rect 2998 118 3002 122
rect 3070 118 3074 122
rect 3454 118 3458 122
rect 3502 118 3506 122
rect 3598 118 3602 122
rect 3822 118 3826 122
rect 4158 118 4162 122
rect 4294 118 4298 122
rect 4374 118 4378 122
rect 4558 118 4562 122
rect 4614 118 4618 122
rect 4766 118 4770 122
rect 5166 118 5170 122
rect 5286 118 5290 122
rect 54 108 58 112
rect 70 108 74 112
rect 1950 108 1954 112
rect 3118 108 3122 112
rect 3958 108 3962 112
rect 5038 108 5042 112
rect 5094 108 5098 112
rect 5126 108 5130 112
rect 5142 108 5146 112
rect 858 103 862 107
rect 865 103 869 107
rect 1874 103 1878 107
rect 1881 103 1885 107
rect 2906 103 2910 107
rect 2913 103 2917 107
rect 3930 103 3934 107
rect 3937 103 3941 107
rect 4954 103 4958 107
rect 4961 103 4965 107
rect 174 98 178 102
rect 518 98 522 102
rect 678 98 682 102
rect 2398 98 2402 102
rect 2734 98 2738 102
rect 2862 98 2866 102
rect 3174 98 3178 102
rect 4654 98 4658 102
rect 4894 98 4898 102
rect 78 88 82 92
rect 94 88 98 92
rect 150 88 154 92
rect 166 88 170 92
rect 454 88 458 92
rect 542 88 546 92
rect 550 88 554 92
rect 558 88 562 92
rect 598 88 602 92
rect 614 88 618 92
rect 702 88 706 92
rect 846 88 850 92
rect 998 88 1002 92
rect 1038 88 1042 92
rect 1086 88 1090 92
rect 1342 88 1346 92
rect 1398 88 1402 92
rect 1462 88 1466 92
rect 1582 88 1586 92
rect 1614 88 1618 92
rect 1702 88 1706 92
rect 1734 88 1738 92
rect 1830 88 1834 92
rect 1854 88 1858 92
rect 2054 88 2058 92
rect 2086 88 2090 92
rect 2334 88 2338 92
rect 2462 88 2466 92
rect 2590 88 2594 92
rect 2614 88 2618 92
rect 2654 88 2658 92
rect 2702 88 2706 92
rect 2750 88 2754 92
rect 2886 88 2890 92
rect 3030 88 3034 92
rect 3230 88 3234 92
rect 3310 88 3314 92
rect 3382 88 3386 92
rect 3774 88 3778 92
rect 3806 88 3810 92
rect 3886 88 3890 92
rect 3942 88 3946 92
rect 3982 88 3986 92
rect 4166 88 4170 92
rect 4262 88 4266 92
rect 4494 88 4498 92
rect 4606 88 4610 92
rect 4838 88 4842 92
rect 4870 88 4874 92
rect 4926 88 4930 92
rect 5022 88 5026 92
rect 5078 88 5082 92
rect 5270 88 5274 92
rect 38 79 42 83
rect 110 79 114 83
rect 174 78 178 82
rect 262 78 266 82
rect 302 78 306 82
rect 438 78 442 82
rect 510 78 514 82
rect 518 78 522 82
rect 662 78 666 82
rect 678 78 682 82
rect 1006 78 1010 82
rect 1022 78 1026 82
rect 78 68 82 72
rect 126 68 130 72
rect 134 66 138 70
rect 174 68 178 72
rect 230 68 234 72
rect 238 68 242 72
rect 270 68 274 72
rect 302 68 306 72
rect 318 68 322 72
rect 366 68 370 72
rect 422 68 426 72
rect 438 68 442 72
rect 470 68 474 72
rect 494 68 498 72
rect 518 68 522 72
rect 526 68 530 72
rect 550 68 554 72
rect 566 68 570 72
rect 606 68 610 72
rect 654 68 658 72
rect 686 68 690 72
rect 750 68 754 72
rect 758 68 762 72
rect 766 68 770 72
rect 790 68 794 72
rect 798 68 802 72
rect 30 58 34 62
rect 70 58 74 62
rect 102 58 106 62
rect 158 58 162 62
rect 182 58 186 62
rect 246 58 250 62
rect 262 58 266 62
rect 390 58 394 62
rect 414 58 418 62
rect 478 58 482 62
rect 486 58 490 62
rect 582 58 586 62
rect 622 58 626 62
rect 662 58 666 62
rect 718 58 722 62
rect 734 58 738 62
rect 806 58 810 62
rect 902 68 906 72
rect 950 68 954 72
rect 990 68 994 72
rect 1006 68 1010 72
rect 1062 78 1066 82
rect 1126 78 1130 82
rect 1166 78 1170 82
rect 1222 78 1226 82
rect 1470 78 1474 82
rect 1502 78 1506 82
rect 1526 78 1530 82
rect 1534 78 1538 82
rect 1678 78 1682 82
rect 1686 78 1690 82
rect 1766 78 1770 82
rect 2078 78 2082 82
rect 2526 78 2530 82
rect 2734 78 2738 82
rect 2798 78 2802 82
rect 2806 78 2810 82
rect 2846 78 2850 82
rect 2862 78 2866 82
rect 2878 78 2882 82
rect 3150 78 3154 82
rect 3174 78 3178 82
rect 3206 78 3210 82
rect 3214 78 3218 82
rect 3294 78 3298 82
rect 3302 78 3306 82
rect 3630 78 3634 82
rect 3646 78 3650 82
rect 3718 78 3722 82
rect 3758 78 3762 82
rect 3766 78 3770 82
rect 3854 78 3858 82
rect 3870 78 3874 82
rect 3910 78 3914 82
rect 1054 68 1058 72
rect 1078 68 1082 72
rect 1118 68 1122 72
rect 1142 68 1146 72
rect 1182 68 1186 72
rect 1222 68 1226 72
rect 1246 68 1250 72
rect 1302 68 1306 72
rect 1310 68 1314 72
rect 1358 68 1362 72
rect 1382 68 1386 72
rect 1430 68 1434 72
rect 1518 68 1522 72
rect 1550 68 1554 72
rect 1630 68 1634 72
rect 1670 68 1674 72
rect 1678 68 1682 72
rect 1726 68 1730 72
rect 1758 68 1762 72
rect 1806 66 1810 70
rect 1814 68 1818 72
rect 1822 68 1826 72
rect 1942 68 1946 72
rect 2038 68 2042 72
rect 2070 68 2074 72
rect 2102 68 2106 72
rect 2366 68 2370 72
rect 2390 68 2394 72
rect 2438 68 2442 72
rect 2446 68 2450 72
rect 2494 68 2498 72
rect 2598 68 2602 72
rect 2646 68 2650 72
rect 2654 68 2658 72
rect 2670 68 2674 72
rect 2726 68 2730 72
rect 2758 68 2762 72
rect 2814 68 2818 72
rect 2838 68 2842 72
rect 3014 68 3018 72
rect 3094 68 3098 72
rect 3158 68 3162 72
rect 3222 68 3226 72
rect 3270 68 3274 72
rect 3286 68 3290 72
rect 3326 68 3330 72
rect 3358 68 3362 72
rect 3366 68 3370 72
rect 3414 68 3418 72
rect 3438 68 3442 72
rect 926 58 930 62
rect 982 58 986 62
rect 1046 58 1050 62
rect 1150 58 1154 62
rect 1166 58 1170 62
rect 1206 58 1210 62
rect 1270 58 1274 62
rect 1438 58 1442 62
rect 1478 58 1482 62
rect 1558 58 1562 62
rect 1582 58 1586 62
rect 1614 58 1618 62
rect 1718 58 1722 62
rect 1750 58 1754 62
rect 1782 58 1786 62
rect 1790 58 1794 62
rect 1918 58 1922 62
rect 2022 59 2026 63
rect 2158 58 2162 62
rect 2190 59 2194 63
rect 2246 59 2250 63
rect 2526 59 2530 63
rect 2678 58 2682 62
rect 2686 58 2690 62
rect 2758 58 2762 62
rect 2782 58 2786 62
rect 2830 58 2834 62
rect 2846 58 2850 62
rect 2894 58 2898 62
rect 2918 58 2922 62
rect 2966 58 2970 62
rect 2990 58 2994 62
rect 3086 58 3090 62
rect 3118 58 3122 62
rect 3134 58 3138 62
rect 3174 58 3178 62
rect 3190 58 3194 62
rect 3222 58 3226 62
rect 3278 58 3282 62
rect 3342 58 3346 62
rect 3430 58 3434 62
rect 3526 68 3530 72
rect 3574 68 3578 72
rect 3614 68 3618 72
rect 3630 68 3634 72
rect 3654 68 3658 72
rect 3702 68 3706 72
rect 3726 68 3730 72
rect 3790 66 3794 70
rect 3798 68 3802 72
rect 3822 68 3826 72
rect 3846 68 3850 72
rect 4318 78 4322 82
rect 4334 78 4338 82
rect 4558 78 4562 82
rect 5070 78 5074 82
rect 5158 78 5162 82
rect 5206 78 5210 82
rect 5238 78 5242 82
rect 3918 68 3922 72
rect 4014 68 4018 72
rect 4118 68 4122 72
rect 4214 68 4218 72
rect 4270 68 4274 72
rect 4302 68 4306 72
rect 4310 68 4314 72
rect 4342 68 4346 72
rect 4414 68 4418 72
rect 4438 68 4442 72
rect 4486 68 4490 72
rect 4590 68 4594 72
rect 4638 68 4642 72
rect 4654 68 4658 72
rect 4790 68 4794 72
rect 4798 68 4802 72
rect 4846 68 4850 72
rect 3550 58 3554 62
rect 3590 58 3594 62
rect 3606 58 3610 62
rect 3646 58 3650 62
rect 3662 58 3666 62
rect 3702 58 3706 62
rect 3742 58 3746 62
rect 3822 58 3826 62
rect 3958 58 3962 62
rect 4022 58 4026 62
rect 4102 59 4106 63
rect 4118 58 4122 62
rect 4214 58 4218 62
rect 4286 58 4290 62
rect 4302 58 4306 62
rect 4470 58 4474 62
rect 4534 58 4538 62
rect 4686 58 4690 62
rect 4758 58 4762 62
rect 4902 68 4906 72
rect 5006 68 5010 72
rect 5038 68 5042 72
rect 5062 68 5066 72
rect 5094 68 5098 72
rect 5102 68 5106 72
rect 5294 68 5298 72
rect 4974 58 4978 62
rect 5038 58 5042 62
rect 5214 58 5218 62
rect 5286 58 5290 62
rect 94 48 98 52
rect 262 48 266 52
rect 294 48 298 52
rect 566 48 570 52
rect 702 48 706 52
rect 710 48 714 52
rect 742 48 746 52
rect 790 48 794 52
rect 822 48 826 52
rect 942 48 946 52
rect 974 48 978 52
rect 1070 48 1074 52
rect 1094 48 1098 52
rect 1102 48 1106 52
rect 1158 48 1162 52
rect 1246 48 1250 52
rect 1286 48 1290 52
rect 1590 48 1594 52
rect 1622 48 1626 52
rect 1630 48 1634 52
rect 1646 48 1650 52
rect 1734 48 1738 52
rect 1838 48 1842 52
rect 2086 48 2090 52
rect 2670 48 2674 52
rect 2742 48 2746 52
rect 2790 48 2794 52
rect 2982 48 2986 52
rect 3070 48 3074 52
rect 3126 48 3130 52
rect 3310 48 3314 52
rect 3326 48 3330 52
rect 3462 48 3466 52
rect 3566 48 3570 52
rect 3598 48 3602 52
rect 3678 48 3682 52
rect 3702 48 3706 52
rect 3750 48 3754 52
rect 3806 48 3810 52
rect 3878 48 3882 52
rect 3886 48 3890 52
rect 4286 48 4290 52
rect 4326 48 4330 52
rect 4358 48 4362 52
rect 5022 48 5026 52
rect 5078 48 5082 52
rect 5118 48 5122 52
rect 5270 48 5274 52
rect 278 38 282 42
rect 958 38 962 42
rect 1142 38 1146 42
rect 1574 38 1578 42
rect 1606 38 1610 42
rect 1654 38 1658 42
rect 1958 38 1962 42
rect 2406 38 2410 42
rect 2694 38 2698 42
rect 2710 38 2714 42
rect 2774 38 2778 42
rect 2998 38 3002 42
rect 3134 38 3138 42
rect 3350 38 3354 42
rect 3486 38 3490 42
rect 3734 38 3738 42
rect 4382 38 4386 42
rect 4598 38 4602 42
rect 4782 38 4786 42
rect 3006 28 3010 32
rect 346 3 350 7
rect 353 3 357 7
rect 1370 3 1374 7
rect 1377 3 1381 7
rect 2394 3 2398 7
rect 2401 3 2405 7
rect 3418 3 3422 7
rect 3425 3 3429 7
rect 4442 3 4446 7
rect 4449 3 4453 7
<< metal2 >>
rect 2206 3728 2210 3732
rect 2686 3728 2690 3732
rect 2718 3728 2722 3732
rect 2758 3731 2762 3732
rect 2750 3728 2762 3731
rect 2942 3728 2946 3732
rect 2982 3731 2986 3732
rect 3166 3731 3170 3732
rect 2974 3728 2986 3731
rect 3158 3728 3170 3731
rect 3286 3728 3290 3732
rect 3302 3728 3306 3732
rect 3374 3731 3378 3732
rect 3398 3731 3402 3732
rect 3630 3731 3634 3732
rect 3374 3728 3385 3731
rect 856 3703 858 3707
rect 862 3703 865 3707
rect 869 3703 872 3707
rect 1872 3703 1874 3707
rect 1878 3703 1881 3707
rect 1885 3703 1888 3707
rect 2206 3702 2209 3728
rect 490 3688 494 3691
rect 6 3679 14 3681
rect 30 3679 38 3681
rect 54 3679 62 3681
rect 78 3679 86 3681
rect 102 3679 110 3681
rect 138 3679 145 3681
rect 6 3678 17 3679
rect 30 3678 41 3679
rect 54 3678 65 3679
rect 78 3678 89 3679
rect 102 3678 113 3679
rect 134 3678 145 3679
rect 162 3679 169 3681
rect 158 3678 169 3679
rect 6 3662 9 3678
rect 30 3662 33 3678
rect 54 3662 57 3678
rect 78 3662 81 3678
rect 102 3662 105 3678
rect 142 3662 145 3678
rect 166 3662 169 3678
rect 198 3679 206 3681
rect 222 3679 230 3681
rect 294 3682 297 3688
rect 198 3678 209 3679
rect 222 3678 233 3679
rect 398 3678 406 3681
rect 198 3662 201 3678
rect 222 3662 225 3678
rect 254 3642 257 3648
rect 262 3642 265 3658
rect 174 3592 177 3638
rect 222 3592 225 3608
rect 170 3568 174 3571
rect 250 3568 254 3571
rect 14 3562 17 3568
rect 262 3562 265 3618
rect 90 3558 94 3561
rect 218 3558 222 3561
rect 118 3552 121 3558
rect 174 3552 177 3558
rect 198 3552 201 3558
rect 218 3548 222 3551
rect 6 3512 9 3528
rect 22 3522 25 3538
rect 6 3472 9 3508
rect 38 3492 41 3548
rect 54 3542 57 3548
rect 126 3542 129 3548
rect 134 3542 137 3548
rect 118 3532 121 3538
rect 230 3532 233 3558
rect 74 3528 78 3531
rect 258 3528 262 3531
rect 62 3488 70 3491
rect 62 3472 65 3488
rect 26 3458 30 3461
rect 54 3392 57 3468
rect 66 3458 70 3461
rect 86 3452 89 3528
rect 150 3522 153 3528
rect 94 3482 97 3518
rect 94 3452 97 3468
rect 102 3462 105 3468
rect 110 3452 113 3478
rect 126 3462 129 3478
rect 142 3471 145 3518
rect 198 3502 201 3528
rect 246 3522 249 3528
rect 142 3468 150 3471
rect 142 3458 150 3461
rect 118 3452 121 3458
rect 54 3362 57 3368
rect 78 3362 81 3368
rect 118 3362 121 3448
rect 134 3442 137 3448
rect 126 3392 129 3418
rect 142 3392 145 3458
rect 174 3392 177 3478
rect 182 3472 185 3478
rect 230 3472 233 3518
rect 246 3472 249 3498
rect 270 3492 273 3648
rect 286 3642 289 3668
rect 310 3652 313 3658
rect 318 3632 321 3678
rect 286 3592 289 3618
rect 326 3601 329 3618
rect 334 3612 337 3638
rect 342 3622 345 3658
rect 350 3632 353 3648
rect 366 3642 369 3668
rect 398 3662 401 3678
rect 374 3622 377 3658
rect 406 3632 409 3668
rect 414 3662 417 3668
rect 422 3662 425 3678
rect 446 3662 449 3678
rect 454 3672 457 3678
rect 478 3675 482 3678
rect 462 3662 465 3668
rect 518 3662 521 3698
rect 538 3678 542 3681
rect 558 3662 561 3698
rect 694 3692 697 3698
rect 1106 3688 1110 3691
rect 1202 3688 1209 3691
rect 834 3678 838 3681
rect 986 3678 990 3681
rect 566 3672 569 3678
rect 622 3672 625 3678
rect 602 3668 606 3671
rect 614 3662 617 3668
rect 344 3603 346 3607
rect 350 3603 353 3607
rect 357 3603 360 3607
rect 318 3598 329 3601
rect 298 3558 302 3561
rect 270 3482 273 3488
rect 202 3458 206 3461
rect 218 3438 222 3441
rect 138 3368 142 3371
rect 162 3368 166 3371
rect 62 3352 65 3358
rect 150 3352 153 3358
rect 182 3352 185 3438
rect 190 3372 193 3418
rect 10 3348 14 3351
rect 6 3312 9 3328
rect 22 3322 25 3338
rect 6 3288 14 3291
rect 6 3272 9 3288
rect 18 3258 22 3261
rect 30 3261 33 3348
rect 54 3332 57 3338
rect 94 3332 97 3338
rect 110 3332 113 3348
rect 126 3332 129 3348
rect 162 3338 166 3341
rect 206 3341 209 3418
rect 202 3338 209 3341
rect 70 3291 73 3318
rect 70 3288 81 3291
rect 54 3282 57 3288
rect 66 3278 70 3281
rect 78 3272 81 3288
rect 50 3268 54 3271
rect 78 3262 81 3268
rect 26 3258 33 3261
rect 38 3252 41 3258
rect 66 3248 70 3251
rect 30 3242 33 3248
rect 86 3242 89 3278
rect 94 3242 97 3328
rect 102 3282 105 3318
rect 110 3272 113 3278
rect 126 3272 129 3288
rect 142 3282 145 3318
rect 134 3272 137 3278
rect 154 3268 158 3271
rect 118 3262 121 3268
rect 166 3262 169 3298
rect 182 3261 185 3328
rect 206 3312 209 3318
rect 206 3272 209 3278
rect 182 3258 190 3261
rect 214 3261 217 3328
rect 222 3302 225 3318
rect 230 3302 233 3468
rect 238 3452 241 3458
rect 246 3352 249 3468
rect 258 3458 262 3461
rect 278 3452 281 3528
rect 286 3522 289 3548
rect 318 3542 321 3598
rect 330 3588 334 3591
rect 430 3562 433 3648
rect 286 3462 289 3518
rect 294 3502 297 3538
rect 306 3528 310 3531
rect 322 3528 326 3531
rect 342 3522 345 3538
rect 326 3472 329 3478
rect 254 3292 257 3348
rect 262 3332 265 3338
rect 270 3332 273 3378
rect 278 3362 281 3448
rect 290 3438 294 3441
rect 286 3362 289 3388
rect 302 3352 305 3468
rect 310 3462 313 3468
rect 318 3462 321 3468
rect 358 3462 361 3468
rect 318 3452 321 3458
rect 374 3432 377 3538
rect 390 3522 393 3558
rect 418 3548 422 3551
rect 398 3542 401 3548
rect 446 3542 449 3618
rect 462 3561 465 3658
rect 542 3592 545 3648
rect 574 3622 577 3648
rect 590 3642 593 3658
rect 606 3632 609 3658
rect 630 3652 633 3678
rect 734 3672 737 3678
rect 670 3662 673 3668
rect 650 3658 654 3661
rect 638 3632 641 3648
rect 654 3642 657 3648
rect 462 3558 470 3561
rect 454 3542 457 3548
rect 470 3542 473 3548
rect 550 3542 553 3578
rect 558 3562 561 3618
rect 622 3592 625 3628
rect 646 3622 649 3628
rect 646 3592 649 3618
rect 670 3572 673 3648
rect 702 3592 705 3668
rect 726 3662 729 3668
rect 742 3622 745 3678
rect 910 3672 913 3678
rect 786 3668 790 3671
rect 774 3652 777 3668
rect 846 3662 849 3668
rect 882 3658 886 3661
rect 798 3652 801 3658
rect 762 3648 766 3651
rect 774 3641 777 3648
rect 766 3638 777 3641
rect 790 3642 793 3648
rect 806 3642 809 3658
rect 822 3652 825 3658
rect 690 3568 694 3571
rect 746 3568 750 3571
rect 758 3562 761 3578
rect 766 3562 769 3638
rect 774 3592 777 3608
rect 806 3591 809 3638
rect 814 3602 817 3638
rect 822 3632 825 3648
rect 830 3612 833 3648
rect 806 3588 817 3591
rect 834 3588 838 3591
rect 642 3558 646 3561
rect 558 3542 561 3548
rect 478 3532 481 3538
rect 506 3518 510 3521
rect 414 3492 417 3498
rect 390 3452 393 3468
rect 438 3462 441 3508
rect 494 3492 497 3518
rect 526 3502 529 3538
rect 534 3532 537 3538
rect 542 3532 545 3538
rect 566 3532 569 3538
rect 574 3482 577 3548
rect 590 3502 593 3518
rect 582 3482 585 3488
rect 606 3482 609 3528
rect 614 3502 617 3538
rect 622 3532 625 3548
rect 630 3491 633 3558
rect 646 3532 649 3548
rect 686 3542 689 3558
rect 714 3548 718 3551
rect 754 3548 758 3551
rect 726 3541 729 3548
rect 718 3538 729 3541
rect 718 3532 721 3538
rect 662 3512 665 3528
rect 718 3492 721 3528
rect 734 3521 737 3538
rect 730 3518 737 3521
rect 630 3488 641 3491
rect 458 3478 462 3481
rect 546 3478 550 3481
rect 446 3472 449 3478
rect 518 3472 521 3478
rect 482 3468 489 3471
rect 450 3458 454 3461
rect 344 3403 346 3407
rect 350 3403 353 3407
rect 357 3403 360 3407
rect 302 3342 305 3348
rect 310 3342 313 3378
rect 358 3352 361 3368
rect 382 3362 385 3368
rect 294 3332 297 3338
rect 314 3328 318 3331
rect 262 3272 265 3318
rect 206 3258 217 3261
rect 266 3258 270 3261
rect 102 3252 105 3258
rect 6 3172 9 3178
rect 14 3132 17 3218
rect 38 3172 41 3178
rect 26 3168 30 3171
rect 30 3142 33 3168
rect 94 3162 97 3168
rect 110 3162 113 3178
rect 134 3172 137 3258
rect 190 3252 193 3258
rect 182 3242 185 3248
rect 166 3182 169 3218
rect 206 3192 209 3258
rect 246 3242 249 3258
rect 270 3232 273 3258
rect 50 3158 54 3161
rect 78 3152 81 3158
rect 58 3148 62 3151
rect 98 3148 102 3151
rect 38 3132 41 3148
rect 54 3132 57 3138
rect 70 3132 73 3138
rect 14 3102 17 3128
rect 54 3082 57 3098
rect 62 3092 65 3118
rect 18 3079 25 3081
rect 14 3078 25 3079
rect 22 3062 25 3078
rect 70 3081 73 3128
rect 62 3078 73 3081
rect 78 3082 81 3148
rect 86 3122 89 3128
rect 54 3052 57 3078
rect 62 3012 65 3078
rect 70 3042 73 3068
rect 82 3058 86 3061
rect 98 3058 102 3061
rect 110 3052 113 3158
rect 122 3148 126 3151
rect 134 3142 137 3168
rect 210 3158 214 3161
rect 142 3142 145 3148
rect 214 3142 217 3158
rect 238 3152 241 3158
rect 270 3142 273 3168
rect 278 3142 281 3308
rect 318 3272 321 3308
rect 326 3292 329 3318
rect 382 3302 385 3358
rect 390 3342 393 3448
rect 398 3412 401 3458
rect 398 3382 401 3408
rect 406 3382 409 3458
rect 478 3422 481 3458
rect 486 3452 489 3468
rect 422 3392 425 3408
rect 446 3382 449 3388
rect 486 3382 489 3448
rect 494 3422 497 3458
rect 506 3438 510 3441
rect 406 3352 409 3378
rect 414 3362 417 3368
rect 410 3338 414 3341
rect 358 3292 361 3298
rect 406 3292 409 3318
rect 422 3302 425 3348
rect 430 3332 433 3368
rect 478 3362 481 3368
rect 518 3362 521 3468
rect 534 3462 537 3478
rect 590 3472 593 3478
rect 614 3472 617 3488
rect 630 3472 633 3478
rect 638 3472 641 3488
rect 702 3488 710 3491
rect 658 3478 662 3481
rect 562 3468 566 3471
rect 550 3462 553 3468
rect 678 3462 681 3478
rect 702 3472 705 3488
rect 766 3472 769 3558
rect 774 3532 777 3588
rect 794 3538 798 3541
rect 634 3458 638 3461
rect 566 3452 569 3458
rect 614 3452 617 3458
rect 670 3452 673 3458
rect 586 3448 590 3451
rect 530 3438 534 3441
rect 526 3392 529 3428
rect 582 3392 585 3418
rect 606 3392 609 3418
rect 562 3378 566 3381
rect 534 3372 537 3378
rect 526 3352 529 3368
rect 550 3362 553 3368
rect 574 3362 577 3368
rect 466 3340 494 3343
rect 550 3342 553 3358
rect 570 3338 574 3341
rect 326 3272 329 3288
rect 414 3282 417 3298
rect 454 3292 457 3338
rect 598 3332 601 3338
rect 478 3322 481 3328
rect 310 3262 313 3268
rect 330 3258 334 3261
rect 286 3192 289 3218
rect 322 3168 326 3171
rect 302 3162 305 3168
rect 314 3158 318 3161
rect 122 3138 126 3141
rect 150 3092 153 3118
rect 174 3112 177 3118
rect 190 3092 193 3138
rect 286 3132 289 3148
rect 306 3128 310 3131
rect 286 3092 289 3128
rect 334 3092 337 3258
rect 350 3222 353 3268
rect 390 3262 393 3278
rect 422 3262 425 3268
rect 446 3262 449 3278
rect 470 3262 473 3268
rect 362 3238 366 3241
rect 344 3203 346 3207
rect 350 3203 353 3207
rect 357 3203 360 3207
rect 374 3192 377 3258
rect 398 3252 401 3258
rect 422 3192 425 3258
rect 366 3172 369 3178
rect 378 3158 382 3161
rect 374 3132 377 3148
rect 398 3142 401 3178
rect 454 3162 457 3168
rect 418 3138 422 3141
rect 346 3128 350 3131
rect 418 3128 422 3131
rect 434 3128 438 3131
rect 258 3088 262 3091
rect 302 3088 310 3091
rect 202 3078 206 3081
rect 254 3072 257 3078
rect 82 3048 86 3051
rect 46 2992 49 3008
rect 94 2992 97 3038
rect 58 2968 62 2971
rect 90 2958 94 2961
rect 46 2952 49 2958
rect 70 2952 73 2958
rect 90 2948 94 2951
rect 6 2931 9 2948
rect 6 2928 14 2931
rect 74 2928 78 2931
rect 22 2892 25 2908
rect 6 2888 14 2891
rect 6 2872 9 2888
rect 54 2862 57 2868
rect 78 2862 81 2928
rect 102 2892 105 2958
rect 118 2952 121 3058
rect 134 3052 137 3058
rect 158 3052 161 3068
rect 174 3062 177 3068
rect 242 3058 246 3061
rect 130 3048 134 3051
rect 174 3042 177 3058
rect 230 3052 233 3058
rect 194 3048 198 3051
rect 218 3048 222 3051
rect 242 3048 249 3051
rect 246 3042 249 3048
rect 222 3032 225 3038
rect 206 3022 209 3028
rect 158 2962 161 2968
rect 190 2962 193 2968
rect 230 2962 233 3028
rect 238 2992 241 3038
rect 254 3032 257 3068
rect 270 3042 273 3068
rect 286 3061 289 3078
rect 294 3072 297 3078
rect 302 3072 305 3088
rect 406 3082 409 3118
rect 414 3092 417 3118
rect 422 3072 425 3078
rect 446 3072 449 3078
rect 394 3068 398 3071
rect 282 3058 289 3061
rect 350 3062 353 3068
rect 454 3062 457 3128
rect 462 3112 465 3258
rect 470 3212 473 3258
rect 486 3242 489 3318
rect 494 3292 497 3328
rect 510 3322 513 3328
rect 574 3282 577 3288
rect 502 3272 505 3278
rect 554 3268 558 3271
rect 554 3258 558 3261
rect 586 3258 590 3261
rect 570 3248 574 3251
rect 494 3242 497 3248
rect 598 3242 601 3328
rect 614 3312 617 3448
rect 630 3412 633 3448
rect 686 3442 689 3468
rect 750 3462 753 3468
rect 758 3422 761 3438
rect 662 3402 665 3418
rect 670 3392 673 3408
rect 630 3372 633 3378
rect 686 3352 689 3388
rect 650 3348 654 3351
rect 678 3348 686 3351
rect 694 3351 697 3418
rect 710 3362 713 3368
rect 694 3348 705 3351
rect 630 3342 633 3348
rect 642 3338 646 3341
rect 678 3332 681 3348
rect 702 3342 705 3348
rect 718 3342 721 3368
rect 766 3362 769 3408
rect 782 3372 785 3498
rect 790 3472 793 3488
rect 806 3482 809 3498
rect 814 3492 817 3588
rect 846 3562 849 3658
rect 854 3582 857 3618
rect 878 3592 881 3638
rect 822 3552 825 3558
rect 822 3492 825 3538
rect 870 3532 873 3558
rect 878 3512 881 3548
rect 856 3503 858 3507
rect 862 3503 865 3507
rect 869 3503 872 3507
rect 842 3478 846 3481
rect 862 3472 865 3488
rect 834 3468 838 3471
rect 846 3468 854 3471
rect 794 3458 798 3461
rect 834 3448 838 3451
rect 814 3442 817 3448
rect 846 3422 849 3468
rect 854 3392 857 3458
rect 798 3362 801 3368
rect 814 3362 817 3368
rect 894 3352 897 3628
rect 902 3552 905 3598
rect 906 3548 910 3551
rect 918 3542 921 3558
rect 934 3552 937 3678
rect 950 3672 953 3678
rect 1046 3672 1049 3678
rect 1078 3672 1081 3688
rect 1206 3672 1209 3688
rect 1214 3682 1217 3688
rect 1222 3682 1225 3688
rect 1446 3682 1449 3698
rect 1566 3688 1574 3691
rect 1738 3688 1742 3691
rect 1778 3688 1782 3691
rect 1274 3678 1281 3681
rect 994 3668 998 3671
rect 1150 3668 1158 3671
rect 958 3662 961 3668
rect 946 3658 950 3661
rect 942 3642 945 3648
rect 966 3622 969 3668
rect 994 3658 998 3661
rect 1050 3658 1054 3661
rect 974 3652 977 3658
rect 1030 3622 1033 3648
rect 1126 3632 1129 3668
rect 1150 3652 1153 3668
rect 1214 3662 1217 3678
rect 1158 3652 1161 3658
rect 1230 3652 1233 3668
rect 1238 3662 1241 3668
rect 1242 3658 1249 3661
rect 910 3532 913 3538
rect 926 3512 929 3548
rect 942 3532 945 3558
rect 966 3552 969 3618
rect 978 3558 982 3561
rect 1030 3552 1033 3618
rect 1158 3592 1161 3648
rect 1190 3592 1193 3618
rect 1222 3592 1225 3628
rect 1230 3622 1233 3648
rect 1230 3571 1233 3618
rect 1238 3602 1241 3618
rect 1230 3568 1241 3571
rect 954 3548 958 3551
rect 994 3548 998 3551
rect 1038 3542 1041 3548
rect 926 3482 929 3488
rect 934 3482 937 3528
rect 950 3512 953 3538
rect 1046 3531 1049 3568
rect 1070 3562 1073 3568
rect 1098 3558 1102 3561
rect 1130 3558 1134 3561
rect 1146 3558 1150 3561
rect 1054 3542 1057 3548
rect 1062 3532 1065 3558
rect 1090 3548 1094 3551
rect 1102 3542 1105 3558
rect 1166 3552 1169 3558
rect 1118 3542 1121 3548
rect 1046 3528 1057 3531
rect 1086 3531 1089 3538
rect 1086 3528 1102 3531
rect 1006 3502 1009 3518
rect 1014 3492 1017 3508
rect 1054 3492 1057 3528
rect 1002 3488 1009 3491
rect 918 3472 921 3478
rect 902 3452 905 3468
rect 942 3452 945 3458
rect 906 3448 910 3451
rect 950 3422 953 3478
rect 1006 3472 1009 3488
rect 1086 3482 1089 3498
rect 1118 3492 1121 3528
rect 1126 3512 1129 3528
rect 1150 3492 1153 3548
rect 1238 3542 1241 3568
rect 1246 3552 1249 3658
rect 1270 3642 1273 3648
rect 1278 3612 1281 3678
rect 1450 3678 1457 3681
rect 1294 3662 1297 3678
rect 1306 3658 1310 3661
rect 1286 3642 1289 3648
rect 1294 3642 1297 3658
rect 1318 3622 1321 3678
rect 1454 3672 1457 3678
rect 1566 3672 1569 3688
rect 1806 3682 1809 3698
rect 1626 3678 1630 3681
rect 1690 3678 1694 3681
rect 1598 3672 1601 3678
rect 1606 3672 1609 3678
rect 1670 3672 1673 3678
rect 1634 3668 1638 3671
rect 1746 3668 1750 3671
rect 1422 3662 1425 3668
rect 1478 3662 1481 3668
rect 1502 3662 1505 3668
rect 1338 3658 1342 3661
rect 1522 3658 1526 3661
rect 1570 3658 1574 3661
rect 1586 3658 1590 3661
rect 1430 3652 1433 3658
rect 1402 3648 1406 3651
rect 1330 3638 1334 3641
rect 1270 3572 1273 3608
rect 1278 3552 1281 3558
rect 1294 3552 1297 3618
rect 1318 3582 1321 3618
rect 1342 3572 1345 3618
rect 1358 3612 1361 3648
rect 1438 3642 1441 3648
rect 1368 3603 1370 3607
rect 1374 3603 1377 3607
rect 1381 3603 1384 3607
rect 1446 3592 1449 3658
rect 1606 3652 1609 3668
rect 1646 3661 1649 3668
rect 1638 3658 1649 3661
rect 1658 3658 1662 3661
rect 1514 3648 1518 3651
rect 1626 3648 1630 3651
rect 1478 3592 1481 3648
rect 1526 3642 1529 3648
rect 1550 3642 1553 3648
rect 1494 3592 1497 3638
rect 1322 3568 1326 3571
rect 1378 3568 1382 3571
rect 1186 3538 1190 3541
rect 1294 3541 1297 3548
rect 1290 3538 1297 3541
rect 1166 3532 1169 3538
rect 1302 3532 1305 3568
rect 1330 3558 1334 3561
rect 1322 3548 1326 3551
rect 1086 3472 1089 3478
rect 1126 3472 1129 3478
rect 1050 3468 1054 3471
rect 958 3432 961 3468
rect 1030 3462 1033 3468
rect 1010 3458 1014 3461
rect 1038 3452 1041 3468
rect 1134 3462 1137 3478
rect 1158 3462 1161 3498
rect 1166 3472 1169 3508
rect 1174 3462 1177 3488
rect 1066 3458 1070 3461
rect 1098 3458 1102 3461
rect 1118 3452 1121 3458
rect 1182 3451 1185 3528
rect 1190 3492 1193 3528
rect 1294 3512 1297 3518
rect 1218 3488 1222 3491
rect 1242 3488 1249 3491
rect 1246 3472 1249 3488
rect 1254 3472 1257 3508
rect 1282 3488 1286 3491
rect 1302 3472 1305 3498
rect 1198 3462 1201 3468
rect 1182 3448 1190 3451
rect 1062 3442 1065 3448
rect 1182 3382 1185 3388
rect 1006 3362 1009 3368
rect 1062 3362 1065 3368
rect 1078 3362 1081 3368
rect 1094 3362 1097 3368
rect 1110 3362 1113 3368
rect 1034 3358 1038 3361
rect 950 3352 953 3358
rect 690 3338 694 3341
rect 730 3340 734 3343
rect 774 3342 777 3348
rect 754 3338 758 3341
rect 874 3338 878 3341
rect 798 3332 801 3338
rect 814 3332 817 3338
rect 714 3328 718 3331
rect 646 3292 649 3318
rect 742 3291 745 3318
rect 734 3288 745 3291
rect 750 3292 753 3328
rect 822 3321 825 3338
rect 822 3318 830 3321
rect 856 3303 858 3307
rect 862 3303 865 3307
rect 869 3303 872 3307
rect 614 3272 617 3278
rect 670 3272 673 3278
rect 606 3252 609 3258
rect 662 3222 665 3268
rect 674 3248 678 3251
rect 690 3238 694 3241
rect 470 3172 473 3178
rect 478 3172 481 3178
rect 526 3162 529 3168
rect 474 3158 478 3161
rect 534 3152 537 3208
rect 566 3192 569 3198
rect 710 3162 713 3228
rect 554 3158 558 3161
rect 478 3142 481 3148
rect 526 3142 529 3148
rect 498 3138 502 3141
rect 510 3132 513 3138
rect 470 3092 473 3128
rect 478 3092 481 3098
rect 494 3062 497 3068
rect 426 3058 430 3061
rect 450 3058 454 3061
rect 278 3052 281 3058
rect 270 2972 273 2978
rect 250 2968 254 2971
rect 130 2958 134 2961
rect 226 2958 230 2961
rect 266 2958 270 2961
rect 146 2948 150 2951
rect 142 2942 145 2948
rect 154 2938 158 2941
rect 118 2932 121 2938
rect 166 2932 169 2958
rect 278 2952 281 3048
rect 398 3032 401 3058
rect 438 3052 441 3058
rect 502 3052 505 3128
rect 534 3122 537 3148
rect 510 3082 513 3098
rect 542 3092 545 3158
rect 582 3142 585 3148
rect 630 3142 633 3148
rect 574 3132 577 3138
rect 638 3132 641 3138
rect 686 3132 689 3138
rect 710 3132 713 3158
rect 574 3092 577 3108
rect 614 3092 617 3118
rect 670 3092 673 3108
rect 718 3092 721 3288
rect 726 3262 729 3278
rect 734 3272 737 3288
rect 782 3272 785 3298
rect 826 3288 830 3291
rect 798 3282 801 3288
rect 866 3278 870 3281
rect 806 3272 809 3278
rect 734 3192 737 3218
rect 782 3152 785 3268
rect 790 3262 793 3268
rect 814 3252 817 3258
rect 794 3248 798 3251
rect 830 3192 833 3278
rect 838 3262 841 3268
rect 854 3242 857 3248
rect 878 3221 881 3258
rect 886 3242 889 3268
rect 878 3218 889 3221
rect 886 3192 889 3218
rect 894 3202 897 3348
rect 918 3332 921 3338
rect 966 3332 969 3338
rect 974 3312 977 3338
rect 990 3332 993 3338
rect 1006 3332 1009 3338
rect 902 3282 905 3298
rect 942 3292 945 3298
rect 966 3292 969 3298
rect 910 3272 913 3278
rect 958 3272 961 3278
rect 982 3272 985 3298
rect 1006 3292 1009 3328
rect 1014 3322 1017 3358
rect 1142 3352 1145 3378
rect 1166 3372 1169 3378
rect 1190 3372 1193 3448
rect 1302 3422 1305 3468
rect 1318 3462 1321 3518
rect 1326 3472 1329 3518
rect 1342 3462 1345 3558
rect 1386 3548 1390 3551
rect 1398 3542 1401 3558
rect 1406 3552 1409 3558
rect 1414 3542 1417 3568
rect 1446 3552 1449 3588
rect 1502 3562 1505 3618
rect 1470 3552 1473 3558
rect 1510 3552 1513 3588
rect 1522 3568 1526 3571
rect 1558 3571 1561 3618
rect 1574 3572 1577 3578
rect 1558 3568 1566 3571
rect 1550 3562 1553 3568
rect 1350 3532 1353 3538
rect 1430 3532 1433 3538
rect 1390 3472 1393 3518
rect 1402 3478 1406 3481
rect 1058 3348 1070 3351
rect 1030 3342 1033 3348
rect 1042 3338 1046 3341
rect 1114 3338 1118 3341
rect 1046 3322 1049 3328
rect 1094 3322 1097 3338
rect 1114 3328 1118 3331
rect 1106 3318 1110 3321
rect 1134 3312 1137 3338
rect 1158 3312 1161 3368
rect 1166 3332 1169 3348
rect 1214 3342 1217 3358
rect 1254 3352 1257 3358
rect 1274 3348 1278 3351
rect 1218 3338 1222 3341
rect 1198 3332 1201 3338
rect 1190 3322 1193 3328
rect 1230 3322 1233 3348
rect 1246 3342 1249 3348
rect 1302 3342 1305 3398
rect 1318 3392 1321 3458
rect 1326 3452 1329 3458
rect 1342 3452 1345 3458
rect 1350 3452 1353 3458
rect 1406 3452 1409 3468
rect 1414 3462 1417 3508
rect 1422 3481 1425 3518
rect 1438 3502 1441 3538
rect 1454 3532 1457 3538
rect 1470 3532 1473 3548
rect 1486 3542 1489 3548
rect 1550 3542 1553 3548
rect 1534 3532 1537 3538
rect 1566 3532 1569 3568
rect 1574 3542 1577 3548
rect 1582 3542 1585 3558
rect 1590 3542 1593 3548
rect 1598 3542 1601 3548
rect 1614 3542 1617 3548
rect 1622 3532 1625 3568
rect 1610 3528 1614 3531
rect 1478 3522 1481 3528
rect 1526 3512 1529 3528
rect 1422 3478 1430 3481
rect 1442 3478 1446 3481
rect 1486 3472 1489 3478
rect 1426 3448 1430 3451
rect 1334 3382 1337 3448
rect 1362 3438 1366 3441
rect 1442 3438 1446 3441
rect 1378 3428 1382 3431
rect 1390 3412 1393 3438
rect 1454 3422 1457 3468
rect 1462 3432 1465 3458
rect 1494 3452 1497 3468
rect 1510 3462 1513 3508
rect 1638 3492 1641 3658
rect 1650 3648 1654 3651
rect 1646 3592 1649 3618
rect 1686 3602 1689 3618
rect 1654 3542 1657 3598
rect 1694 3582 1697 3668
rect 1798 3662 1801 3668
rect 1822 3662 1825 3678
rect 1950 3672 1953 3698
rect 1982 3692 1985 3698
rect 2686 3692 2689 3728
rect 2718 3702 2721 3728
rect 2750 3692 2753 3728
rect 2904 3703 2906 3707
rect 2910 3703 2913 3707
rect 2917 3703 2920 3707
rect 2942 3692 2945 3728
rect 2974 3692 2977 3728
rect 3158 3692 3161 3728
rect 3286 3702 3289 3728
rect 3302 3692 3305 3728
rect 3382 3692 3385 3728
rect 3390 3728 3402 3731
rect 3622 3728 3634 3731
rect 3654 3731 3658 3732
rect 3678 3731 3682 3732
rect 3790 3731 3794 3732
rect 3654 3728 3665 3731
rect 3678 3728 3689 3731
rect 3390 3692 3393 3728
rect 3622 3692 3625 3728
rect 3662 3692 3665 3728
rect 3686 3692 3689 3728
rect 3782 3728 3794 3731
rect 3958 3728 3962 3732
rect 3974 3731 3978 3732
rect 3974 3728 3985 3731
rect 1958 3688 1966 3691
rect 2274 3688 2278 3691
rect 1958 3672 1961 3688
rect 2042 3679 2049 3681
rect 2038 3678 2049 3679
rect 1882 3668 1886 3671
rect 1862 3662 1865 3668
rect 1746 3658 1750 3661
rect 1842 3658 1846 3661
rect 1726 3652 1729 3658
rect 1822 3652 1825 3658
rect 1902 3652 1905 3668
rect 1910 3662 1913 3668
rect 1966 3662 1969 3678
rect 1998 3671 2001 3678
rect 1990 3668 2001 3671
rect 1982 3662 1985 3668
rect 1954 3658 1958 3661
rect 1934 3652 1937 3658
rect 1858 3648 1862 3651
rect 1990 3651 1993 3668
rect 2046 3662 2049 3678
rect 2070 3679 2078 3681
rect 2070 3678 2081 3679
rect 2206 3679 2214 3681
rect 2230 3682 2233 3688
rect 2254 3682 2257 3688
rect 2310 3682 2313 3688
rect 2550 3682 2553 3688
rect 2206 3678 2217 3679
rect 2450 3678 2454 3681
rect 2590 3679 2598 3681
rect 2614 3679 2622 3681
rect 2638 3682 2641 3688
rect 3110 3682 3113 3688
rect 3318 3682 3321 3688
rect 2590 3678 2601 3679
rect 2614 3678 2625 3679
rect 2002 3658 2006 3661
rect 1986 3648 1993 3651
rect 1830 3642 1833 3648
rect 1838 3642 1841 3648
rect 1850 3638 1854 3641
rect 1686 3562 1689 3568
rect 1726 3562 1729 3638
rect 1742 3562 1745 3588
rect 1806 3572 1809 3638
rect 1750 3562 1753 3568
rect 1662 3552 1665 3558
rect 1646 3491 1649 3518
rect 1662 3512 1665 3548
rect 1710 3542 1713 3548
rect 1718 3542 1721 3548
rect 1726 3542 1729 3558
rect 1758 3552 1761 3568
rect 1766 3562 1769 3568
rect 1786 3548 1790 3551
rect 1742 3532 1745 3538
rect 1758 3532 1761 3538
rect 1686 3492 1689 3518
rect 1646 3488 1657 3491
rect 1518 3472 1521 3478
rect 1622 3475 1626 3478
rect 1578 3468 1582 3471
rect 1526 3451 1529 3468
rect 1598 3462 1601 3468
rect 1514 3448 1529 3451
rect 1486 3432 1489 3448
rect 1368 3403 1370 3407
rect 1374 3403 1377 3407
rect 1381 3403 1384 3407
rect 1422 3352 1425 3358
rect 1430 3342 1433 3418
rect 1462 3392 1465 3408
rect 1494 3402 1497 3448
rect 1554 3438 1558 3441
rect 1558 3392 1561 3428
rect 1446 3352 1449 3388
rect 1454 3342 1457 3358
rect 1486 3352 1489 3388
rect 1518 3382 1521 3388
rect 1566 3362 1569 3368
rect 1538 3358 1542 3361
rect 1578 3358 1582 3361
rect 1498 3348 1502 3351
rect 1478 3342 1481 3348
rect 1354 3338 1358 3341
rect 1370 3338 1374 3341
rect 1238 3332 1241 3338
rect 1470 3332 1473 3338
rect 1510 3332 1513 3358
rect 1550 3352 1553 3358
rect 1542 3342 1545 3348
rect 1558 3342 1561 3348
rect 1590 3342 1593 3458
rect 1606 3452 1609 3468
rect 1654 3462 1657 3488
rect 1662 3482 1665 3488
rect 1694 3482 1697 3518
rect 1678 3472 1681 3478
rect 1686 3472 1689 3478
rect 1694 3472 1697 3478
rect 1666 3468 1670 3471
rect 1710 3462 1713 3478
rect 1738 3468 1742 3471
rect 1682 3458 1686 3461
rect 1730 3458 1734 3461
rect 1750 3452 1753 3458
rect 1602 3448 1606 3451
rect 1718 3442 1721 3448
rect 1758 3442 1761 3518
rect 1766 3462 1769 3508
rect 1782 3482 1785 3518
rect 1790 3462 1793 3498
rect 1806 3492 1809 3568
rect 1814 3542 1817 3548
rect 1838 3542 1841 3618
rect 1890 3558 1894 3561
rect 1846 3552 1849 3558
rect 1858 3548 1862 3551
rect 1902 3542 1905 3568
rect 1926 3552 1929 3618
rect 1934 3562 1937 3568
rect 1910 3542 1913 3548
rect 1866 3538 1870 3541
rect 1822 3532 1825 3538
rect 1838 3532 1841 3538
rect 1814 3482 1817 3528
rect 1830 3462 1833 3498
rect 1846 3482 1849 3498
rect 1854 3492 1857 3538
rect 1918 3532 1921 3548
rect 1872 3503 1874 3507
rect 1878 3503 1881 3507
rect 1885 3503 1888 3507
rect 1918 3492 1921 3528
rect 1926 3482 1929 3538
rect 1942 3532 1945 3548
rect 1950 3532 1953 3548
rect 1958 3542 1961 3558
rect 1962 3518 1966 3521
rect 1990 3502 1993 3648
rect 2006 3622 2009 3658
rect 2054 3632 2057 3678
rect 2070 3662 2073 3678
rect 2094 3672 2097 3678
rect 2194 3668 2198 3671
rect 2206 3662 2209 3678
rect 2098 3658 2102 3661
rect 2122 3658 2126 3661
rect 2142 3652 2145 3658
rect 2062 3642 2065 3648
rect 2134 3642 2137 3648
rect 2150 3642 2153 3658
rect 2174 3652 2177 3658
rect 2114 3638 2118 3641
rect 2126 3582 2129 3618
rect 2014 3552 2017 3558
rect 2030 3552 2033 3558
rect 2046 3542 2049 3548
rect 2070 3542 2073 3548
rect 2134 3541 2137 3598
rect 2150 3571 2153 3618
rect 2158 3592 2161 3638
rect 2150 3568 2161 3571
rect 2170 3568 2174 3571
rect 2130 3538 2137 3541
rect 2006 3532 2009 3538
rect 2062 3492 2065 3498
rect 1966 3482 1969 3488
rect 1858 3478 1862 3481
rect 1902 3470 1905 3478
rect 2022 3472 2025 3488
rect 2078 3472 2081 3508
rect 1854 3462 1857 3468
rect 1814 3452 1817 3458
rect 1778 3448 1782 3451
rect 1598 3352 1601 3398
rect 1662 3382 1665 3418
rect 1734 3372 1737 3418
rect 1714 3348 1718 3351
rect 1622 3342 1625 3348
rect 1630 3342 1633 3348
rect 1734 3342 1737 3368
rect 1774 3362 1777 3368
rect 1774 3342 1777 3348
rect 1782 3342 1785 3378
rect 1798 3342 1801 3348
rect 1814 3342 1817 3438
rect 1870 3392 1873 3468
rect 1894 3462 1897 3468
rect 1962 3468 1966 3471
rect 1942 3452 1945 3458
rect 1958 3382 1961 3418
rect 2006 3372 2009 3418
rect 2030 3402 2033 3468
rect 2086 3462 2089 3468
rect 2086 3392 2089 3458
rect 2094 3402 2097 3518
rect 2118 3512 2121 3538
rect 2142 3522 2145 3558
rect 2150 3552 2153 3558
rect 2158 3552 2161 3568
rect 2182 3562 2185 3658
rect 2190 3632 2193 3658
rect 2182 3552 2185 3558
rect 2190 3552 2193 3628
rect 2158 3532 2161 3548
rect 2162 3518 2166 3521
rect 2134 3482 2137 3518
rect 2142 3482 2145 3518
rect 2158 3492 2161 3508
rect 2182 3491 2185 3548
rect 2190 3532 2193 3538
rect 2206 3532 2209 3558
rect 2214 3542 2217 3668
rect 2234 3648 2238 3651
rect 2246 3622 2249 3668
rect 2254 3662 2257 3678
rect 2274 3668 2278 3671
rect 2286 3662 2289 3678
rect 2294 3662 2297 3678
rect 2318 3662 2321 3678
rect 2358 3672 2361 3678
rect 2442 3668 2446 3671
rect 2270 3652 2273 3658
rect 2302 3652 2305 3658
rect 2342 3652 2345 3658
rect 2390 3652 2393 3658
rect 2398 3652 2401 3658
rect 2422 3652 2425 3658
rect 2362 3648 2366 3651
rect 2318 3642 2321 3648
rect 2330 3638 2334 3641
rect 2378 3638 2382 3641
rect 2342 3622 2345 3628
rect 2394 3618 2398 3621
rect 2270 3592 2273 3598
rect 2238 3562 2241 3588
rect 2286 3582 2289 3618
rect 2392 3603 2394 3607
rect 2398 3603 2401 3607
rect 2405 3603 2408 3607
rect 2298 3588 2302 3591
rect 2422 3582 2425 3648
rect 2430 3632 2433 3668
rect 2450 3648 2454 3651
rect 2462 3632 2465 3658
rect 2470 3642 2473 3678
rect 2494 3652 2497 3678
rect 2546 3668 2553 3671
rect 2514 3658 2518 3661
rect 2538 3658 2542 3661
rect 2530 3648 2534 3651
rect 2474 3638 2478 3641
rect 2490 3638 2494 3641
rect 2482 3628 2486 3631
rect 2510 3622 2513 3638
rect 2550 3622 2553 3668
rect 2558 3652 2561 3678
rect 2590 3662 2593 3678
rect 2614 3662 2617 3678
rect 2918 3672 2921 3678
rect 2654 3662 2657 3668
rect 2678 3662 2681 3668
rect 2642 3658 2646 3661
rect 2518 3612 2521 3618
rect 2558 3592 2561 3648
rect 2662 3632 2665 3648
rect 2662 3602 2665 3628
rect 2678 3612 2681 3618
rect 2278 3572 2281 3578
rect 2626 3568 2630 3571
rect 2666 3568 2670 3571
rect 2278 3562 2281 3568
rect 2366 3562 2369 3568
rect 2250 3558 2254 3561
rect 2262 3552 2265 3558
rect 2226 3548 2230 3551
rect 2254 3548 2262 3551
rect 2198 3492 2201 3518
rect 2214 3512 2217 3538
rect 2254 3532 2257 3548
rect 2270 3532 2273 3548
rect 2298 3528 2302 3531
rect 2238 3522 2241 3528
rect 2310 3522 2313 3548
rect 2318 3542 2321 3558
rect 2362 3548 2366 3551
rect 2402 3548 2406 3551
rect 2334 3532 2337 3548
rect 2342 3521 2345 3538
rect 2350 3532 2353 3548
rect 2414 3542 2417 3558
rect 2438 3552 2441 3558
rect 2446 3552 2449 3558
rect 2454 3532 2457 3568
rect 2514 3558 2518 3561
rect 2494 3552 2497 3558
rect 2394 3528 2398 3531
rect 2426 3528 2430 3531
rect 2342 3518 2350 3521
rect 2182 3488 2193 3491
rect 2258 3488 2262 3491
rect 2106 3468 2110 3471
rect 2122 3468 2129 3471
rect 2138 3468 2142 3471
rect 2106 3458 2110 3461
rect 2126 3452 2129 3468
rect 2106 3448 2110 3451
rect 2126 3392 2129 3448
rect 2134 3442 2137 3448
rect 1842 3368 1846 3371
rect 2086 3368 2094 3371
rect 2138 3368 2142 3371
rect 2154 3368 2158 3371
rect 1826 3358 1830 3361
rect 2074 3358 2078 3361
rect 1862 3352 1865 3358
rect 1902 3352 1905 3358
rect 2058 3348 2062 3351
rect 2074 3348 2078 3351
rect 1634 3338 1641 3341
rect 1590 3332 1593 3338
rect 1638 3332 1641 3338
rect 1746 3338 1750 3341
rect 1610 3328 1614 3331
rect 1046 3292 1049 3308
rect 1134 3292 1137 3298
rect 1034 3288 1038 3291
rect 1078 3282 1081 3288
rect 994 3278 998 3281
rect 1014 3272 1017 3278
rect 902 3262 905 3268
rect 910 3262 913 3268
rect 1022 3262 1025 3268
rect 1066 3258 1070 3261
rect 1098 3258 1102 3261
rect 966 3242 969 3248
rect 926 3192 929 3238
rect 858 3188 862 3191
rect 774 3142 777 3148
rect 798 3142 801 3188
rect 938 3168 942 3171
rect 954 3168 958 3171
rect 614 3072 617 3078
rect 674 3068 678 3071
rect 746 3068 750 3071
rect 418 3048 422 3051
rect 474 3048 478 3051
rect 344 3003 346 3007
rect 350 3003 353 3007
rect 357 3003 360 3007
rect 382 2962 385 2968
rect 290 2958 294 2961
rect 194 2948 198 2951
rect 242 2948 246 2951
rect 330 2948 334 2951
rect 386 2948 390 2951
rect 198 2932 201 2938
rect 150 2892 153 2918
rect 166 2892 169 2928
rect 206 2922 209 2948
rect 194 2888 198 2891
rect 146 2878 150 2881
rect 86 2872 89 2878
rect 158 2872 161 2878
rect 146 2868 153 2871
rect 102 2842 105 2858
rect 102 2832 105 2838
rect 82 2768 86 2771
rect 98 2768 102 2771
rect 54 2762 57 2768
rect 62 2752 65 2758
rect 22 2701 25 2748
rect 30 2731 33 2748
rect 70 2742 73 2748
rect 42 2738 46 2741
rect 30 2728 41 2731
rect 58 2728 62 2731
rect 22 2698 30 2701
rect 30 2682 33 2698
rect 6 2612 9 2658
rect 30 2562 33 2568
rect 38 2552 41 2728
rect 70 2721 73 2738
rect 78 2732 81 2768
rect 110 2752 113 2758
rect 134 2752 137 2848
rect 86 2742 89 2748
rect 142 2742 145 2758
rect 102 2732 105 2738
rect 62 2718 73 2721
rect 62 2692 65 2718
rect 118 2692 121 2738
rect 150 2732 153 2868
rect 162 2858 166 2861
rect 170 2848 174 2851
rect 174 2752 177 2758
rect 182 2752 185 2858
rect 190 2822 193 2868
rect 78 2688 86 2691
rect 70 2672 73 2678
rect 78 2672 81 2688
rect 166 2682 169 2718
rect 110 2672 113 2678
rect 118 2672 121 2678
rect 138 2668 142 2671
rect 46 2552 49 2658
rect 54 2652 57 2668
rect 82 2658 86 2661
rect 98 2658 102 2661
rect 118 2622 121 2668
rect 158 2662 161 2668
rect 166 2652 169 2658
rect 174 2652 177 2738
rect 190 2732 193 2818
rect 210 2738 214 2741
rect 182 2692 185 2728
rect 222 2712 225 2758
rect 230 2692 233 2948
rect 278 2932 281 2938
rect 278 2872 281 2888
rect 294 2882 297 2938
rect 314 2928 318 2931
rect 342 2922 345 2948
rect 398 2942 401 3028
rect 406 2992 409 3038
rect 438 2992 441 3048
rect 510 2992 513 3048
rect 450 2958 454 2961
rect 390 2938 398 2941
rect 390 2932 393 2938
rect 378 2928 382 2931
rect 310 2892 313 2898
rect 390 2892 393 2928
rect 398 2882 401 2908
rect 406 2892 409 2958
rect 422 2942 425 2958
rect 526 2952 529 3058
rect 534 3052 537 3068
rect 550 3062 553 3068
rect 550 2992 553 3058
rect 558 3032 561 3068
rect 574 2992 577 3048
rect 594 2988 598 2991
rect 586 2958 590 2961
rect 434 2938 441 2941
rect 438 2912 441 2938
rect 422 2882 425 2908
rect 294 2872 297 2878
rect 422 2872 425 2878
rect 438 2872 441 2908
rect 342 2862 345 2868
rect 254 2792 257 2848
rect 262 2821 265 2859
rect 262 2818 273 2821
rect 262 2772 265 2778
rect 238 2762 241 2768
rect 246 2742 249 2758
rect 254 2712 257 2748
rect 262 2682 265 2748
rect 198 2662 201 2668
rect 186 2648 190 2651
rect 126 2642 129 2648
rect 142 2642 145 2648
rect 154 2638 158 2641
rect 94 2592 97 2608
rect 118 2572 121 2618
rect 18 2548 22 2551
rect 6 2521 9 2538
rect 54 2532 57 2548
rect 62 2542 65 2558
rect 118 2542 121 2548
rect 126 2531 129 2548
rect 122 2528 129 2531
rect 134 2532 137 2538
rect 6 2518 14 2521
rect 6 2479 14 2481
rect 30 2482 33 2518
rect 38 2492 41 2528
rect 106 2518 110 2521
rect 118 2492 121 2528
rect 142 2492 145 2558
rect 166 2552 169 2628
rect 206 2612 209 2668
rect 254 2632 257 2668
rect 262 2652 265 2678
rect 270 2582 273 2818
rect 278 2792 281 2858
rect 366 2811 369 2868
rect 434 2858 438 2861
rect 374 2822 377 2858
rect 446 2852 449 2928
rect 478 2892 481 2948
rect 486 2922 489 2928
rect 494 2912 497 2938
rect 542 2932 545 2938
rect 502 2872 505 2908
rect 510 2892 513 2908
rect 366 2808 377 2811
rect 344 2803 346 2807
rect 350 2803 353 2807
rect 357 2803 360 2807
rect 374 2792 377 2808
rect 446 2802 449 2848
rect 302 2772 305 2778
rect 278 2752 281 2758
rect 350 2752 353 2768
rect 338 2748 342 2751
rect 278 2652 281 2748
rect 366 2742 369 2748
rect 298 2728 302 2731
rect 310 2722 313 2738
rect 342 2732 345 2738
rect 390 2732 393 2758
rect 414 2742 417 2768
rect 426 2748 430 2751
rect 322 2728 326 2731
rect 418 2728 422 2731
rect 298 2668 302 2671
rect 298 2658 302 2661
rect 314 2658 318 2661
rect 306 2648 310 2651
rect 326 2642 329 2688
rect 358 2682 361 2718
rect 390 2692 393 2708
rect 414 2692 417 2718
rect 454 2692 457 2868
rect 470 2792 473 2818
rect 550 2792 553 2938
rect 558 2932 561 2958
rect 570 2948 574 2951
rect 566 2921 569 2938
rect 606 2922 609 3068
rect 666 3058 670 3061
rect 670 3042 673 3048
rect 686 2972 689 3068
rect 694 2981 697 3068
rect 746 3058 750 3061
rect 754 3038 758 3041
rect 702 2992 705 3038
rect 766 2992 769 3138
rect 790 3072 793 3128
rect 798 3091 801 3138
rect 798 3088 809 3091
rect 778 3068 782 3071
rect 778 3058 782 3061
rect 798 3052 801 3078
rect 806 3072 809 3088
rect 822 3072 825 3118
rect 830 3102 833 3118
rect 846 3102 849 3138
rect 878 3132 881 3138
rect 856 3103 858 3107
rect 862 3103 865 3107
rect 869 3103 872 3107
rect 878 3092 881 3128
rect 894 3092 897 3168
rect 902 3132 905 3148
rect 910 3102 913 3158
rect 918 3122 921 3158
rect 982 3152 985 3248
rect 990 3242 993 3248
rect 1006 3242 1009 3258
rect 1046 3252 1049 3258
rect 990 3171 993 3238
rect 1038 3222 1041 3248
rect 1134 3192 1137 3218
rect 1142 3192 1145 3238
rect 1150 3222 1153 3268
rect 1158 3252 1161 3258
rect 1190 3252 1193 3318
rect 1262 3292 1265 3328
rect 1270 3322 1273 3328
rect 1654 3322 1657 3338
rect 1702 3332 1705 3338
rect 1774 3332 1777 3338
rect 1330 3318 1334 3321
rect 1286 3292 1289 3318
rect 1350 3292 1353 3298
rect 1246 3282 1249 3288
rect 1254 3282 1257 3288
rect 1198 3232 1201 3268
rect 1206 3242 1209 3278
rect 1350 3275 1354 3278
rect 1390 3272 1393 3288
rect 1454 3282 1457 3288
rect 1470 3282 1473 3318
rect 1442 3278 1446 3281
rect 1222 3262 1225 3268
rect 1222 3182 1225 3258
rect 1230 3192 1233 3258
rect 1250 3248 1254 3251
rect 1262 3192 1265 3248
rect 1270 3222 1273 3268
rect 1278 3252 1281 3258
rect 1286 3242 1289 3268
rect 1294 3252 1297 3258
rect 1294 3232 1297 3248
rect 1310 3192 1313 3248
rect 1318 3192 1321 3258
rect 1366 3241 1369 3268
rect 1358 3238 1369 3241
rect 1358 3192 1361 3238
rect 1368 3203 1370 3207
rect 1374 3203 1377 3207
rect 1381 3203 1384 3207
rect 1182 3172 1185 3178
rect 990 3168 998 3171
rect 1194 3168 1198 3171
rect 1210 3168 1214 3171
rect 998 3152 1001 3168
rect 1190 3162 1193 3168
rect 926 3142 929 3148
rect 966 3142 969 3148
rect 1006 3142 1009 3148
rect 1062 3142 1065 3158
rect 958 3102 961 3128
rect 974 3122 977 3138
rect 990 3102 993 3138
rect 942 3092 945 3098
rect 1006 3092 1009 3128
rect 1054 3121 1057 3138
rect 1050 3118 1057 3121
rect 1038 3102 1041 3118
rect 1078 3092 1081 3118
rect 838 3072 841 3078
rect 810 3058 814 3061
rect 846 3052 849 3078
rect 918 3072 921 3078
rect 910 3052 913 3068
rect 926 3062 929 3088
rect 950 3082 953 3088
rect 962 3068 966 3071
rect 974 3062 977 3088
rect 1038 3082 1041 3088
rect 1094 3082 1097 3118
rect 1110 3092 1113 3138
rect 1142 3132 1145 3158
rect 1166 3142 1169 3148
rect 1174 3141 1177 3158
rect 1214 3152 1217 3158
rect 1238 3152 1241 3178
rect 1274 3168 1278 3171
rect 1290 3168 1294 3171
rect 1250 3158 1254 3161
rect 1270 3152 1273 3168
rect 1170 3138 1177 3141
rect 1158 3132 1161 3138
rect 1182 3132 1185 3148
rect 1122 3128 1129 3131
rect 1126 3092 1129 3128
rect 1134 3082 1137 3118
rect 1034 3078 1038 3081
rect 990 3062 993 3068
rect 1038 3062 1041 3068
rect 1094 3062 1097 3068
rect 1110 3062 1113 3068
rect 962 3058 966 3061
rect 1010 3058 1014 3061
rect 1058 3058 1062 3061
rect 834 3048 838 3051
rect 994 3048 998 3051
rect 886 3042 889 3048
rect 902 2992 905 3018
rect 786 2988 790 2991
rect 742 2982 745 2988
rect 694 2978 705 2981
rect 694 2952 697 2958
rect 662 2942 665 2947
rect 566 2918 574 2921
rect 630 2892 633 2938
rect 694 2922 697 2938
rect 590 2872 593 2888
rect 658 2868 662 2871
rect 574 2822 577 2859
rect 482 2768 486 2771
rect 538 2768 542 2771
rect 462 2722 465 2758
rect 494 2752 497 2758
rect 374 2672 377 2678
rect 414 2672 417 2678
rect 430 2672 433 2678
rect 462 2672 465 2708
rect 470 2702 473 2748
rect 514 2740 518 2743
rect 526 2742 529 2758
rect 590 2752 593 2868
rect 606 2832 609 2868
rect 626 2858 630 2861
rect 658 2858 662 2861
rect 678 2842 681 2878
rect 642 2788 646 2791
rect 678 2752 681 2758
rect 546 2738 550 2741
rect 486 2692 489 2738
rect 526 2732 529 2738
rect 518 2692 521 2728
rect 558 2692 561 2698
rect 606 2692 609 2728
rect 614 2711 617 2747
rect 614 2708 625 2711
rect 506 2688 513 2691
rect 578 2688 582 2691
rect 346 2668 350 2671
rect 442 2668 446 2671
rect 382 2662 385 2668
rect 406 2662 409 2668
rect 466 2658 470 2661
rect 438 2652 441 2658
rect 454 2652 457 2658
rect 478 2652 481 2678
rect 510 2672 513 2688
rect 614 2682 617 2698
rect 614 2672 617 2678
rect 586 2668 590 2671
rect 534 2662 537 2668
rect 502 2652 505 2658
rect 542 2652 545 2668
rect 550 2662 553 2668
rect 394 2648 398 2651
rect 418 2648 422 2651
rect 278 2572 281 2618
rect 190 2558 198 2561
rect 274 2558 278 2561
rect 154 2548 158 2551
rect 170 2538 174 2541
rect 150 2532 153 2538
rect 190 2532 193 2558
rect 310 2552 313 2568
rect 318 2552 321 2618
rect 344 2603 346 2607
rect 350 2603 353 2607
rect 357 2603 360 2607
rect 446 2592 449 2648
rect 346 2588 350 2591
rect 414 2552 417 2558
rect 454 2552 457 2648
rect 478 2642 481 2648
rect 542 2592 545 2648
rect 550 2592 553 2658
rect 562 2648 566 2651
rect 574 2592 577 2668
rect 602 2658 614 2661
rect 486 2582 489 2588
rect 586 2558 590 2561
rect 546 2548 550 2551
rect 262 2542 265 2548
rect 302 2542 305 2548
rect 202 2538 206 2541
rect 314 2538 318 2541
rect 6 2478 17 2479
rect 90 2478 94 2481
rect 6 2462 9 2478
rect 78 2472 81 2478
rect 38 2468 46 2471
rect 38 2442 41 2468
rect 58 2458 62 2461
rect 66 2438 70 2441
rect 78 2441 81 2458
rect 86 2452 89 2478
rect 110 2472 113 2478
rect 118 2468 126 2471
rect 118 2452 121 2468
rect 142 2462 145 2488
rect 78 2438 89 2441
rect 14 2362 17 2368
rect 14 2332 17 2338
rect 22 2292 25 2408
rect 38 2392 41 2438
rect 86 2392 89 2438
rect 118 2392 121 2448
rect 134 2442 137 2458
rect 150 2442 153 2478
rect 170 2468 174 2471
rect 158 2452 161 2458
rect 190 2452 193 2458
rect 166 2442 169 2448
rect 30 2372 33 2378
rect 74 2368 110 2371
rect 118 2362 121 2368
rect 166 2362 169 2438
rect 198 2422 201 2518
rect 206 2492 209 2528
rect 254 2521 257 2538
rect 246 2518 257 2521
rect 246 2492 249 2518
rect 294 2492 297 2518
rect 314 2478 318 2481
rect 362 2478 366 2481
rect 214 2472 217 2478
rect 294 2472 297 2478
rect 322 2468 326 2471
rect 246 2462 249 2468
rect 222 2412 225 2458
rect 270 2452 273 2458
rect 278 2452 281 2468
rect 278 2441 281 2448
rect 270 2438 281 2441
rect 294 2442 297 2468
rect 366 2462 369 2478
rect 374 2472 377 2488
rect 306 2458 310 2461
rect 334 2452 337 2458
rect 198 2392 201 2408
rect 270 2392 273 2438
rect 302 2372 305 2418
rect 310 2392 313 2438
rect 382 2422 385 2428
rect 346 2418 350 2421
rect 38 2352 41 2358
rect 54 2332 57 2358
rect 166 2352 169 2358
rect 154 2348 158 2351
rect 86 2342 89 2348
rect 118 2342 121 2348
rect 154 2338 161 2341
rect 54 2312 57 2328
rect 6 2288 14 2291
rect 6 2272 9 2288
rect 54 2262 57 2268
rect 62 2262 65 2288
rect 94 2271 97 2338
rect 158 2332 161 2338
rect 142 2292 145 2318
rect 114 2288 118 2291
rect 158 2272 161 2328
rect 174 2312 177 2358
rect 190 2292 193 2368
rect 198 2362 201 2368
rect 282 2358 286 2361
rect 202 2348 206 2351
rect 234 2348 238 2351
rect 222 2342 225 2348
rect 186 2278 190 2281
rect 206 2272 209 2308
rect 214 2302 217 2338
rect 254 2332 257 2358
rect 270 2342 273 2348
rect 302 2342 305 2368
rect 326 2361 329 2418
rect 344 2403 346 2407
rect 350 2403 353 2407
rect 357 2403 360 2407
rect 382 2392 385 2408
rect 390 2392 393 2548
rect 438 2512 441 2528
rect 454 2522 457 2548
rect 454 2492 457 2508
rect 478 2502 481 2548
rect 502 2542 505 2548
rect 518 2532 521 2548
rect 498 2528 502 2531
rect 510 2492 513 2518
rect 518 2492 521 2518
rect 526 2512 529 2528
rect 542 2472 545 2508
rect 486 2462 489 2468
rect 494 2462 497 2468
rect 398 2412 401 2448
rect 414 2442 417 2458
rect 322 2358 329 2361
rect 326 2352 329 2358
rect 490 2388 494 2391
rect 314 2348 318 2351
rect 330 2338 334 2341
rect 246 2302 249 2318
rect 254 2312 257 2328
rect 218 2278 222 2281
rect 230 2272 233 2298
rect 262 2292 265 2338
rect 270 2292 273 2298
rect 350 2292 353 2388
rect 418 2368 422 2371
rect 478 2362 481 2388
rect 502 2372 505 2418
rect 486 2362 489 2368
rect 434 2348 438 2351
rect 362 2338 366 2341
rect 374 2332 377 2348
rect 374 2322 377 2328
rect 390 2292 393 2338
rect 414 2332 417 2348
rect 426 2338 430 2341
rect 402 2318 406 2321
rect 414 2292 417 2328
rect 454 2322 457 2358
rect 518 2352 521 2358
rect 498 2348 502 2351
rect 502 2338 510 2341
rect 286 2272 289 2288
rect 314 2278 318 2281
rect 402 2278 406 2281
rect 478 2281 481 2318
rect 502 2292 505 2338
rect 518 2322 521 2328
rect 526 2292 529 2458
rect 550 2392 553 2548
rect 558 2532 561 2558
rect 570 2548 574 2551
rect 566 2521 569 2538
rect 598 2532 601 2538
rect 566 2518 574 2521
rect 606 2492 609 2658
rect 622 2612 625 2708
rect 638 2672 641 2718
rect 654 2692 657 2738
rect 686 2692 689 2918
rect 702 2892 705 2978
rect 710 2942 713 2978
rect 766 2972 769 2978
rect 722 2948 726 2951
rect 762 2948 766 2951
rect 718 2932 721 2938
rect 734 2892 737 2948
rect 762 2938 766 2941
rect 782 2932 785 2958
rect 854 2942 857 2947
rect 870 2942 873 2948
rect 754 2928 758 2931
rect 822 2922 825 2938
rect 856 2903 858 2907
rect 862 2903 865 2907
rect 869 2903 872 2907
rect 910 2902 913 3048
rect 1006 3042 1009 3048
rect 1014 3042 1017 3058
rect 1050 3038 1054 3041
rect 934 2932 937 2938
rect 942 2932 945 3038
rect 1006 2992 1009 3038
rect 1062 3032 1065 3038
rect 1014 2992 1017 2998
rect 966 2951 969 2958
rect 1070 2942 1073 3048
rect 1082 3038 1086 3041
rect 1102 3032 1105 3048
rect 1118 3042 1121 3068
rect 1134 3032 1137 3078
rect 1142 3072 1145 3108
rect 1174 3082 1177 3098
rect 1150 3062 1153 3078
rect 1174 3062 1177 3068
rect 1190 3062 1193 3098
rect 1118 2992 1121 3028
rect 1138 2958 1142 2961
rect 1122 2948 1126 2951
rect 1150 2951 1153 3058
rect 1166 2972 1169 3048
rect 1190 3042 1193 3048
rect 1146 2948 1153 2951
rect 1078 2942 1081 2947
rect 1158 2942 1161 2948
rect 982 2912 985 2938
rect 998 2932 1001 2938
rect 838 2892 841 2898
rect 934 2892 937 2898
rect 1038 2892 1041 2908
rect 1070 2892 1073 2938
rect 762 2888 766 2891
rect 1078 2882 1081 2928
rect 1110 2902 1113 2938
rect 1166 2932 1169 2958
rect 1198 2952 1201 2958
rect 1206 2952 1209 3138
rect 1214 3132 1217 3148
rect 1226 3138 1230 3141
rect 1246 3132 1249 3148
rect 1262 3142 1265 3148
rect 1302 3132 1305 3138
rect 1334 3132 1337 3138
rect 1274 3128 1278 3131
rect 1214 3122 1217 3128
rect 1294 3122 1297 3128
rect 1214 3092 1217 3108
rect 1238 3062 1241 3098
rect 1262 3072 1265 3118
rect 1270 3062 1273 3098
rect 1218 3058 1222 3061
rect 1254 3052 1257 3058
rect 1286 3052 1289 3058
rect 1226 3048 1230 3051
rect 1238 3042 1241 3048
rect 1294 3042 1297 3118
rect 1342 3112 1345 3148
rect 1350 3142 1353 3158
rect 1390 3152 1393 3248
rect 1426 3188 1430 3191
rect 1398 3158 1406 3161
rect 1350 3092 1353 3128
rect 1366 3112 1369 3138
rect 1374 3122 1377 3138
rect 1390 3132 1393 3148
rect 1398 3092 1401 3158
rect 1406 3152 1409 3158
rect 1362 3078 1366 3081
rect 1302 3072 1305 3078
rect 1406 3072 1409 3138
rect 1414 3122 1417 3158
rect 1422 3152 1425 3158
rect 1430 3142 1433 3168
rect 1438 3102 1441 3268
rect 1446 3262 1449 3268
rect 1486 3262 1489 3268
rect 1462 3252 1465 3258
rect 1510 3252 1513 3258
rect 1470 3192 1473 3218
rect 1494 3192 1497 3248
rect 1526 3232 1529 3278
rect 1534 3272 1537 3318
rect 1646 3282 1649 3318
rect 1686 3312 1689 3318
rect 1710 3292 1713 3328
rect 1734 3322 1737 3328
rect 1682 3278 1686 3281
rect 1646 3272 1649 3278
rect 1694 3272 1697 3278
rect 1578 3268 1582 3271
rect 1666 3268 1670 3271
rect 1542 3262 1545 3268
rect 1566 3262 1569 3268
rect 1638 3262 1641 3268
rect 1582 3252 1585 3258
rect 1562 3248 1566 3251
rect 1658 3248 1662 3251
rect 1618 3238 1622 3241
rect 1558 3232 1561 3238
rect 1686 3192 1689 3268
rect 1718 3262 1721 3278
rect 1742 3271 1745 3318
rect 1738 3268 1745 3271
rect 1738 3258 1742 3261
rect 1694 3252 1697 3258
rect 1722 3248 1726 3251
rect 1458 3148 1462 3151
rect 1446 3122 1449 3128
rect 1470 3112 1473 3148
rect 1478 3112 1481 3168
rect 1490 3148 1494 3151
rect 1534 3142 1537 3148
rect 1514 3138 1518 3141
rect 1514 3128 1518 3131
rect 1454 3082 1457 3098
rect 1510 3092 1513 3118
rect 1526 3082 1529 3138
rect 1534 3092 1537 3128
rect 1550 3122 1553 3148
rect 1582 3142 1585 3148
rect 1578 3138 1582 3141
rect 1590 3132 1593 3158
rect 1634 3148 1638 3151
rect 1582 3112 1585 3118
rect 1594 3088 1601 3091
rect 1422 3072 1425 3078
rect 1302 3062 1305 3068
rect 1382 3062 1385 3068
rect 1414 3062 1417 3068
rect 1438 3062 1441 3068
rect 1318 3058 1326 3061
rect 1310 3052 1313 3058
rect 1318 3052 1321 3058
rect 1446 3052 1449 3058
rect 1394 3048 1398 3051
rect 1326 3042 1329 3048
rect 1214 2992 1217 3038
rect 1230 2992 1233 3018
rect 1368 3003 1370 3007
rect 1374 3003 1377 3007
rect 1381 3003 1384 3007
rect 1430 2972 1433 3038
rect 1462 2992 1465 3068
rect 1478 3052 1481 3068
rect 1490 3066 1494 3069
rect 1534 3062 1537 3068
rect 1542 3052 1545 3078
rect 1550 3072 1553 3088
rect 1598 3072 1601 3088
rect 1614 3062 1617 3138
rect 1622 3122 1625 3138
rect 1630 3052 1633 3108
rect 1646 3092 1649 3178
rect 1718 3162 1721 3168
rect 1658 3158 1662 3161
rect 1742 3152 1745 3158
rect 1750 3152 1753 3258
rect 1766 3251 1769 3278
rect 1778 3258 1782 3261
rect 1786 3258 1790 3261
rect 1762 3248 1769 3251
rect 1778 3248 1782 3251
rect 1758 3242 1761 3248
rect 1798 3242 1801 3338
rect 1838 3332 1841 3348
rect 1894 3342 1897 3348
rect 1862 3332 1865 3338
rect 1818 3328 1822 3331
rect 1872 3303 1874 3307
rect 1878 3303 1881 3307
rect 1885 3303 1888 3307
rect 1830 3282 1833 3298
rect 1810 3258 1814 3261
rect 1806 3162 1809 3218
rect 1830 3152 1833 3278
rect 1838 3272 1841 3278
rect 1886 3262 1889 3268
rect 1838 3252 1841 3258
rect 1870 3242 1873 3248
rect 1670 3132 1673 3148
rect 1694 3142 1697 3148
rect 1710 3142 1713 3148
rect 1730 3140 1734 3143
rect 1742 3142 1745 3148
rect 1766 3142 1769 3148
rect 1782 3142 1785 3148
rect 1806 3142 1809 3148
rect 1862 3142 1865 3158
rect 1870 3152 1873 3178
rect 1918 3172 1921 3318
rect 1926 3292 1929 3348
rect 1950 3321 1953 3338
rect 1950 3318 1958 3321
rect 1982 3282 1985 3318
rect 1998 3291 2001 3338
rect 1994 3288 2001 3291
rect 2006 3322 2009 3348
rect 1990 3272 1993 3288
rect 1926 3182 1929 3258
rect 1934 3252 1937 3268
rect 1966 3252 1969 3258
rect 1982 3252 1985 3268
rect 2006 3261 2009 3318
rect 2022 3292 2025 3328
rect 2038 3312 2041 3318
rect 2046 3292 2049 3338
rect 2054 3332 2057 3338
rect 2002 3258 2009 3261
rect 2034 3288 2038 3291
rect 1998 3242 2001 3248
rect 1926 3162 1929 3178
rect 1942 3152 1945 3158
rect 1958 3142 1961 3148
rect 1966 3142 1969 3168
rect 2014 3142 2017 3288
rect 2054 3262 2057 3278
rect 2062 3262 2065 3348
rect 2078 3282 2081 3338
rect 2086 3292 2089 3368
rect 2098 3348 2102 3351
rect 2110 3342 2113 3358
rect 2126 3332 2129 3358
rect 2138 3348 2142 3351
rect 2078 3272 2081 3278
rect 2022 3252 2025 3258
rect 2042 3248 2046 3251
rect 2086 3242 2089 3248
rect 2094 3152 2097 3318
rect 2126 3272 2129 3328
rect 2150 3292 2153 3358
rect 2158 3332 2161 3338
rect 2166 3292 2169 3348
rect 2190 3342 2193 3488
rect 2198 3452 2201 3478
rect 2214 3462 2217 3488
rect 2326 3482 2329 3518
rect 2306 3478 2310 3481
rect 2362 3478 2366 3481
rect 2222 3472 2225 3478
rect 2358 3472 2361 3478
rect 2306 3468 2310 3471
rect 2230 3452 2233 3468
rect 2278 3452 2281 3468
rect 2286 3462 2289 3468
rect 2294 3452 2297 3458
rect 2350 3452 2353 3458
rect 2322 3448 2326 3451
rect 2198 3352 2201 3448
rect 2206 3382 2209 3428
rect 2206 3342 2209 3378
rect 2174 3332 2177 3338
rect 2186 3328 2190 3331
rect 2194 3288 2198 3291
rect 2114 3268 2118 3271
rect 2102 3252 2105 3268
rect 2114 3258 2118 3261
rect 2142 3252 2145 3278
rect 2174 3242 2177 3248
rect 2098 3148 2105 3151
rect 1906 3138 1910 3141
rect 1710 3112 1713 3128
rect 1750 3101 1753 3118
rect 1782 3112 1785 3128
rect 1814 3121 1817 3138
rect 1814 3118 1822 3121
rect 1742 3098 1753 3101
rect 1830 3102 1833 3118
rect 1872 3103 1874 3107
rect 1878 3103 1881 3107
rect 1885 3103 1888 3107
rect 1658 3088 1662 3091
rect 1742 3072 1745 3098
rect 1754 3088 1758 3091
rect 1854 3082 1857 3098
rect 1998 3092 2001 3118
rect 2022 3102 2025 3138
rect 1986 3088 1990 3091
rect 1990 3072 1993 3078
rect 1654 3052 1657 3068
rect 1718 3052 1721 3058
rect 1726 3052 1729 3068
rect 1790 3052 1793 3058
rect 1474 3048 1478 3051
rect 1522 3038 1526 3041
rect 1470 3032 1473 3038
rect 1474 2988 1478 2991
rect 1578 2988 1582 2991
rect 1342 2962 1345 2968
rect 1222 2942 1225 2958
rect 1406 2951 1409 2958
rect 1294 2942 1297 2947
rect 1198 2938 1206 2941
rect 1158 2912 1161 2928
rect 1198 2892 1201 2938
rect 1098 2888 1102 2891
rect 1226 2888 1230 2891
rect 1286 2882 1289 2938
rect 742 2872 745 2878
rect 918 2872 921 2878
rect 1014 2872 1017 2878
rect 1182 2872 1185 2878
rect 1254 2872 1257 2878
rect 802 2868 806 2871
rect 1378 2868 1382 2871
rect 734 2772 737 2868
rect 774 2792 777 2848
rect 746 2748 750 2751
rect 770 2748 774 2751
rect 710 2742 713 2747
rect 742 2722 745 2728
rect 766 2692 769 2708
rect 782 2692 785 2768
rect 790 2722 793 2868
rect 798 2852 801 2858
rect 822 2792 825 2868
rect 902 2852 905 2859
rect 998 2852 1001 2859
rect 1094 2842 1097 2868
rect 1214 2862 1217 2868
rect 1302 2862 1305 2868
rect 1166 2852 1169 2859
rect 918 2792 921 2838
rect 798 2762 801 2768
rect 850 2758 854 2761
rect 806 2742 809 2758
rect 1118 2752 1121 2758
rect 814 2748 822 2751
rect 898 2748 902 2751
rect 954 2748 958 2751
rect 978 2748 982 2751
rect 1082 2748 1086 2751
rect 814 2732 817 2748
rect 830 2732 833 2738
rect 802 2728 806 2731
rect 814 2692 817 2728
rect 838 2692 841 2738
rect 902 2732 905 2738
rect 866 2718 870 2721
rect 846 2691 849 2718
rect 856 2703 858 2707
rect 862 2703 865 2707
rect 869 2703 872 2707
rect 894 2692 897 2698
rect 846 2688 854 2691
rect 658 2678 662 2681
rect 738 2678 742 2681
rect 646 2652 649 2678
rect 822 2672 825 2678
rect 894 2672 897 2688
rect 926 2682 929 2718
rect 934 2692 937 2708
rect 950 2692 953 2738
rect 962 2728 966 2731
rect 982 2722 985 2728
rect 842 2668 846 2671
rect 614 2532 617 2558
rect 626 2548 630 2551
rect 638 2542 641 2558
rect 622 2472 625 2508
rect 646 2492 649 2628
rect 662 2592 665 2668
rect 670 2662 673 2668
rect 718 2662 721 2668
rect 694 2592 697 2658
rect 742 2652 745 2668
rect 742 2602 745 2648
rect 798 2602 801 2668
rect 806 2652 809 2658
rect 718 2592 721 2598
rect 790 2582 793 2588
rect 738 2578 742 2581
rect 758 2572 761 2578
rect 798 2572 801 2598
rect 822 2592 825 2668
rect 918 2662 921 2668
rect 942 2662 945 2668
rect 974 2662 977 2718
rect 990 2671 993 2718
rect 998 2702 1001 2748
rect 1006 2692 1009 2698
rect 1002 2678 1006 2681
rect 1022 2672 1025 2738
rect 1086 2692 1089 2738
rect 1094 2692 1097 2728
rect 1042 2688 1046 2691
rect 1110 2682 1113 2748
rect 1158 2742 1161 2748
rect 1118 2732 1121 2738
rect 1138 2728 1142 2731
rect 1118 2692 1121 2718
rect 1158 2712 1161 2728
rect 1166 2722 1169 2728
rect 1058 2678 1062 2681
rect 1158 2672 1161 2678
rect 1166 2672 1169 2718
rect 1174 2681 1177 2818
rect 1182 2752 1185 2758
rect 1190 2742 1193 2758
rect 1198 2752 1201 2848
rect 1230 2792 1233 2858
rect 1186 2738 1190 2741
rect 1182 2692 1185 2708
rect 1198 2692 1201 2748
rect 1206 2742 1209 2758
rect 1246 2752 1249 2758
rect 1226 2748 1230 2751
rect 1210 2738 1214 2741
rect 1250 2738 1254 2741
rect 1222 2721 1225 2738
rect 1262 2732 1265 2748
rect 1270 2732 1273 2738
rect 1222 2718 1230 2721
rect 1262 2712 1265 2728
rect 1174 2678 1185 2681
rect 990 2668 1001 2671
rect 1034 2668 1038 2671
rect 1082 2668 1086 2671
rect 954 2658 958 2661
rect 986 2658 990 2661
rect 830 2652 833 2658
rect 886 2632 889 2658
rect 846 2592 849 2598
rect 894 2592 897 2658
rect 670 2552 673 2558
rect 654 2502 657 2538
rect 678 2532 681 2558
rect 686 2492 689 2538
rect 702 2512 705 2548
rect 710 2542 713 2568
rect 742 2562 745 2568
rect 778 2558 782 2561
rect 858 2558 862 2561
rect 770 2548 774 2551
rect 786 2548 793 2551
rect 742 2532 745 2538
rect 730 2528 737 2531
rect 734 2492 737 2528
rect 766 2492 769 2508
rect 630 2472 633 2488
rect 738 2478 742 2481
rect 574 2462 577 2468
rect 678 2462 681 2468
rect 714 2458 718 2461
rect 690 2438 694 2441
rect 638 2392 641 2438
rect 678 2392 681 2428
rect 594 2368 598 2371
rect 626 2368 630 2371
rect 674 2368 678 2371
rect 614 2352 617 2358
rect 646 2352 649 2358
rect 634 2348 638 2351
rect 638 2342 641 2348
rect 654 2342 657 2358
rect 662 2352 665 2368
rect 694 2352 697 2358
rect 702 2352 705 2458
rect 714 2448 718 2451
rect 726 2442 729 2468
rect 734 2452 737 2478
rect 774 2472 777 2478
rect 750 2452 753 2458
rect 714 2368 718 2371
rect 750 2362 753 2448
rect 758 2432 761 2468
rect 782 2452 785 2538
rect 790 2532 793 2548
rect 806 2542 809 2558
rect 858 2548 862 2551
rect 898 2548 902 2551
rect 806 2532 809 2538
rect 790 2492 793 2528
rect 814 2492 817 2548
rect 906 2538 910 2541
rect 838 2532 841 2538
rect 830 2492 833 2528
rect 856 2503 858 2507
rect 862 2503 865 2507
rect 869 2503 872 2507
rect 910 2492 913 2528
rect 854 2482 857 2488
rect 778 2448 782 2451
rect 790 2432 793 2458
rect 798 2442 801 2468
rect 802 2438 806 2441
rect 814 2432 817 2478
rect 838 2472 841 2478
rect 898 2468 902 2471
rect 822 2442 825 2448
rect 770 2388 774 2391
rect 786 2368 790 2371
rect 766 2362 769 2368
rect 742 2352 745 2358
rect 750 2352 753 2358
rect 682 2338 686 2341
rect 534 2332 537 2338
rect 582 2321 585 2338
rect 578 2318 585 2321
rect 590 2312 593 2328
rect 614 2322 617 2328
rect 630 2292 633 2328
rect 678 2322 681 2338
rect 694 2312 697 2348
rect 726 2332 729 2348
rect 738 2338 742 2341
rect 758 2332 761 2358
rect 778 2348 782 2351
rect 798 2342 801 2378
rect 830 2362 833 2418
rect 838 2392 841 2468
rect 862 2372 865 2458
rect 902 2452 905 2468
rect 890 2448 894 2451
rect 918 2442 921 2658
rect 998 2652 1001 2668
rect 1054 2662 1057 2668
rect 966 2642 969 2648
rect 954 2628 958 2631
rect 950 2542 953 2578
rect 966 2532 969 2628
rect 1006 2592 1009 2608
rect 1022 2592 1025 2658
rect 982 2552 985 2558
rect 990 2542 993 2548
rect 966 2492 969 2518
rect 954 2478 958 2481
rect 934 2472 937 2478
rect 818 2348 822 2351
rect 730 2328 734 2331
rect 806 2312 809 2348
rect 894 2342 897 2438
rect 926 2422 929 2458
rect 934 2382 937 2468
rect 942 2442 945 2448
rect 910 2351 913 2358
rect 958 2352 961 2428
rect 974 2352 977 2538
rect 998 2522 1001 2558
rect 998 2392 1001 2518
rect 1014 2442 1017 2528
rect 1022 2522 1025 2528
rect 1038 2522 1041 2648
rect 1046 2552 1049 2658
rect 1062 2652 1065 2668
rect 1110 2662 1113 2668
rect 1082 2658 1086 2661
rect 1098 2648 1105 2651
rect 1062 2552 1065 2648
rect 1078 2592 1081 2608
rect 1102 2592 1105 2648
rect 1110 2612 1113 2658
rect 1118 2632 1121 2668
rect 1134 2642 1137 2658
rect 1142 2652 1145 2658
rect 1126 2611 1129 2618
rect 1126 2608 1134 2611
rect 1182 2592 1185 2678
rect 1254 2672 1257 2678
rect 1218 2668 1222 2671
rect 1242 2668 1246 2671
rect 1218 2658 1222 2661
rect 1230 2652 1233 2668
rect 1254 2662 1257 2668
rect 1262 2662 1265 2668
rect 1198 2641 1201 2648
rect 1206 2641 1209 2648
rect 1198 2638 1209 2641
rect 1078 2582 1081 2588
rect 1102 2562 1105 2588
rect 1198 2582 1201 2588
rect 1110 2572 1113 2578
rect 1066 2548 1078 2551
rect 1074 2538 1078 2541
rect 1054 2532 1057 2538
rect 1086 2512 1089 2558
rect 1094 2542 1097 2558
rect 1094 2492 1097 2538
rect 1102 2512 1105 2548
rect 1206 2542 1209 2638
rect 1214 2592 1217 2618
rect 1246 2592 1249 2658
rect 1270 2632 1273 2658
rect 1278 2622 1281 2858
rect 1318 2842 1321 2868
rect 1390 2862 1393 2938
rect 1438 2932 1441 2938
rect 1454 2932 1457 2968
rect 1570 2958 1574 2961
rect 1726 2952 1729 3048
rect 1822 3042 1825 3059
rect 1870 3042 1873 3058
rect 1902 3052 1905 3068
rect 1918 3052 1921 3059
rect 2006 3052 2009 3068
rect 2022 3062 2025 3078
rect 2038 3052 2041 3118
rect 2078 3102 2081 3128
rect 2094 3122 2097 3138
rect 2046 3052 2049 3058
rect 2054 3052 2057 3058
rect 2062 3052 2065 3078
rect 2086 3072 2089 3118
rect 2094 3072 2097 3098
rect 2086 3062 2089 3068
rect 2102 3062 2105 3148
rect 2150 3142 2153 3218
rect 2158 3152 2161 3158
rect 2174 3132 2177 3168
rect 2206 3162 2209 3338
rect 2238 3302 2241 3318
rect 2234 3288 2238 3291
rect 2222 3282 2225 3288
rect 2254 3272 2257 3448
rect 2334 3442 2337 3448
rect 2374 3441 2377 3528
rect 2422 3512 2425 3518
rect 2394 3468 2398 3471
rect 2406 3462 2409 3468
rect 2382 3452 2385 3458
rect 2454 3451 2457 3518
rect 2470 3502 2473 3548
rect 2486 3542 2489 3548
rect 2534 3542 2537 3568
rect 2550 3562 2553 3568
rect 2590 3562 2593 3568
rect 2654 3562 2657 3568
rect 2686 3562 2689 3578
rect 2594 3558 2601 3561
rect 2610 3558 2614 3561
rect 2634 3558 2638 3561
rect 2694 3561 2697 3668
rect 2742 3662 2745 3668
rect 2726 3582 2729 3618
rect 2742 3572 2745 3658
rect 2838 3652 2841 3659
rect 2854 3642 2857 3668
rect 2910 3662 2913 3668
rect 3062 3663 3065 3678
rect 3118 3672 3121 3678
rect 2870 3652 2873 3658
rect 2902 3652 2905 3658
rect 2778 3628 2782 3631
rect 2966 3622 2969 3658
rect 2990 3612 2993 3658
rect 3078 3642 3081 3668
rect 3110 3662 3113 3668
rect 3214 3662 3217 3678
rect 3326 3672 3329 3678
rect 3726 3672 3729 3678
rect 3738 3668 3742 3671
rect 3002 3618 3006 3621
rect 2706 3568 2718 3571
rect 2694 3558 2705 3561
rect 2586 3548 2590 3551
rect 2562 3538 2566 3541
rect 2486 3512 2489 3528
rect 2510 3522 2513 3538
rect 2534 3532 2537 3538
rect 2542 3532 2545 3538
rect 2462 3472 2465 3478
rect 2494 3472 2497 3508
rect 2466 3458 2470 3461
rect 2454 3448 2462 3451
rect 2374 3438 2385 3441
rect 2322 3418 2326 3421
rect 2318 3382 2321 3388
rect 2278 3352 2281 3378
rect 2350 3372 2353 3418
rect 2382 3372 2385 3438
rect 2392 3403 2394 3407
rect 2398 3403 2401 3407
rect 2405 3403 2408 3407
rect 2330 3368 2334 3371
rect 2318 3362 2321 3368
rect 2342 3352 2345 3358
rect 2290 3338 2294 3341
rect 2302 3332 2305 3348
rect 2318 3332 2321 3348
rect 2350 3342 2353 3368
rect 2298 3328 2302 3331
rect 2362 3328 2366 3331
rect 2318 3322 2321 3328
rect 2262 3292 2265 3318
rect 2358 3312 2361 3318
rect 2270 3282 2273 3288
rect 2226 3268 2238 3271
rect 2234 3258 2238 3261
rect 2214 3252 2217 3258
rect 2254 3152 2257 3268
rect 2302 3262 2305 3288
rect 2310 3272 2313 3308
rect 2282 3258 2286 3261
rect 2318 3252 2321 3278
rect 2330 3258 2342 3261
rect 2282 3248 2286 3251
rect 2330 3248 2334 3251
rect 2350 3242 2353 3248
rect 2170 3128 2174 3131
rect 2210 3118 2214 3121
rect 2106 3048 2110 3051
rect 1790 2962 1793 2968
rect 1814 2962 1817 2968
rect 1806 2952 1809 2958
rect 1838 2952 1841 3038
rect 1862 2972 1865 3018
rect 1846 2962 1849 2968
rect 1846 2952 1849 2958
rect 1286 2692 1289 2828
rect 1318 2732 1321 2838
rect 1326 2792 1329 2858
rect 1368 2803 1370 2807
rect 1374 2803 1377 2807
rect 1381 2803 1384 2807
rect 1354 2788 1358 2791
rect 1398 2692 1401 2918
rect 1410 2888 1414 2891
rect 1438 2862 1441 2868
rect 1446 2862 1449 2928
rect 1454 2762 1457 2928
rect 1502 2872 1505 2948
rect 1510 2892 1513 2948
rect 1550 2942 1553 2948
rect 1614 2942 1617 2948
rect 1646 2942 1649 2947
rect 1710 2942 1713 2948
rect 1862 2942 1865 2958
rect 1902 2952 1905 3038
rect 2038 3032 2041 3038
rect 1998 3022 2001 3028
rect 2014 2972 2017 3018
rect 1954 2958 1958 2961
rect 1858 2938 1862 2941
rect 1774 2932 1777 2938
rect 1526 2882 1529 2898
rect 1574 2892 1577 2928
rect 1598 2888 1606 2891
rect 1542 2872 1545 2888
rect 1598 2872 1601 2888
rect 1586 2868 1590 2871
rect 1470 2822 1473 2859
rect 1502 2852 1505 2858
rect 1422 2711 1425 2747
rect 1438 2742 1441 2748
rect 1454 2742 1457 2748
rect 1422 2708 1433 2711
rect 1302 2662 1305 2688
rect 1326 2682 1329 2688
rect 1370 2668 1374 2671
rect 1342 2662 1345 2668
rect 1290 2648 1294 2651
rect 1310 2642 1313 2648
rect 1302 2632 1305 2638
rect 1310 2592 1313 2618
rect 1342 2592 1345 2658
rect 1358 2652 1361 2668
rect 1370 2648 1374 2651
rect 1350 2592 1353 2638
rect 1106 2488 1113 2491
rect 1110 2472 1113 2488
rect 1126 2482 1129 2538
rect 1174 2521 1177 2538
rect 1170 2518 1177 2521
rect 1190 2522 1193 2528
rect 1158 2502 1161 2518
rect 1134 2472 1137 2488
rect 1150 2482 1153 2498
rect 1174 2492 1177 2508
rect 1206 2492 1209 2538
rect 1254 2492 1257 2528
rect 1278 2512 1281 2547
rect 1294 2542 1297 2548
rect 1326 2532 1329 2538
rect 1318 2521 1321 2528
rect 1318 2518 1329 2521
rect 1214 2488 1222 2491
rect 1202 2478 1206 2481
rect 1030 2392 1033 2459
rect 1010 2368 1014 2371
rect 1026 2368 1030 2371
rect 946 2348 950 2351
rect 962 2348 966 2351
rect 970 2338 974 2341
rect 666 2288 670 2291
rect 478 2278 489 2281
rect 382 2272 385 2278
rect 486 2272 489 2278
rect 730 2279 737 2281
rect 726 2278 737 2279
rect 754 2279 761 2281
rect 750 2278 761 2279
rect 542 2272 545 2278
rect 654 2272 657 2278
rect 94 2268 102 2271
rect 338 2268 342 2271
rect 426 2268 430 2271
rect 562 2268 566 2271
rect 102 2262 105 2268
rect 110 2262 113 2268
rect 6 2152 9 2198
rect 158 2182 161 2268
rect 238 2262 241 2268
rect 170 2258 174 2261
rect 314 2258 318 2261
rect 190 2252 193 2258
rect 210 2248 214 2251
rect 366 2242 369 2258
rect 326 2192 329 2228
rect 344 2203 346 2207
rect 350 2203 353 2207
rect 357 2203 360 2207
rect 366 2192 369 2218
rect 374 2212 377 2268
rect 478 2262 481 2268
rect 426 2258 430 2261
rect 450 2258 454 2261
rect 402 2248 406 2251
rect 414 2172 417 2238
rect 534 2232 537 2268
rect 542 2222 545 2268
rect 598 2262 601 2268
rect 554 2258 558 2261
rect 590 2252 593 2258
rect 646 2252 649 2268
rect 710 2262 713 2278
rect 734 2262 737 2278
rect 758 2262 761 2278
rect 766 2262 769 2308
rect 856 2303 858 2307
rect 862 2303 865 2307
rect 869 2303 872 2307
rect 790 2292 793 2298
rect 886 2272 889 2338
rect 894 2292 897 2338
rect 926 2322 929 2338
rect 982 2332 985 2368
rect 998 2352 1001 2358
rect 954 2328 958 2331
rect 970 2288 977 2291
rect 926 2272 929 2278
rect 974 2272 977 2288
rect 982 2272 985 2308
rect 678 2242 681 2248
rect 554 2238 558 2241
rect 566 2192 569 2208
rect 486 2182 489 2188
rect 154 2168 158 2171
rect 170 2168 174 2171
rect 54 2162 57 2168
rect 66 2158 70 2161
rect 106 2148 110 2151
rect 30 2112 33 2128
rect 46 2112 49 2148
rect 74 2138 78 2141
rect 106 2138 110 2141
rect 54 2132 57 2138
rect 94 2132 97 2138
rect 126 2132 129 2168
rect 178 2158 182 2161
rect 134 2152 137 2158
rect 158 2152 161 2158
rect 202 2148 206 2151
rect 114 2128 118 2131
rect 6 2088 14 2091
rect 6 2072 9 2088
rect 22 2061 25 2108
rect 30 2092 33 2098
rect 70 2092 73 2128
rect 38 2088 46 2091
rect 38 2072 41 2088
rect 78 2082 81 2128
rect 86 2082 89 2118
rect 110 2092 113 2108
rect 134 2102 137 2148
rect 142 2142 145 2148
rect 174 2102 177 2128
rect 166 2098 174 2101
rect 62 2062 65 2068
rect 18 2058 30 2061
rect 6 1972 9 1978
rect 14 1932 17 2018
rect 14 1902 17 1928
rect 22 1892 25 2058
rect 78 2052 81 2078
rect 34 2048 38 2051
rect 86 1982 89 2068
rect 134 2042 137 2068
rect 142 2041 145 2078
rect 150 2062 153 2068
rect 158 2062 161 2068
rect 166 2052 169 2098
rect 190 2082 193 2138
rect 206 2132 209 2138
rect 214 2132 217 2158
rect 174 2062 177 2078
rect 206 2062 209 2078
rect 214 2052 217 2128
rect 230 2092 233 2118
rect 238 2092 241 2138
rect 262 2132 265 2148
rect 246 2082 249 2118
rect 270 2112 273 2138
rect 278 2132 281 2168
rect 394 2158 398 2161
rect 390 2152 393 2158
rect 290 2138 294 2141
rect 346 2138 350 2141
rect 366 2132 369 2148
rect 382 2142 385 2148
rect 254 2082 257 2088
rect 318 2082 321 2108
rect 342 2092 345 2128
rect 350 2082 353 2118
rect 406 2112 409 2148
rect 414 2142 417 2168
rect 454 2162 457 2178
rect 462 2172 465 2178
rect 470 2158 478 2161
rect 422 2152 425 2158
rect 374 2082 377 2098
rect 422 2092 425 2148
rect 438 2142 441 2158
rect 450 2148 454 2151
rect 438 2132 441 2138
rect 438 2102 441 2128
rect 402 2088 406 2091
rect 430 2082 433 2088
rect 438 2072 441 2078
rect 454 2072 457 2088
rect 470 2082 473 2158
rect 478 2142 481 2158
rect 534 2152 537 2178
rect 618 2158 622 2161
rect 522 2148 526 2151
rect 534 2142 537 2148
rect 558 2142 561 2148
rect 582 2142 585 2158
rect 638 2152 641 2178
rect 662 2172 665 2178
rect 674 2168 678 2171
rect 686 2162 689 2168
rect 658 2158 662 2161
rect 602 2148 606 2151
rect 618 2148 622 2151
rect 646 2142 649 2148
rect 594 2138 598 2141
rect 542 2132 545 2138
rect 494 2112 497 2118
rect 482 2088 486 2091
rect 542 2072 545 2108
rect 566 2092 569 2128
rect 606 2122 609 2138
rect 662 2132 665 2148
rect 694 2141 697 2178
rect 758 2171 761 2248
rect 798 2232 801 2268
rect 854 2232 857 2259
rect 766 2182 769 2188
rect 758 2168 769 2171
rect 742 2162 745 2168
rect 758 2152 761 2158
rect 690 2138 697 2141
rect 718 2148 726 2151
rect 702 2142 705 2148
rect 622 2092 625 2118
rect 710 2112 713 2128
rect 718 2092 721 2148
rect 726 2122 729 2138
rect 582 2082 585 2088
rect 570 2078 582 2081
rect 266 2068 270 2071
rect 246 2062 249 2068
rect 274 2058 278 2061
rect 290 2058 294 2061
rect 402 2058 409 2061
rect 290 2048 294 2051
rect 222 2042 225 2048
rect 230 2042 233 2048
rect 302 2042 305 2058
rect 318 2052 321 2058
rect 142 2038 150 2041
rect 162 2038 166 2041
rect 394 2038 398 2041
rect 30 1972 33 1978
rect 38 1972 41 1978
rect 30 1932 33 1968
rect 50 1958 54 1961
rect 78 1952 81 1958
rect 86 1952 89 1978
rect 58 1948 62 1951
rect 98 1948 102 1951
rect 38 1942 41 1948
rect 78 1942 81 1948
rect 110 1942 113 2038
rect 174 1992 177 2028
rect 206 1992 209 2018
rect 254 1982 257 2018
rect 138 1968 145 1971
rect 134 1962 137 1968
rect 142 1962 145 1968
rect 214 1962 217 1978
rect 226 1968 230 1971
rect 242 1968 246 1971
rect 266 1968 270 1971
rect 294 1961 297 2018
rect 406 2012 409 2058
rect 414 2052 417 2068
rect 450 2058 454 2061
rect 422 2042 425 2048
rect 470 2032 473 2038
rect 494 2022 497 2058
rect 344 2003 346 2007
rect 350 2003 353 2007
rect 357 2003 360 2007
rect 398 1992 401 1998
rect 286 1958 297 1961
rect 66 1938 70 1941
rect 50 1928 54 1931
rect 82 1928 86 1931
rect 6 1888 14 1891
rect 6 1872 9 1888
rect 62 1882 65 1898
rect 70 1892 73 1928
rect 54 1841 57 1868
rect 62 1852 65 1878
rect 110 1872 113 1878
rect 122 1868 126 1871
rect 46 1838 57 1841
rect 78 1842 81 1868
rect 106 1858 110 1861
rect 38 1792 41 1838
rect 6 1772 9 1778
rect 14 1732 17 1778
rect 26 1768 30 1771
rect 30 1762 33 1768
rect 38 1752 41 1768
rect 46 1692 49 1838
rect 78 1792 81 1838
rect 86 1792 89 1858
rect 142 1852 145 1958
rect 262 1952 265 1958
rect 158 1892 161 1908
rect 166 1872 169 1898
rect 190 1892 193 1938
rect 206 1922 209 1938
rect 214 1932 217 1938
rect 222 1922 225 1928
rect 182 1862 185 1868
rect 114 1848 118 1851
rect 98 1838 102 1841
rect 122 1788 126 1791
rect 70 1762 73 1778
rect 90 1768 94 1771
rect 138 1768 142 1771
rect 78 1752 81 1768
rect 98 1758 102 1761
rect 86 1748 94 1751
rect 122 1748 126 1751
rect 54 1738 62 1741
rect 46 1662 49 1688
rect 54 1672 57 1738
rect 62 1732 65 1738
rect 86 1692 89 1748
rect 130 1738 134 1741
rect 142 1732 145 1748
rect 150 1742 153 1818
rect 158 1792 161 1848
rect 182 1832 185 1858
rect 198 1852 201 1898
rect 206 1852 209 1918
rect 238 1902 241 1918
rect 254 1912 257 1948
rect 286 1942 289 1958
rect 302 1952 305 1958
rect 318 1952 321 1958
rect 294 1942 297 1948
rect 326 1942 329 1948
rect 266 1928 270 1931
rect 310 1922 313 1938
rect 334 1892 337 1938
rect 342 1912 345 1948
rect 214 1862 217 1868
rect 206 1842 209 1848
rect 222 1842 225 1878
rect 238 1872 241 1888
rect 334 1882 337 1888
rect 342 1882 345 1908
rect 270 1872 273 1878
rect 302 1872 305 1878
rect 326 1872 329 1878
rect 290 1868 294 1871
rect 198 1792 201 1838
rect 214 1832 217 1838
rect 174 1772 177 1778
rect 238 1742 241 1868
rect 254 1862 257 1868
rect 350 1862 353 1948
rect 358 1912 361 1958
rect 390 1952 393 1958
rect 370 1948 374 1951
rect 382 1942 385 1948
rect 398 1941 401 1968
rect 394 1938 401 1941
rect 358 1872 361 1908
rect 406 1892 409 2008
rect 446 1962 449 1968
rect 438 1932 441 1958
rect 430 1922 433 1928
rect 454 1892 457 2018
rect 470 1992 473 2018
rect 502 2002 505 2068
rect 514 2058 518 2061
rect 514 2048 518 2051
rect 526 2012 529 2058
rect 566 2052 569 2078
rect 586 2068 590 2071
rect 578 2048 582 2051
rect 638 2051 641 2068
rect 646 2062 649 2078
rect 742 2072 745 2108
rect 766 2092 769 2168
rect 774 2152 777 2188
rect 782 2152 785 2158
rect 774 2132 777 2148
rect 798 2132 801 2228
rect 886 2192 889 2248
rect 826 2148 830 2151
rect 806 2142 809 2148
rect 854 2142 857 2148
rect 878 2142 881 2158
rect 918 2152 921 2268
rect 926 2182 929 2268
rect 990 2262 993 2308
rect 998 2272 1001 2348
rect 1006 2342 1009 2348
rect 1006 2252 1009 2328
rect 1014 2292 1017 2358
rect 1030 2312 1033 2348
rect 1038 2332 1041 2398
rect 1046 2322 1049 2468
rect 1062 2382 1065 2468
rect 1122 2458 1126 2461
rect 1110 2392 1113 2458
rect 1142 2452 1145 2478
rect 1214 2472 1217 2488
rect 1246 2482 1249 2488
rect 1302 2482 1305 2488
rect 1294 2472 1297 2478
rect 1162 2458 1166 2461
rect 1174 2452 1177 2468
rect 1246 2462 1249 2468
rect 1294 2462 1297 2468
rect 1318 2462 1321 2498
rect 1210 2458 1214 2461
rect 1266 2458 1270 2461
rect 1234 2448 1238 2451
rect 1174 2442 1177 2448
rect 1206 2442 1209 2448
rect 1278 2442 1281 2448
rect 1294 2442 1297 2448
rect 1126 2402 1129 2418
rect 1098 2378 1102 2381
rect 1118 2372 1121 2378
rect 1126 2362 1129 2398
rect 1294 2391 1297 2438
rect 1326 2422 1329 2518
rect 1334 2472 1337 2488
rect 1350 2482 1353 2498
rect 1358 2472 1361 2648
rect 1430 2622 1433 2708
rect 1368 2603 1370 2607
rect 1374 2603 1377 2607
rect 1381 2603 1384 2607
rect 1390 2511 1393 2548
rect 1382 2508 1393 2511
rect 1382 2492 1385 2508
rect 1382 2432 1385 2438
rect 1290 2388 1297 2391
rect 1186 2368 1190 2371
rect 1082 2358 1086 2361
rect 1062 2352 1065 2358
rect 1170 2348 1174 2351
rect 1078 2342 1081 2348
rect 1126 2342 1129 2348
rect 1058 2338 1062 2341
rect 1102 2332 1105 2338
rect 1034 2288 1038 2291
rect 1030 2252 1033 2268
rect 1014 2242 1017 2248
rect 894 2142 897 2148
rect 910 2142 913 2148
rect 926 2142 929 2158
rect 950 2152 953 2178
rect 990 2152 993 2218
rect 938 2148 942 2151
rect 782 2091 785 2128
rect 774 2088 785 2091
rect 830 2092 833 2138
rect 858 2128 862 2131
rect 838 2112 841 2128
rect 902 2121 905 2138
rect 942 2132 945 2138
rect 902 2118 910 2121
rect 856 2103 858 2107
rect 862 2103 865 2107
rect 869 2103 872 2107
rect 850 2088 857 2091
rect 774 2078 777 2088
rect 806 2072 809 2078
rect 854 2072 857 2088
rect 878 2088 886 2091
rect 878 2072 881 2088
rect 694 2062 697 2068
rect 638 2048 649 2051
rect 462 1972 465 1988
rect 474 1958 478 1961
rect 470 1932 473 1948
rect 494 1942 497 1988
rect 502 1892 505 1988
rect 574 1972 577 1998
rect 646 1992 649 2048
rect 694 2032 697 2058
rect 534 1962 537 1968
rect 582 1962 585 1968
rect 638 1962 641 1968
rect 522 1958 526 1961
rect 570 1948 574 1951
rect 594 1948 598 1951
rect 518 1942 521 1948
rect 594 1938 598 1941
rect 510 1932 513 1938
rect 534 1892 537 1938
rect 614 1932 617 1948
rect 390 1888 398 1891
rect 382 1882 385 1888
rect 370 1878 374 1881
rect 390 1872 393 1888
rect 550 1882 553 1928
rect 598 1922 601 1928
rect 630 1922 633 1958
rect 726 1951 729 1988
rect 638 1942 641 1948
rect 742 1942 745 2038
rect 758 1992 761 2028
rect 650 1938 654 1941
rect 662 1912 665 1918
rect 562 1878 566 1881
rect 526 1872 529 1878
rect 466 1868 470 1871
rect 438 1862 441 1868
rect 246 1842 249 1858
rect 262 1852 265 1858
rect 286 1852 289 1858
rect 326 1852 329 1858
rect 274 1848 278 1851
rect 350 1842 353 1858
rect 344 1803 346 1807
rect 350 1803 353 1807
rect 357 1803 360 1807
rect 330 1788 334 1791
rect 394 1768 398 1771
rect 418 1768 422 1771
rect 182 1732 185 1738
rect 142 1692 145 1728
rect 198 1692 201 1708
rect 222 1692 225 1718
rect 238 1712 241 1728
rect 254 1712 257 1748
rect 262 1742 265 1758
rect 278 1742 281 1768
rect 286 1762 289 1768
rect 294 1752 297 1768
rect 314 1758 318 1761
rect 386 1758 390 1761
rect 286 1742 289 1748
rect 334 1742 337 1748
rect 342 1722 345 1738
rect 210 1688 217 1691
rect 110 1672 113 1678
rect 166 1672 169 1678
rect 214 1672 217 1688
rect 22 1622 25 1658
rect 50 1548 54 1551
rect 10 1538 14 1541
rect 6 1512 9 1528
rect 22 1522 25 1538
rect 38 1522 41 1548
rect 6 1462 9 1478
rect 38 1472 41 1498
rect 46 1452 49 1458
rect 22 1422 25 1428
rect 46 1412 49 1448
rect 22 1392 25 1408
rect 42 1368 46 1371
rect 6 1288 14 1291
rect 6 1272 9 1288
rect 22 1272 25 1348
rect 30 1321 33 1368
rect 54 1362 57 1548
rect 62 1542 65 1558
rect 78 1542 81 1558
rect 86 1552 89 1568
rect 102 1512 105 1668
rect 158 1632 161 1668
rect 238 1652 241 1658
rect 110 1582 113 1588
rect 130 1568 134 1571
rect 158 1562 161 1588
rect 130 1548 137 1551
rect 110 1532 113 1538
rect 118 1521 121 1538
rect 134 1522 137 1548
rect 158 1532 161 1558
rect 118 1518 126 1521
rect 70 1472 73 1478
rect 94 1462 97 1488
rect 102 1462 105 1468
rect 138 1458 142 1461
rect 70 1452 73 1458
rect 70 1392 73 1448
rect 94 1382 97 1418
rect 62 1372 65 1378
rect 102 1371 105 1458
rect 126 1401 129 1449
rect 126 1398 137 1401
rect 94 1368 105 1371
rect 42 1358 46 1361
rect 38 1332 41 1358
rect 62 1332 65 1368
rect 82 1358 86 1361
rect 94 1352 97 1368
rect 110 1352 113 1358
rect 70 1342 73 1348
rect 98 1338 102 1341
rect 30 1318 41 1321
rect 38 1292 41 1318
rect 70 1292 73 1338
rect 82 1328 86 1331
rect 110 1321 113 1348
rect 118 1332 121 1378
rect 110 1318 121 1321
rect 102 1288 110 1291
rect 94 1272 97 1278
rect 102 1272 105 1288
rect 118 1282 121 1318
rect 118 1272 121 1278
rect 126 1272 129 1388
rect 134 1362 137 1398
rect 158 1392 161 1508
rect 166 1482 169 1648
rect 246 1612 249 1668
rect 262 1662 265 1718
rect 310 1681 313 1718
rect 366 1712 369 1748
rect 374 1742 377 1748
rect 398 1732 401 1758
rect 446 1752 449 1868
rect 466 1848 473 1851
rect 470 1792 473 1848
rect 518 1792 521 1868
rect 654 1862 657 1868
rect 550 1852 553 1858
rect 638 1852 641 1859
rect 546 1848 550 1851
rect 574 1782 577 1818
rect 582 1792 585 1838
rect 670 1792 673 1868
rect 726 1862 729 1928
rect 774 1882 777 1948
rect 782 1942 785 1948
rect 462 1762 465 1768
rect 438 1742 441 1748
rect 426 1738 430 1741
rect 406 1732 409 1738
rect 454 1732 457 1758
rect 550 1742 553 1768
rect 686 1752 689 1818
rect 702 1752 705 1798
rect 726 1782 729 1848
rect 742 1822 745 1868
rect 734 1761 737 1808
rect 750 1782 753 1878
rect 726 1758 737 1761
rect 742 1762 745 1778
rect 726 1742 729 1758
rect 758 1752 761 1788
rect 766 1752 769 1818
rect 774 1752 777 1878
rect 782 1872 785 1918
rect 790 1822 793 1858
rect 798 1832 801 2068
rect 898 2058 902 2061
rect 926 2012 929 2068
rect 934 1972 937 2018
rect 942 1982 945 2128
rect 994 2118 998 2121
rect 1046 2112 1049 2318
rect 1054 2312 1057 2328
rect 1150 2312 1153 2348
rect 1162 2338 1166 2341
rect 1182 2332 1185 2338
rect 1130 2288 1134 2291
rect 1118 2272 1121 2278
rect 1166 2272 1169 2278
rect 1102 2252 1105 2259
rect 1182 2222 1185 2328
rect 1198 2282 1201 2338
rect 1254 2292 1257 2347
rect 1270 2342 1273 2348
rect 1278 2272 1281 2308
rect 1318 2292 1321 2378
rect 1342 2302 1345 2348
rect 1350 2342 1353 2428
rect 1422 2412 1425 2547
rect 1438 2542 1441 2658
rect 1454 2592 1457 2708
rect 1494 2692 1497 2758
rect 1462 2602 1465 2659
rect 1502 2592 1505 2848
rect 1518 2732 1521 2738
rect 1526 2692 1529 2868
rect 1562 2858 1566 2861
rect 1610 2858 1614 2861
rect 1626 2848 1630 2851
rect 1558 2842 1561 2848
rect 1638 2842 1641 2868
rect 1646 2862 1649 2888
rect 1654 2852 1657 2878
rect 1662 2872 1665 2878
rect 1678 2872 1681 2888
rect 1790 2882 1793 2928
rect 1798 2892 1801 2918
rect 1694 2862 1697 2878
rect 1714 2868 1718 2871
rect 1666 2858 1670 2861
rect 1722 2858 1726 2861
rect 1734 2852 1737 2868
rect 1542 2772 1545 2818
rect 1582 2762 1585 2838
rect 1606 2752 1609 2818
rect 1646 2802 1649 2818
rect 1654 2792 1657 2828
rect 1678 2792 1681 2848
rect 1742 2832 1745 2878
rect 1806 2872 1809 2918
rect 1806 2862 1809 2868
rect 1822 2862 1825 2938
rect 1838 2921 1841 2938
rect 1834 2918 1841 2921
rect 1846 2872 1849 2918
rect 1872 2903 1874 2907
rect 1878 2903 1881 2907
rect 1885 2903 1888 2907
rect 1866 2888 1870 2891
rect 1894 2882 1897 2938
rect 1910 2902 1913 2938
rect 1918 2932 1921 2938
rect 1926 2922 1929 2948
rect 1942 2932 1945 2958
rect 1974 2952 1977 2968
rect 2006 2952 2009 2958
rect 2022 2952 2025 2998
rect 2030 2972 2033 3018
rect 2034 2958 2038 2961
rect 2034 2948 2038 2951
rect 1950 2942 1953 2948
rect 1982 2942 1985 2948
rect 2002 2928 2009 2931
rect 1990 2922 1993 2928
rect 1950 2892 1953 2918
rect 2006 2892 2009 2928
rect 2038 2892 2041 2938
rect 2046 2932 2049 2948
rect 2054 2892 2057 3048
rect 2118 3042 2121 3118
rect 2230 3112 2233 3138
rect 2262 3132 2265 3148
rect 2226 3078 2230 3081
rect 2126 3072 2129 3078
rect 2182 3072 2185 3078
rect 2246 3062 2249 3108
rect 2270 3072 2273 3188
rect 2294 3132 2297 3158
rect 2302 3142 2305 3218
rect 2342 3162 2345 3218
rect 2318 3152 2321 3158
rect 2302 3112 2305 3118
rect 2318 3072 2321 3138
rect 2326 3082 2329 3158
rect 2350 3142 2353 3178
rect 2358 3152 2361 3298
rect 2366 3272 2369 3308
rect 2374 3262 2377 3278
rect 2382 3272 2385 3368
rect 2418 3348 2422 3351
rect 2430 3342 2433 3348
rect 2438 3342 2441 3418
rect 2462 3352 2465 3448
rect 2478 3402 2481 3458
rect 2494 3452 2497 3458
rect 2518 3442 2521 3518
rect 2526 3462 2529 3508
rect 2574 3492 2577 3548
rect 2598 3542 2601 3558
rect 2674 3548 2678 3551
rect 2630 3532 2633 3538
rect 2590 3482 2593 3528
rect 2598 3492 2601 3518
rect 2614 3482 2617 3518
rect 2486 3342 2489 3358
rect 2510 3342 2513 3408
rect 2526 3352 2529 3388
rect 2534 3382 2537 3468
rect 2542 3452 2545 3478
rect 2578 3458 2582 3461
rect 2562 3438 2566 3441
rect 2574 3401 2577 3418
rect 2566 3398 2577 3401
rect 2566 3352 2569 3398
rect 2582 3391 2585 3448
rect 2574 3388 2585 3391
rect 2574 3372 2577 3388
rect 2590 3382 2593 3478
rect 2622 3462 2625 3498
rect 2630 3472 2633 3508
rect 2638 3472 2641 3538
rect 2654 3532 2657 3538
rect 2678 3532 2681 3538
rect 2694 3532 2697 3548
rect 2638 3462 2641 3468
rect 2646 3462 2649 3488
rect 2610 3458 2614 3461
rect 2654 3451 2657 3528
rect 2662 3492 2665 3518
rect 2702 3492 2705 3558
rect 2718 3542 2721 3548
rect 2726 3512 2729 3548
rect 2734 3522 2737 3558
rect 2774 3552 2777 3598
rect 2798 3562 2801 3598
rect 2742 3512 2745 3548
rect 2782 3542 2785 3558
rect 2854 3552 2857 3558
rect 2822 3542 2825 3548
rect 2830 3542 2833 3548
rect 2862 3542 2865 3608
rect 2950 3562 2953 3568
rect 2966 3552 2969 3558
rect 2850 3538 2854 3541
rect 2914 3538 2918 3541
rect 2750 3522 2753 3538
rect 2766 3532 2769 3538
rect 2958 3532 2961 3548
rect 2974 3532 2977 3538
rect 2990 3532 2993 3548
rect 3014 3542 3017 3548
rect 2726 3482 2729 3508
rect 2766 3502 2769 3518
rect 2814 3512 2817 3518
rect 2722 3478 2726 3481
rect 2782 3472 2785 3508
rect 2822 3492 2825 3528
rect 2890 3518 2894 3521
rect 2838 3472 2841 3508
rect 2904 3503 2906 3507
rect 2910 3503 2913 3507
rect 2917 3503 2920 3507
rect 2878 3482 2881 3498
rect 2950 3492 2953 3518
rect 2974 3512 2977 3528
rect 2906 3488 2910 3491
rect 2966 3482 2969 3488
rect 2898 3478 2902 3481
rect 2870 3472 2873 3478
rect 2730 3468 2734 3471
rect 2694 3462 2697 3468
rect 2654 3448 2662 3451
rect 2622 3392 2625 3398
rect 2630 3392 2633 3408
rect 2654 3381 2657 3448
rect 2686 3432 2689 3458
rect 2726 3422 2729 3428
rect 2654 3378 2662 3381
rect 2582 3372 2585 3378
rect 2574 3352 2577 3368
rect 2518 3342 2521 3348
rect 2498 3338 2502 3341
rect 2390 3322 2393 3338
rect 2526 3332 2529 3348
rect 2566 3342 2569 3348
rect 2574 3342 2577 3348
rect 2546 3338 2550 3341
rect 2490 3328 2494 3331
rect 2558 3331 2561 3338
rect 2550 3328 2561 3331
rect 2590 3332 2593 3358
rect 2598 3352 2601 3358
rect 2606 3332 2609 3348
rect 2390 3242 2393 3318
rect 2414 3282 2417 3298
rect 2430 3272 2433 3288
rect 2446 3262 2449 3278
rect 2406 3252 2409 3258
rect 2430 3242 2433 3248
rect 2454 3232 2457 3318
rect 2502 3292 2505 3328
rect 2550 3292 2553 3328
rect 2462 3282 2465 3288
rect 2478 3262 2481 3278
rect 2510 3262 2513 3268
rect 2534 3262 2537 3278
rect 2614 3272 2617 3368
rect 2638 3362 2641 3368
rect 2678 3362 2681 3388
rect 2698 3358 2702 3361
rect 2622 3292 2625 3358
rect 2654 3352 2657 3358
rect 2646 3342 2649 3348
rect 2702 3342 2705 3348
rect 2650 3338 2662 3341
rect 2682 3338 2686 3341
rect 2718 3332 2721 3368
rect 2726 3362 2729 3398
rect 2742 3352 2745 3368
rect 2750 3342 2753 3448
rect 2790 3442 2793 3468
rect 2878 3462 2881 3478
rect 2958 3472 2961 3478
rect 2990 3472 2993 3488
rect 2978 3468 2982 3471
rect 2966 3462 2969 3468
rect 2998 3462 3001 3538
rect 3006 3462 3009 3528
rect 3022 3492 3025 3588
rect 3042 3558 3046 3561
rect 3066 3558 3070 3561
rect 3078 3552 3081 3628
rect 3094 3592 3097 3658
rect 3118 3652 3121 3658
rect 3118 3552 3121 3558
rect 3050 3538 3054 3541
rect 3074 3538 3078 3541
rect 3030 3481 3033 3538
rect 3022 3478 3033 3481
rect 2914 3458 2918 3461
rect 2986 3458 2990 3461
rect 2766 3382 2769 3418
rect 2814 3362 2817 3368
rect 2758 3352 2761 3358
rect 2830 3352 2833 3438
rect 2846 3432 2849 3448
rect 2862 3372 2865 3418
rect 2834 3348 2838 3351
rect 2730 3338 2734 3341
rect 2754 3338 2761 3341
rect 2682 3328 2686 3331
rect 2646 3292 2649 3328
rect 2726 3282 2729 3288
rect 2622 3272 2625 3278
rect 2630 3272 2633 3278
rect 2586 3268 2590 3271
rect 2618 3268 2622 3271
rect 2498 3248 2502 3251
rect 2522 3248 2526 3251
rect 2392 3203 2394 3207
rect 2398 3203 2401 3207
rect 2405 3203 2408 3207
rect 2442 3188 2446 3191
rect 2358 3132 2361 3138
rect 2374 3132 2377 3178
rect 2394 3158 2398 3161
rect 2382 3142 2385 3148
rect 2390 3142 2393 3148
rect 2398 3112 2401 3138
rect 2478 3132 2481 3218
rect 2446 3092 2449 3108
rect 2486 3092 2489 3168
rect 2550 3162 2553 3238
rect 2498 3148 2502 3151
rect 2530 3148 2534 3151
rect 2550 3142 2553 3158
rect 2558 3142 2561 3268
rect 2566 3262 2569 3268
rect 2614 3232 2617 3258
rect 2646 3252 2649 3258
rect 2646 3162 2649 3248
rect 2654 3182 2657 3258
rect 2670 3212 2673 3268
rect 2678 3262 2681 3268
rect 2686 3262 2689 3278
rect 2714 3268 2718 3271
rect 2678 3232 2681 3258
rect 2710 3252 2713 3258
rect 2746 3248 2750 3251
rect 2622 3142 2625 3148
rect 2498 3138 2502 3141
rect 2326 3072 2329 3078
rect 2334 3062 2337 3088
rect 2346 3068 2350 3071
rect 2358 3062 2361 3088
rect 2370 3078 2374 3081
rect 2382 3062 2385 3078
rect 2510 3072 2513 3118
rect 2518 3072 2521 3078
rect 2574 3072 2577 3088
rect 2590 3082 2593 3098
rect 2598 3072 2601 3108
rect 2606 3102 2609 3138
rect 2638 3132 2641 3158
rect 2654 3092 2657 3148
rect 2662 3122 2665 3168
rect 2686 3162 2689 3218
rect 2702 3212 2705 3248
rect 2710 3192 2713 3248
rect 2670 3152 2673 3158
rect 2742 3151 2745 3158
rect 2758 3152 2761 3338
rect 2834 3338 2838 3341
rect 2774 3332 2777 3338
rect 2782 3332 2785 3338
rect 2766 3262 2769 3318
rect 2774 3292 2777 3318
rect 2790 3272 2793 3278
rect 2830 3271 2833 3328
rect 2826 3268 2833 3271
rect 2846 3272 2849 3368
rect 2894 3362 2897 3458
rect 2930 3448 2934 3451
rect 2950 3371 2953 3418
rect 2958 3402 2961 3458
rect 3014 3452 3017 3458
rect 3022 3452 3025 3478
rect 3038 3471 3041 3518
rect 3110 3502 3113 3548
rect 3082 3488 3086 3491
rect 3030 3468 3041 3471
rect 3074 3468 3078 3471
rect 2950 3368 2958 3371
rect 2954 3358 2958 3361
rect 2862 3352 2865 3358
rect 2858 3268 2862 3271
rect 2814 3262 2817 3268
rect 2790 3252 2793 3258
rect 2826 3248 2830 3251
rect 2766 3192 2769 3228
rect 2798 3172 2801 3248
rect 2814 3202 2817 3218
rect 2838 3192 2841 3258
rect 2846 3242 2849 3268
rect 2870 3262 2873 3288
rect 2886 3231 2889 3358
rect 2898 3338 2902 3341
rect 2966 3322 2969 3348
rect 2974 3342 2977 3358
rect 2990 3352 2993 3358
rect 2986 3338 2990 3341
rect 3006 3332 3009 3338
rect 3014 3322 3017 3328
rect 2904 3303 2906 3307
rect 2910 3303 2913 3307
rect 2917 3303 2920 3307
rect 2926 3282 2929 3298
rect 2934 3272 2937 3318
rect 2974 3292 2977 3318
rect 3022 3292 3025 3448
rect 3030 3441 3033 3468
rect 3042 3458 3046 3461
rect 3054 3442 3057 3448
rect 3030 3438 3038 3441
rect 3046 3432 3049 3438
rect 3062 3432 3065 3458
rect 3102 3432 3105 3478
rect 3110 3452 3113 3488
rect 3118 3462 3121 3538
rect 3126 3492 3129 3548
rect 3150 3542 3153 3658
rect 3158 3552 3161 3618
rect 3134 3532 3137 3538
rect 3142 3532 3145 3538
rect 3150 3521 3153 3528
rect 3142 3518 3153 3521
rect 3142 3462 3145 3518
rect 3174 3512 3177 3658
rect 3222 3642 3225 3668
rect 3222 3572 3225 3638
rect 3274 3618 3278 3621
rect 3202 3568 3206 3571
rect 3190 3552 3193 3568
rect 3198 3552 3201 3558
rect 3302 3552 3305 3618
rect 3318 3592 3321 3668
rect 3370 3658 3374 3661
rect 3326 3652 3329 3658
rect 3326 3552 3329 3648
rect 3434 3618 3438 3621
rect 3350 3552 3353 3558
rect 3398 3552 3401 3608
rect 3416 3603 3418 3607
rect 3422 3603 3425 3607
rect 3429 3603 3432 3607
rect 3158 3482 3161 3488
rect 3142 3452 3145 3458
rect 3114 3448 3118 3451
rect 3126 3442 3129 3448
rect 3150 3442 3153 3478
rect 3182 3472 3185 3528
rect 3190 3492 3193 3498
rect 3254 3482 3257 3538
rect 3270 3482 3273 3547
rect 3030 3392 3033 3428
rect 3062 3382 3065 3428
rect 3134 3422 3137 3428
rect 3030 3292 3033 3368
rect 3046 3352 3049 3378
rect 3038 3302 3041 3338
rect 2998 3282 3001 3288
rect 3026 3278 3030 3281
rect 2950 3272 2953 3278
rect 2894 3262 2897 3268
rect 2886 3228 2897 3231
rect 2894 3222 2897 3228
rect 2818 3188 2822 3191
rect 2854 3172 2857 3218
rect 2886 3172 2889 3218
rect 2742 3148 2750 3151
rect 2678 3142 2681 3148
rect 2702 3142 2705 3148
rect 2738 3138 2742 3141
rect 2766 3141 2769 3158
rect 2778 3148 2782 3151
rect 2766 3138 2774 3141
rect 2806 3132 2809 3168
rect 2838 3162 2841 3168
rect 2894 3142 2897 3218
rect 2818 3138 2822 3141
rect 2722 3128 2726 3131
rect 2902 3131 2905 3228
rect 2918 3142 2921 3258
rect 2958 3252 2961 3268
rect 2966 3262 2969 3268
rect 3022 3262 3025 3268
rect 3030 3262 3033 3278
rect 3054 3272 3057 3338
rect 3062 3332 3065 3358
rect 3082 3348 3086 3351
rect 3094 3342 3097 3358
rect 3134 3351 3137 3358
rect 3134 3348 3142 3351
rect 3130 3338 3134 3341
rect 3114 3328 3118 3331
rect 3070 3312 3073 3328
rect 3094 3302 3097 3318
rect 3062 3282 3065 3288
rect 3102 3272 3105 3288
rect 3090 3268 3094 3271
rect 2970 3258 2977 3261
rect 2930 3248 2934 3251
rect 2942 3162 2945 3218
rect 2974 3192 2977 3258
rect 2966 3142 2969 3168
rect 2998 3152 3001 3258
rect 3054 3252 3057 3268
rect 3110 3262 3113 3278
rect 3126 3262 3129 3328
rect 3142 3262 3145 3268
rect 3066 3248 3070 3251
rect 3078 3242 3081 3258
rect 3126 3252 3129 3258
rect 3090 3238 3094 3241
rect 2894 3128 2905 3131
rect 2982 3132 2985 3148
rect 2694 3112 2697 3128
rect 2706 3118 2710 3121
rect 2718 3092 2721 3108
rect 2742 3092 2745 3128
rect 2798 3092 2801 3118
rect 2678 3072 2681 3078
rect 2450 3068 2454 3071
rect 2722 3068 2726 3071
rect 2570 3058 2574 3061
rect 2602 3058 2606 3061
rect 2158 3052 2161 3058
rect 2198 3052 2201 3058
rect 2350 3052 2353 3058
rect 2622 3052 2625 3068
rect 2694 3062 2697 3068
rect 2654 3052 2657 3058
rect 2226 3048 2230 3051
rect 2426 3048 2430 3051
rect 2650 3048 2654 3051
rect 2702 3051 2705 3058
rect 2698 3048 2705 3051
rect 2254 3042 2257 3048
rect 2366 3042 2369 3048
rect 2582 3042 2585 3048
rect 2062 2962 2065 2988
rect 2062 2942 2065 2958
rect 2070 2952 2073 2998
rect 2078 2992 2081 3018
rect 2150 3002 2153 3018
rect 2118 2982 2121 2988
rect 2086 2972 2089 2978
rect 2106 2958 2110 2961
rect 2130 2958 2134 2961
rect 2150 2952 2153 2968
rect 2166 2962 2169 2978
rect 2214 2962 2217 3018
rect 2230 2962 2233 2978
rect 2158 2952 2161 2958
rect 2082 2948 2086 2951
rect 2070 2902 2073 2938
rect 2110 2932 2113 2948
rect 2158 2942 2161 2948
rect 2182 2942 2185 2948
rect 2134 2932 2137 2938
rect 2198 2932 2201 2958
rect 2218 2948 2222 2951
rect 2230 2931 2233 2958
rect 2238 2952 2241 3018
rect 2254 2962 2257 3038
rect 2286 2982 2289 3018
rect 2392 3003 2394 3007
rect 2398 3003 2401 3007
rect 2405 3003 2408 3007
rect 2414 2992 2417 3018
rect 2266 2968 2270 2971
rect 2286 2962 2289 2968
rect 2298 2958 2302 2961
rect 2310 2942 2313 2968
rect 2242 2938 2246 2941
rect 2282 2938 2286 2941
rect 2318 2932 2321 2948
rect 2390 2942 2393 2988
rect 2638 2982 2641 3018
rect 2710 2992 2713 3068
rect 2750 3062 2753 3088
rect 2830 3082 2833 3118
rect 2862 3072 2865 3118
rect 2894 3092 2897 3128
rect 2904 3103 2906 3107
rect 2910 3103 2913 3107
rect 2917 3103 2920 3107
rect 2950 3102 2953 3118
rect 2990 3102 2993 3138
rect 2950 3072 2953 3078
rect 2974 3072 2977 3078
rect 2962 3068 2966 3071
rect 2746 3048 2753 3051
rect 2750 2992 2753 3048
rect 2774 3032 2777 3068
rect 2846 3062 2849 3068
rect 2806 3042 2809 3058
rect 2854 3012 2857 3068
rect 2902 3062 2905 3068
rect 2862 3052 2865 3058
rect 2562 2968 2566 2971
rect 2586 2958 2590 2961
rect 2230 2928 2238 2931
rect 2158 2922 2161 2928
rect 1918 2872 1921 2888
rect 1966 2878 1993 2881
rect 1966 2872 1969 2878
rect 1990 2872 1993 2878
rect 1762 2858 1766 2861
rect 1794 2858 1798 2861
rect 1650 2778 1654 2781
rect 1546 2748 1550 2751
rect 1566 2742 1569 2748
rect 1550 2672 1553 2738
rect 1582 2711 1585 2747
rect 1574 2708 1585 2711
rect 1510 2542 1513 2638
rect 1558 2592 1561 2659
rect 1518 2551 1521 2558
rect 1368 2403 1370 2407
rect 1374 2403 1377 2407
rect 1381 2403 1384 2407
rect 1394 2368 1398 2371
rect 1390 2302 1393 2318
rect 1390 2292 1393 2298
rect 1438 2278 1441 2488
rect 1446 2472 1449 2478
rect 1518 2472 1521 2478
rect 1526 2472 1529 2498
rect 1542 2492 1545 2518
rect 1462 2351 1465 2358
rect 1478 2342 1481 2358
rect 1502 2352 1505 2418
rect 1518 2392 1521 2438
rect 1494 2302 1497 2348
rect 1502 2302 1505 2338
rect 1518 2322 1521 2328
rect 1526 2312 1529 2468
rect 1550 2442 1553 2528
rect 1574 2521 1577 2708
rect 1590 2692 1593 2698
rect 1630 2682 1633 2768
rect 1702 2762 1705 2768
rect 1758 2762 1761 2768
rect 1670 2732 1673 2758
rect 1730 2748 1734 2751
rect 1766 2742 1769 2838
rect 1774 2792 1777 2848
rect 1782 2802 1785 2848
rect 1814 2842 1817 2848
rect 1830 2842 1833 2868
rect 1846 2852 1849 2858
rect 1854 2842 1857 2868
rect 1974 2862 1977 2868
rect 1982 2862 1985 2868
rect 1938 2858 1942 2861
rect 1898 2848 1902 2851
rect 1790 2792 1793 2818
rect 1774 2752 1777 2788
rect 1814 2762 1817 2838
rect 1822 2782 1825 2818
rect 1862 2792 1865 2848
rect 2006 2842 2009 2848
rect 1834 2788 1838 2791
rect 1826 2768 1830 2771
rect 1838 2762 1841 2778
rect 1782 2742 1785 2758
rect 1814 2742 1817 2748
rect 1706 2738 1710 2741
rect 1830 2741 1833 2758
rect 1838 2752 1841 2758
rect 1830 2738 1838 2741
rect 1726 2732 1729 2738
rect 1662 2721 1665 2728
rect 1742 2722 1745 2738
rect 1878 2732 1881 2798
rect 1902 2762 1905 2788
rect 1918 2752 1921 2778
rect 1914 2748 1918 2751
rect 1926 2742 1929 2828
rect 1934 2762 1937 2798
rect 1998 2792 2001 2838
rect 2022 2822 2025 2868
rect 2030 2852 2033 2888
rect 2066 2878 2070 2881
rect 2082 2868 2086 2871
rect 2094 2862 2097 2868
rect 2102 2862 2105 2888
rect 2126 2882 2129 2898
rect 2142 2892 2145 2898
rect 2258 2888 2262 2891
rect 2138 2878 2142 2881
rect 2110 2862 2113 2868
rect 2126 2862 2129 2868
rect 2042 2858 2046 2861
rect 2050 2838 2054 2841
rect 2066 2838 2070 2841
rect 2038 2832 2041 2838
rect 2094 2832 2097 2858
rect 2150 2842 2153 2868
rect 2158 2862 2161 2868
rect 2166 2852 2169 2878
rect 2174 2872 2177 2878
rect 2174 2862 2177 2868
rect 2198 2862 2201 2868
rect 2246 2862 2249 2868
rect 2286 2862 2289 2868
rect 2294 2862 2297 2908
rect 2302 2902 2305 2918
rect 2342 2882 2345 2908
rect 2302 2872 2305 2878
rect 2334 2872 2337 2878
rect 2334 2862 2337 2868
rect 2358 2862 2361 2918
rect 2422 2892 2425 2938
rect 2462 2892 2465 2958
rect 2510 2952 2513 2958
rect 2526 2952 2529 2958
rect 2614 2952 2617 2958
rect 2622 2952 2625 2958
rect 2374 2872 2377 2878
rect 2314 2848 2318 2851
rect 2186 2838 2190 2841
rect 2178 2818 2182 2821
rect 2054 2792 2057 2798
rect 2122 2788 2126 2791
rect 2222 2782 2225 2818
rect 1954 2768 1958 2771
rect 1938 2748 1942 2751
rect 1950 2742 1953 2758
rect 1930 2738 1934 2741
rect 1910 2732 1913 2738
rect 1662 2718 1673 2721
rect 1714 2718 1718 2721
rect 1566 2518 1577 2521
rect 1566 2492 1569 2518
rect 1598 2492 1601 2668
rect 1630 2662 1633 2678
rect 1606 2542 1609 2638
rect 1614 2542 1617 2548
rect 1646 2522 1649 2658
rect 1654 2592 1657 2658
rect 1670 2652 1673 2718
rect 1758 2692 1761 2728
rect 1798 2722 1801 2728
rect 1958 2722 1961 2728
rect 1966 2712 1969 2738
rect 1974 2732 1977 2778
rect 1994 2768 1998 2771
rect 2006 2762 2009 2768
rect 1998 2752 2001 2758
rect 2022 2752 2025 2768
rect 2070 2742 2073 2748
rect 2038 2712 2041 2728
rect 1698 2679 1705 2681
rect 1694 2678 1705 2679
rect 1702 2662 1705 2678
rect 1718 2672 1721 2678
rect 1702 2642 1705 2648
rect 1662 2562 1665 2568
rect 1682 2538 1686 2541
rect 1694 2532 1697 2628
rect 1702 2592 1705 2638
rect 1734 2621 1737 2659
rect 1726 2618 1737 2621
rect 1726 2592 1729 2618
rect 1734 2592 1737 2598
rect 1750 2592 1753 2598
rect 1682 2528 1686 2531
rect 1694 2521 1697 2528
rect 1686 2518 1697 2521
rect 1606 2472 1609 2478
rect 1674 2468 1678 2471
rect 1558 2392 1561 2438
rect 1566 2432 1569 2458
rect 1574 2442 1577 2448
rect 1598 2432 1601 2448
rect 1678 2442 1681 2458
rect 1566 2382 1569 2428
rect 1614 2392 1617 2428
rect 1662 2362 1665 2418
rect 1670 2352 1673 2358
rect 1582 2342 1585 2348
rect 1686 2342 1689 2518
rect 1710 2412 1713 2548
rect 1746 2528 1750 2531
rect 1718 2512 1721 2528
rect 1722 2468 1726 2471
rect 1738 2459 1742 2462
rect 1758 2402 1761 2458
rect 1774 2432 1777 2478
rect 1758 2392 1761 2398
rect 1710 2382 1713 2388
rect 1698 2368 1702 2371
rect 1726 2362 1729 2378
rect 1742 2362 1745 2368
rect 1750 2362 1753 2378
rect 1766 2362 1769 2368
rect 1718 2352 1721 2358
rect 1634 2338 1638 2341
rect 1574 2331 1577 2338
rect 1574 2328 1585 2331
rect 1478 2292 1481 2298
rect 1518 2292 1521 2298
rect 1286 2272 1289 2278
rect 1558 2272 1561 2318
rect 1354 2268 1358 2271
rect 1538 2268 1542 2271
rect 1570 2268 1574 2271
rect 1198 2252 1201 2259
rect 1282 2258 1286 2261
rect 1186 2188 1190 2191
rect 1334 2162 1337 2268
rect 1342 2262 1345 2268
rect 1290 2158 1294 2161
rect 1062 2151 1065 2158
rect 1158 2151 1161 2158
rect 1358 2152 1361 2268
rect 1394 2258 1398 2261
rect 1382 2252 1385 2258
rect 1402 2238 1406 2241
rect 1368 2203 1370 2207
rect 1374 2203 1377 2207
rect 1381 2203 1384 2207
rect 1414 2202 1417 2268
rect 1430 2242 1433 2258
rect 1438 2192 1441 2218
rect 1462 2202 1465 2268
rect 1510 2262 1513 2268
rect 1558 2262 1561 2268
rect 1546 2258 1550 2261
rect 1562 2248 1566 2251
rect 1470 2242 1473 2248
rect 1470 2182 1473 2238
rect 1526 2222 1529 2248
rect 1542 2212 1545 2218
rect 1566 2182 1569 2188
rect 1542 2172 1545 2178
rect 1550 2158 1558 2161
rect 1542 2152 1545 2158
rect 1222 2142 1225 2148
rect 1250 2147 1254 2150
rect 1394 2148 1398 2151
rect 1490 2148 1494 2151
rect 1078 2132 1081 2138
rect 1094 2122 1097 2128
rect 982 2082 985 2098
rect 1086 2092 1089 2098
rect 1038 2088 1046 2091
rect 1018 2078 1022 2081
rect 1030 2072 1033 2078
rect 1038 2072 1041 2088
rect 1150 2082 1153 2138
rect 1318 2131 1321 2148
rect 1422 2142 1425 2148
rect 1502 2142 1505 2148
rect 1054 2072 1057 2078
rect 1070 2072 1073 2078
rect 1010 2068 1014 2071
rect 950 2062 953 2068
rect 962 2058 966 2061
rect 1026 2058 1030 2061
rect 1078 2052 1081 2078
rect 1214 2072 1217 2108
rect 1274 2088 1278 2091
rect 1262 2072 1265 2078
rect 1066 2048 1070 2051
rect 1118 2042 1121 2058
rect 994 1968 998 1971
rect 870 1962 873 1968
rect 822 1952 825 1958
rect 834 1948 838 1951
rect 834 1938 838 1941
rect 854 1932 857 1958
rect 886 1942 889 1948
rect 902 1942 905 1968
rect 930 1958 934 1961
rect 986 1958 990 1961
rect 910 1952 913 1958
rect 914 1948 918 1951
rect 926 1942 929 1948
rect 942 1942 945 1958
rect 806 1842 809 1918
rect 856 1903 858 1907
rect 862 1903 865 1907
rect 869 1903 872 1907
rect 918 1892 921 1938
rect 874 1888 878 1891
rect 814 1822 817 1858
rect 798 1812 801 1818
rect 822 1752 825 1888
rect 838 1882 841 1888
rect 886 1881 889 1888
rect 882 1878 889 1881
rect 918 1862 921 1868
rect 886 1852 889 1858
rect 846 1802 849 1818
rect 910 1781 913 1848
rect 926 1842 929 1938
rect 958 1922 961 1928
rect 966 1892 969 1938
rect 974 1932 977 1948
rect 990 1942 993 1948
rect 1006 1942 1009 2038
rect 1150 2032 1153 2059
rect 1246 2052 1249 2059
rect 1182 2042 1185 2048
rect 1278 1992 1281 2048
rect 1294 1992 1297 2128
rect 1314 2128 1321 2131
rect 1338 2118 1342 2121
rect 1310 2072 1313 2078
rect 1358 2072 1361 2138
rect 1470 2092 1473 2108
rect 1486 2092 1489 2118
rect 1418 2088 1422 2091
rect 1334 2062 1337 2068
rect 1146 1988 1150 1991
rect 1058 1968 1062 1971
rect 1114 1968 1118 1971
rect 1154 1968 1158 1971
rect 1018 1948 1022 1951
rect 1034 1948 1038 1951
rect 1046 1942 1049 1958
rect 1062 1952 1065 1958
rect 1042 1938 1046 1941
rect 1078 1932 1081 1968
rect 1110 1952 1113 1958
rect 1130 1948 1134 1951
rect 1086 1942 1089 1948
rect 1102 1942 1105 1948
rect 990 1882 993 1898
rect 998 1882 1001 1918
rect 1014 1892 1017 1928
rect 1086 1912 1089 1928
rect 1134 1902 1137 1938
rect 1154 1928 1158 1931
rect 1166 1892 1169 1948
rect 1206 1892 1209 1978
rect 1222 1951 1225 1958
rect 1254 1952 1257 1958
rect 1034 1888 1041 1891
rect 1038 1872 1041 1888
rect 1094 1888 1102 1891
rect 1194 1888 1201 1891
rect 1054 1872 1057 1878
rect 1094 1872 1097 1888
rect 1198 1872 1201 1888
rect 1238 1872 1241 1938
rect 1262 1932 1265 1968
rect 1290 1958 1294 1961
rect 1302 1952 1305 2018
rect 1318 1952 1321 1958
rect 1282 1948 1286 1951
rect 1294 1948 1302 1951
rect 1294 1942 1297 1948
rect 1310 1942 1313 1948
rect 1274 1938 1278 1941
rect 1314 1938 1318 1941
rect 1330 1938 1334 1941
rect 1270 1892 1273 1938
rect 1342 1932 1345 2068
rect 1390 2022 1393 2068
rect 1438 2062 1441 2068
rect 1368 2003 1370 2007
rect 1374 2003 1377 2007
rect 1381 2003 1384 2007
rect 1446 1992 1449 2068
rect 1478 2062 1481 2088
rect 1494 2082 1497 2098
rect 1502 2092 1505 2128
rect 1534 2092 1537 2138
rect 1458 2058 1462 2061
rect 1478 1992 1481 2038
rect 1354 1988 1358 1991
rect 1418 1978 1422 1981
rect 1494 1952 1497 2078
rect 1518 2062 1521 2078
rect 1550 2062 1553 2158
rect 1558 2152 1561 2158
rect 1574 2132 1577 2138
rect 1582 2132 1585 2328
rect 1598 2292 1601 2335
rect 1622 2292 1625 2298
rect 1606 2282 1609 2288
rect 1594 2278 1598 2281
rect 1630 2272 1633 2308
rect 1594 2268 1598 2271
rect 1590 2252 1593 2258
rect 1618 2248 1625 2251
rect 1614 2152 1617 2168
rect 1590 2142 1593 2148
rect 1582 2121 1585 2128
rect 1574 2118 1585 2121
rect 1562 2078 1566 2081
rect 1562 2068 1566 2071
rect 1554 2058 1558 2061
rect 1502 1992 1505 2048
rect 1502 1972 1505 1988
rect 1558 1962 1561 2018
rect 1566 1992 1569 2058
rect 1574 2052 1577 2118
rect 1586 2088 1590 2091
rect 1582 2072 1585 2078
rect 1582 2062 1585 2068
rect 1590 2051 1593 2078
rect 1582 2048 1593 2051
rect 1582 1992 1585 2048
rect 1622 1992 1625 2248
rect 1574 1972 1577 1978
rect 1630 1962 1633 2268
rect 1638 2242 1641 2248
rect 1654 2182 1657 2332
rect 1710 2312 1713 2348
rect 1726 2342 1729 2358
rect 1738 2328 1742 2331
rect 1734 2292 1737 2298
rect 1718 2272 1721 2278
rect 1702 2252 1705 2259
rect 1766 2252 1769 2348
rect 1774 2342 1777 2428
rect 1782 2392 1785 2708
rect 1872 2703 1874 2707
rect 1878 2703 1881 2707
rect 1885 2703 1888 2707
rect 1798 2692 1801 2698
rect 1894 2692 1897 2698
rect 1934 2692 1937 2708
rect 1966 2682 1969 2698
rect 2046 2692 2049 2738
rect 2118 2732 2121 2738
rect 2058 2728 2062 2731
rect 2078 2692 2081 2708
rect 2102 2702 2105 2718
rect 2046 2682 2049 2688
rect 1814 2672 1817 2678
rect 1830 2663 1833 2668
rect 1918 2662 1921 2678
rect 1926 2672 1929 2678
rect 1966 2672 1969 2678
rect 1986 2668 1990 2671
rect 1954 2658 1958 2661
rect 1986 2658 1990 2661
rect 1934 2652 1937 2658
rect 2006 2652 2009 2668
rect 2018 2666 2022 2669
rect 2062 2662 2065 2668
rect 2038 2652 2041 2658
rect 2070 2652 2073 2688
rect 2126 2672 2129 2718
rect 2142 2692 2145 2758
rect 2178 2748 2182 2751
rect 2230 2692 2233 2818
rect 2254 2792 2257 2838
rect 2306 2788 2310 2791
rect 2310 2762 2313 2788
rect 2334 2772 2337 2848
rect 2366 2842 2369 2848
rect 2342 2792 2345 2838
rect 2350 2772 2353 2818
rect 2366 2791 2369 2828
rect 2374 2802 2377 2868
rect 2382 2862 2385 2868
rect 2392 2803 2394 2807
rect 2398 2803 2401 2807
rect 2405 2803 2408 2807
rect 2366 2788 2374 2791
rect 2338 2768 2342 2771
rect 2378 2768 2382 2771
rect 2330 2758 2334 2761
rect 2246 2751 2249 2758
rect 2342 2752 2345 2758
rect 2350 2752 2353 2768
rect 2370 2758 2374 2761
rect 2402 2758 2406 2761
rect 2370 2748 2374 2751
rect 2094 2662 2097 2668
rect 2126 2662 2129 2668
rect 2090 2658 2094 2661
rect 2134 2652 2137 2678
rect 2170 2668 2174 2671
rect 2214 2670 2217 2678
rect 2178 2658 2182 2661
rect 2238 2652 2241 2658
rect 2002 2648 2006 2651
rect 2202 2648 2206 2651
rect 1990 2642 1993 2648
rect 2054 2632 2057 2638
rect 2246 2632 2249 2728
rect 2310 2682 2313 2698
rect 2342 2692 2345 2708
rect 2414 2692 2417 2748
rect 2422 2732 2425 2878
rect 2430 2852 2433 2878
rect 2458 2848 2462 2851
rect 2430 2772 2433 2848
rect 2478 2782 2481 2947
rect 2630 2942 2633 2948
rect 2522 2938 2526 2941
rect 2586 2938 2590 2941
rect 2610 2938 2614 2941
rect 2494 2882 2497 2938
rect 2594 2928 2598 2931
rect 2562 2888 2566 2891
rect 2614 2872 2617 2908
rect 2638 2882 2641 2978
rect 2758 2972 2761 3008
rect 2838 2992 2841 3008
rect 2878 2992 2881 3048
rect 2934 3012 2937 3018
rect 2958 2992 2961 3068
rect 2982 3062 2985 3098
rect 3006 3082 3009 3178
rect 3038 3162 3041 3238
rect 3150 3212 3153 3438
rect 3158 3432 3161 3448
rect 3166 3351 3169 3468
rect 3174 3362 3177 3458
rect 3182 3412 3185 3468
rect 3254 3452 3257 3459
rect 3202 3388 3206 3391
rect 3202 3368 3206 3371
rect 3190 3352 3193 3358
rect 3166 3348 3177 3351
rect 3166 3332 3169 3338
rect 3158 3292 3161 3318
rect 3174 3292 3177 3348
rect 3190 3332 3193 3338
rect 3166 3252 3169 3278
rect 3182 3242 3185 3268
rect 3198 3262 3201 3358
rect 3214 3352 3217 3378
rect 3226 3358 3230 3361
rect 3246 3352 3249 3358
rect 3270 3342 3273 3378
rect 3286 3362 3289 3428
rect 3318 3352 3321 3408
rect 3306 3338 3310 3341
rect 3262 3332 3265 3338
rect 3226 3328 3230 3331
rect 3254 3328 3262 3331
rect 3162 3218 3166 3221
rect 3034 3158 3038 3161
rect 3014 3152 3017 3158
rect 3094 3142 3097 3148
rect 3102 3142 3105 3208
rect 3174 3192 3177 3208
rect 3190 3192 3193 3258
rect 3198 3252 3201 3258
rect 3206 3242 3209 3278
rect 3246 3262 3249 3328
rect 3254 3282 3257 3328
rect 3294 3292 3297 3318
rect 3254 3262 3257 3278
rect 3286 3272 3289 3278
rect 3302 3272 3305 3328
rect 3326 3292 3329 3458
rect 3334 3392 3337 3548
rect 3342 3462 3345 3498
rect 3358 3492 3361 3548
rect 3398 3492 3401 3548
rect 3418 3538 3422 3541
rect 3370 3488 3374 3491
rect 3342 3392 3345 3398
rect 3358 3352 3361 3478
rect 3446 3472 3449 3548
rect 3454 3542 3457 3548
rect 3462 3532 3465 3668
rect 3670 3662 3673 3668
rect 3494 3632 3497 3659
rect 3650 3658 3654 3661
rect 3558 3652 3561 3658
rect 3582 3642 3585 3658
rect 3638 3622 3641 3658
rect 3618 3618 3622 3621
rect 3598 3552 3601 3618
rect 3638 3552 3641 3558
rect 3494 3531 3497 3548
rect 3626 3548 3630 3551
rect 3642 3548 3646 3551
rect 3454 3462 3457 3518
rect 3462 3482 3465 3528
rect 3490 3528 3497 3531
rect 3502 3512 3505 3518
rect 3534 3502 3537 3538
rect 3566 3522 3569 3547
rect 3582 3532 3585 3538
rect 3618 3528 3622 3531
rect 3654 3521 3657 3628
rect 3674 3548 3681 3551
rect 3662 3532 3665 3538
rect 3670 3522 3673 3528
rect 3678 3522 3681 3548
rect 3654 3518 3662 3521
rect 3478 3472 3481 3498
rect 3606 3492 3609 3498
rect 3630 3492 3633 3518
rect 3694 3512 3697 3658
rect 3494 3479 3502 3481
rect 3494 3478 3505 3479
rect 3634 3478 3638 3481
rect 3494 3462 3497 3478
rect 3630 3462 3633 3468
rect 3638 3462 3641 3468
rect 3398 3392 3401 3458
rect 3542 3412 3545 3459
rect 3574 3452 3577 3458
rect 3416 3403 3418 3407
rect 3422 3403 3425 3407
rect 3429 3403 3432 3407
rect 3570 3388 3574 3391
rect 3590 3372 3593 3448
rect 3546 3368 3550 3371
rect 3630 3352 3633 3368
rect 3670 3352 3673 3508
rect 3702 3502 3705 3658
rect 3750 3561 3753 3648
rect 3758 3642 3761 3648
rect 3758 3552 3761 3618
rect 3686 3482 3689 3488
rect 3710 3472 3713 3538
rect 3718 3522 3721 3548
rect 3730 3538 3734 3541
rect 3762 3538 3766 3541
rect 3718 3482 3721 3518
rect 3686 3392 3689 3458
rect 3702 3452 3705 3458
rect 3726 3402 3729 3528
rect 3782 3492 3785 3728
rect 3928 3703 3930 3707
rect 3934 3703 3937 3707
rect 3941 3703 3944 3707
rect 3958 3702 3961 3728
rect 3982 3692 3985 3728
rect 3998 3728 4002 3732
rect 4078 3728 4082 3732
rect 4110 3731 4114 3732
rect 4110 3728 4121 3731
rect 3998 3702 4001 3728
rect 4078 3702 4081 3728
rect 3858 3688 3862 3691
rect 3806 3663 3809 3688
rect 4086 3682 4089 3688
rect 4102 3682 4105 3688
rect 3822 3652 3825 3668
rect 3846 3662 3849 3678
rect 3854 3672 3857 3678
rect 3954 3668 3958 3671
rect 4054 3663 4057 3678
rect 3862 3642 3865 3658
rect 3806 3552 3809 3568
rect 3890 3558 3894 3561
rect 3902 3552 3905 3658
rect 3910 3632 3913 3658
rect 3966 3642 3969 3658
rect 4006 3642 4009 3648
rect 4070 3642 4073 3668
rect 4086 3662 4089 3678
rect 4098 3668 4102 3671
rect 4110 3652 4113 3658
rect 3986 3638 3990 3641
rect 3814 3512 3817 3548
rect 3822 3542 3825 3548
rect 3846 3542 3849 3548
rect 3854 3531 3857 3548
rect 3854 3528 3862 3531
rect 3886 3522 3889 3548
rect 3870 3492 3873 3508
rect 3774 3442 3777 3468
rect 3714 3348 3718 3351
rect 3358 3302 3361 3348
rect 3434 3338 3438 3341
rect 3482 3338 3486 3341
rect 3382 3311 3385 3338
rect 3374 3308 3385 3311
rect 3310 3272 3313 3288
rect 3358 3272 3361 3278
rect 3298 3268 3302 3271
rect 3290 3258 3294 3261
rect 3214 3242 3217 3258
rect 3274 3248 3278 3251
rect 3198 3192 3201 3238
rect 3222 3212 3225 3248
rect 3246 3242 3249 3248
rect 3246 3192 3249 3238
rect 3254 3182 3257 3218
rect 3134 3152 3137 3158
rect 3158 3142 3161 3158
rect 3174 3152 3177 3158
rect 3230 3152 3233 3158
rect 3190 3142 3193 3148
rect 3238 3142 3241 3158
rect 3278 3152 3281 3188
rect 3038 3112 3041 3118
rect 3046 3092 3049 3138
rect 3150 3121 3153 3138
rect 3146 3118 3161 3121
rect 3182 3121 3185 3138
rect 3262 3132 3265 3138
rect 3178 3118 3185 3121
rect 3058 3078 3062 3081
rect 2970 3058 2974 3061
rect 2990 3051 2993 3078
rect 3006 3072 3009 3078
rect 3018 3068 3022 3071
rect 2986 3048 2993 3051
rect 2998 3052 3001 3058
rect 3034 3048 3038 3051
rect 2974 2992 2977 3038
rect 2982 3022 2985 3048
rect 3070 3032 3073 3118
rect 3126 3072 3129 3078
rect 3022 3022 3025 3028
rect 2686 2962 2689 2968
rect 2694 2962 2697 2968
rect 2706 2948 2710 2951
rect 2654 2932 2657 2938
rect 2670 2932 2673 2938
rect 2686 2932 2689 2948
rect 2718 2942 2721 2948
rect 2726 2932 2729 2968
rect 2738 2958 2742 2961
rect 2738 2948 2742 2951
rect 2746 2948 2750 2951
rect 2802 2948 2806 2951
rect 2866 2948 2870 2951
rect 2778 2938 2782 2941
rect 2794 2938 2798 2941
rect 2770 2928 2774 2931
rect 2802 2928 2806 2931
rect 2646 2922 2649 2928
rect 2846 2922 2849 2938
rect 2854 2932 2857 2948
rect 2878 2932 2881 2948
rect 2886 2942 2889 2968
rect 2886 2932 2889 2938
rect 2702 2892 2705 2918
rect 2562 2868 2566 2871
rect 2458 2747 2462 2750
rect 2282 2678 2286 2681
rect 2254 2670 2257 2678
rect 2274 2668 2278 2671
rect 2262 2662 2265 2668
rect 2286 2662 2289 2668
rect 2302 2652 2305 2678
rect 2310 2662 2313 2668
rect 2326 2662 2329 2668
rect 2334 2652 2337 2678
rect 2398 2672 2401 2688
rect 2422 2682 2425 2728
rect 2406 2672 2409 2678
rect 2438 2672 2441 2738
rect 2374 2662 2377 2668
rect 2378 2658 2382 2661
rect 2290 2648 2294 2651
rect 2354 2648 2358 2651
rect 2418 2648 2422 2651
rect 1998 2622 2001 2628
rect 1950 2592 1953 2598
rect 1954 2578 1958 2581
rect 1798 2492 1801 2578
rect 1814 2551 1817 2568
rect 1806 2472 1809 2538
rect 1822 2492 1825 2498
rect 1794 2458 1798 2461
rect 1790 2442 1793 2448
rect 1798 2442 1801 2448
rect 1806 2381 1809 2468
rect 1814 2392 1817 2468
rect 1806 2378 1817 2381
rect 1802 2368 1806 2371
rect 1790 2262 1793 2328
rect 1798 2322 1801 2328
rect 1806 2301 1809 2338
rect 1798 2298 1809 2301
rect 1798 2282 1801 2298
rect 1718 2192 1721 2238
rect 1766 2192 1769 2238
rect 1798 2221 1801 2259
rect 1798 2218 1809 2221
rect 1806 2182 1809 2218
rect 1650 2168 1654 2171
rect 1646 2152 1649 2158
rect 1654 2152 1657 2158
rect 1638 2132 1641 2138
rect 1654 2132 1657 2138
rect 1662 2122 1665 2168
rect 1702 2162 1705 2168
rect 1678 2142 1681 2148
rect 1682 2138 1689 2141
rect 1594 1958 1598 1961
rect 1554 1948 1558 1951
rect 1586 1948 1590 1951
rect 1594 1948 1598 1951
rect 1350 1942 1353 1948
rect 1446 1942 1449 1948
rect 1498 1938 1502 1941
rect 1390 1932 1393 1938
rect 1358 1928 1366 1931
rect 1326 1922 1329 1928
rect 1294 1902 1297 1918
rect 1318 1882 1321 1888
rect 986 1868 990 1871
rect 942 1862 945 1868
rect 958 1862 961 1868
rect 1018 1858 1022 1861
rect 1034 1858 1038 1861
rect 1054 1852 1057 1868
rect 1142 1862 1145 1868
rect 1082 1858 1086 1861
rect 946 1848 950 1851
rect 970 1848 974 1851
rect 1018 1848 1022 1851
rect 1042 1848 1046 1851
rect 998 1842 1001 1848
rect 918 1792 921 1818
rect 1006 1792 1009 1818
rect 1078 1782 1081 1818
rect 1150 1782 1153 1868
rect 1254 1792 1257 1868
rect 1310 1862 1313 1878
rect 1350 1862 1353 1868
rect 1270 1842 1273 1859
rect 1302 1852 1305 1858
rect 1318 1792 1321 1798
rect 910 1778 918 1781
rect 894 1772 897 1778
rect 902 1762 905 1768
rect 738 1748 742 1751
rect 798 1742 801 1748
rect 822 1742 825 1748
rect 830 1742 833 1748
rect 498 1738 502 1741
rect 778 1738 782 1741
rect 490 1728 494 1731
rect 374 1682 377 1698
rect 310 1678 318 1681
rect 302 1672 305 1678
rect 366 1672 369 1678
rect 310 1662 313 1668
rect 322 1666 326 1669
rect 346 1668 350 1671
rect 370 1658 374 1661
rect 394 1658 398 1661
rect 286 1652 289 1658
rect 254 1572 257 1648
rect 262 1632 265 1648
rect 398 1642 401 1648
rect 274 1638 278 1641
rect 298 1638 302 1641
rect 406 1631 409 1728
rect 422 1672 425 1708
rect 542 1692 545 1708
rect 558 1702 561 1738
rect 606 1721 609 1738
rect 614 1732 617 1738
rect 686 1732 689 1738
rect 698 1728 702 1731
rect 598 1718 609 1721
rect 598 1692 601 1718
rect 670 1692 673 1728
rect 694 1702 697 1718
rect 718 1692 721 1718
rect 430 1688 438 1691
rect 430 1672 433 1688
rect 694 1682 697 1688
rect 750 1682 753 1738
rect 766 1732 769 1738
rect 822 1702 825 1718
rect 856 1703 858 1707
rect 862 1703 865 1707
rect 869 1703 872 1707
rect 662 1678 686 1681
rect 706 1678 710 1681
rect 486 1672 489 1678
rect 622 1672 625 1678
rect 538 1668 542 1671
rect 662 1671 665 1678
rect 750 1672 753 1678
rect 758 1672 761 1698
rect 886 1692 889 1758
rect 898 1748 902 1751
rect 918 1732 921 1778
rect 926 1762 929 1768
rect 998 1762 1001 1778
rect 1146 1768 1150 1771
rect 966 1758 974 1761
rect 966 1752 969 1758
rect 950 1742 953 1748
rect 938 1738 942 1741
rect 958 1722 961 1738
rect 938 1688 942 1691
rect 814 1682 817 1688
rect 822 1682 825 1688
rect 886 1682 889 1688
rect 966 1682 969 1748
rect 974 1742 977 1748
rect 990 1732 993 1758
rect 1006 1752 1009 1758
rect 1014 1722 1017 1768
rect 1038 1762 1041 1768
rect 1086 1752 1089 1758
rect 1022 1748 1030 1751
rect 1022 1742 1025 1748
rect 1094 1742 1097 1758
rect 1182 1752 1185 1758
rect 1214 1751 1217 1758
rect 1102 1742 1105 1748
rect 1022 1692 1025 1738
rect 1030 1702 1033 1738
rect 1070 1732 1073 1738
rect 1142 1732 1145 1738
rect 1118 1712 1121 1728
rect 1130 1718 1134 1721
rect 990 1688 998 1691
rect 786 1678 790 1681
rect 842 1678 846 1681
rect 866 1678 870 1681
rect 930 1678 934 1681
rect 658 1668 665 1671
rect 698 1668 702 1671
rect 786 1668 793 1671
rect 478 1662 481 1668
rect 418 1658 422 1661
rect 398 1628 409 1631
rect 178 1558 182 1561
rect 182 1542 185 1548
rect 190 1542 193 1548
rect 206 1542 209 1558
rect 214 1552 217 1558
rect 230 1552 233 1568
rect 222 1542 225 1548
rect 254 1532 257 1568
rect 182 1462 185 1478
rect 134 1352 137 1358
rect 134 1272 137 1328
rect 58 1268 62 1271
rect 14 1212 17 1258
rect 30 1252 33 1258
rect 78 1252 81 1258
rect 58 1248 62 1251
rect 38 1202 41 1248
rect 110 1212 113 1258
rect 126 1252 129 1268
rect 142 1262 145 1328
rect 190 1292 193 1498
rect 198 1452 201 1488
rect 206 1482 209 1518
rect 222 1492 225 1518
rect 206 1462 209 1468
rect 218 1458 222 1461
rect 230 1452 233 1458
rect 246 1441 249 1518
rect 278 1492 281 1618
rect 326 1592 329 1608
rect 334 1571 337 1618
rect 344 1603 346 1607
rect 350 1603 353 1607
rect 357 1603 360 1607
rect 334 1568 345 1571
rect 314 1558 318 1561
rect 286 1542 289 1548
rect 294 1532 297 1558
rect 342 1552 345 1568
rect 382 1562 385 1568
rect 330 1548 334 1551
rect 302 1542 305 1548
rect 342 1542 345 1548
rect 358 1542 361 1558
rect 318 1492 321 1528
rect 282 1488 286 1491
rect 366 1482 369 1558
rect 378 1548 382 1551
rect 390 1542 393 1568
rect 398 1532 401 1628
rect 414 1572 417 1618
rect 446 1592 449 1658
rect 542 1632 545 1648
rect 506 1628 510 1631
rect 558 1562 561 1668
rect 566 1652 569 1668
rect 614 1662 617 1668
rect 634 1658 638 1661
rect 670 1652 673 1668
rect 718 1662 721 1668
rect 758 1662 761 1668
rect 682 1658 686 1661
rect 778 1658 782 1661
rect 630 1642 633 1648
rect 574 1592 577 1638
rect 630 1592 633 1628
rect 646 1612 649 1648
rect 742 1642 745 1658
rect 778 1648 782 1651
rect 426 1548 430 1551
rect 430 1542 433 1548
rect 590 1542 593 1558
rect 478 1532 481 1538
rect 486 1521 489 1538
rect 534 1532 537 1538
rect 486 1518 494 1521
rect 506 1518 510 1521
rect 542 1521 545 1538
rect 598 1532 601 1548
rect 638 1542 641 1578
rect 678 1572 681 1578
rect 654 1562 657 1568
rect 658 1548 662 1551
rect 650 1538 654 1541
rect 614 1532 617 1538
rect 670 1532 673 1558
rect 710 1552 713 1578
rect 790 1572 793 1668
rect 898 1668 902 1671
rect 798 1632 801 1668
rect 846 1662 849 1668
rect 806 1622 809 1658
rect 886 1652 889 1668
rect 918 1662 921 1668
rect 898 1658 902 1661
rect 850 1648 854 1651
rect 814 1602 817 1618
rect 830 1612 833 1648
rect 818 1578 822 1581
rect 818 1568 822 1571
rect 746 1548 750 1551
rect 718 1542 721 1548
rect 726 1542 729 1548
rect 734 1542 737 1548
rect 534 1518 545 1521
rect 590 1528 598 1531
rect 682 1528 686 1531
rect 462 1492 465 1508
rect 534 1492 537 1518
rect 590 1492 593 1528
rect 470 1482 473 1488
rect 482 1478 486 1481
rect 254 1472 257 1478
rect 310 1472 313 1478
rect 422 1472 425 1478
rect 550 1472 553 1488
rect 606 1472 609 1518
rect 686 1512 689 1528
rect 698 1518 702 1521
rect 306 1468 310 1471
rect 330 1458 334 1461
rect 242 1438 249 1441
rect 374 1442 377 1468
rect 422 1452 425 1458
rect 222 1352 225 1418
rect 198 1332 201 1348
rect 214 1342 217 1348
rect 230 1342 233 1418
rect 344 1403 346 1407
rect 350 1403 353 1407
rect 357 1403 360 1407
rect 446 1382 449 1458
rect 454 1452 457 1458
rect 254 1352 257 1358
rect 278 1342 281 1378
rect 430 1372 433 1378
rect 302 1362 305 1368
rect 310 1362 313 1368
rect 286 1352 289 1358
rect 310 1342 313 1358
rect 366 1352 369 1358
rect 382 1352 385 1358
rect 354 1348 358 1351
rect 390 1342 393 1368
rect 438 1362 441 1368
rect 426 1358 430 1361
rect 466 1358 470 1361
rect 490 1358 494 1361
rect 402 1348 406 1351
rect 362 1338 366 1341
rect 270 1332 273 1338
rect 414 1332 417 1358
rect 218 1328 225 1331
rect 214 1272 217 1318
rect 222 1312 225 1328
rect 314 1328 318 1331
rect 378 1328 382 1331
rect 230 1292 233 1328
rect 238 1292 241 1318
rect 290 1278 294 1281
rect 222 1262 225 1278
rect 238 1252 241 1268
rect 246 1262 249 1268
rect 246 1251 249 1258
rect 262 1252 265 1258
rect 246 1248 254 1251
rect 290 1248 294 1251
rect 158 1242 161 1248
rect 238 1232 241 1248
rect 22 1192 25 1198
rect 46 1192 49 1208
rect 158 1192 161 1228
rect 214 1192 217 1198
rect 122 1188 126 1191
rect 154 1168 158 1171
rect 90 1148 94 1151
rect 114 1148 118 1151
rect 126 1142 129 1158
rect 134 1152 137 1158
rect 142 1152 145 1168
rect 174 1162 177 1168
rect 166 1152 169 1158
rect 146 1148 150 1151
rect 6 1112 9 1128
rect 22 1122 25 1138
rect 6 1079 14 1081
rect 6 1078 17 1079
rect 6 1062 9 1078
rect 30 1042 33 1078
rect 38 1062 41 1068
rect 54 1042 57 1098
rect 78 1082 81 1138
rect 174 1132 177 1148
rect 190 1132 193 1138
rect 90 1128 94 1131
rect 86 1082 89 1088
rect 126 1072 129 1118
rect 182 1092 185 1108
rect 214 1082 217 1168
rect 246 1152 249 1248
rect 270 1242 273 1248
rect 262 1232 265 1238
rect 254 1162 257 1218
rect 234 1148 238 1151
rect 254 1142 257 1158
rect 286 1152 289 1178
rect 302 1172 305 1318
rect 310 1292 313 1308
rect 390 1292 393 1328
rect 310 1192 313 1208
rect 318 1192 321 1268
rect 326 1202 329 1258
rect 342 1242 345 1268
rect 350 1252 353 1278
rect 414 1272 417 1328
rect 446 1302 449 1348
rect 454 1322 457 1358
rect 462 1342 465 1348
rect 482 1338 486 1341
rect 478 1328 486 1331
rect 478 1292 481 1328
rect 494 1302 497 1318
rect 502 1292 505 1458
rect 558 1432 561 1468
rect 622 1442 625 1498
rect 718 1492 721 1528
rect 742 1502 745 1548
rect 766 1532 769 1548
rect 790 1542 793 1568
rect 810 1558 814 1561
rect 830 1552 833 1608
rect 878 1572 881 1598
rect 842 1558 846 1561
rect 886 1552 889 1628
rect 894 1562 897 1618
rect 902 1602 905 1648
rect 918 1612 921 1658
rect 942 1652 945 1668
rect 954 1658 958 1661
rect 966 1652 969 1678
rect 990 1672 993 1688
rect 1046 1682 1049 1708
rect 1142 1702 1145 1728
rect 974 1662 977 1668
rect 974 1642 977 1648
rect 1038 1642 1041 1668
rect 1050 1658 1054 1661
rect 1074 1658 1078 1661
rect 1106 1658 1110 1661
rect 1094 1652 1097 1658
rect 1134 1652 1137 1678
rect 1142 1662 1145 1668
rect 1158 1662 1161 1688
rect 1166 1672 1169 1708
rect 1182 1682 1185 1688
rect 1206 1662 1209 1688
rect 1214 1672 1217 1708
rect 1222 1692 1225 1698
rect 1170 1658 1174 1661
rect 1082 1648 1086 1651
rect 1062 1642 1065 1648
rect 1182 1642 1185 1648
rect 1074 1638 1078 1641
rect 966 1612 969 1618
rect 950 1592 953 1598
rect 998 1592 1001 1598
rect 1038 1582 1041 1638
rect 1102 1632 1105 1638
rect 1110 1632 1113 1638
rect 1126 1632 1129 1638
rect 962 1568 966 1571
rect 978 1568 982 1571
rect 1010 1568 1014 1571
rect 1058 1568 1062 1571
rect 898 1558 902 1561
rect 994 1558 998 1561
rect 1026 1558 1033 1561
rect 810 1548 814 1551
rect 866 1548 870 1551
rect 898 1548 902 1551
rect 910 1542 913 1558
rect 942 1552 945 1558
rect 1002 1548 1006 1551
rect 918 1542 921 1548
rect 926 1542 929 1548
rect 934 1542 937 1548
rect 950 1542 953 1548
rect 846 1532 849 1538
rect 982 1532 985 1548
rect 1022 1542 1025 1548
rect 1030 1532 1033 1558
rect 1046 1551 1049 1558
rect 1046 1548 1057 1551
rect 1042 1538 1046 1541
rect 1054 1532 1057 1548
rect 1070 1542 1073 1568
rect 1142 1562 1145 1568
rect 1206 1562 1209 1618
rect 1230 1552 1233 1768
rect 1350 1752 1353 1858
rect 1306 1738 1310 1741
rect 1254 1672 1257 1718
rect 1358 1692 1361 1928
rect 1382 1863 1385 1898
rect 1430 1892 1433 1908
rect 1438 1882 1441 1938
rect 1446 1922 1449 1938
rect 1510 1931 1513 1948
rect 1542 1942 1545 1948
rect 1522 1938 1526 1941
rect 1506 1928 1513 1931
rect 1534 1932 1537 1938
rect 1368 1803 1370 1807
rect 1374 1803 1377 1807
rect 1381 1803 1384 1807
rect 1430 1762 1433 1768
rect 1382 1742 1385 1747
rect 1422 1742 1425 1748
rect 1330 1678 1337 1681
rect 1326 1662 1329 1668
rect 1286 1652 1289 1659
rect 1322 1648 1326 1651
rect 1270 1592 1273 1648
rect 1334 1642 1337 1678
rect 1398 1672 1401 1718
rect 1402 1618 1406 1621
rect 1368 1603 1370 1607
rect 1374 1603 1377 1607
rect 1381 1603 1384 1607
rect 1122 1548 1126 1551
rect 1162 1548 1166 1551
rect 1322 1548 1326 1551
rect 1078 1542 1081 1548
rect 1086 1542 1089 1548
rect 1114 1538 1118 1541
rect 1146 1538 1150 1541
rect 1170 1538 1174 1541
rect 1314 1538 1318 1541
rect 1134 1532 1137 1538
rect 762 1528 766 1531
rect 1122 1528 1126 1531
rect 1138 1528 1142 1531
rect 782 1522 785 1528
rect 762 1488 766 1491
rect 646 1462 649 1468
rect 634 1458 638 1461
rect 642 1448 646 1451
rect 654 1451 657 1478
rect 686 1472 689 1478
rect 694 1472 697 1478
rect 726 1472 729 1488
rect 790 1482 793 1528
rect 856 1503 858 1507
rect 862 1503 865 1507
rect 869 1503 872 1507
rect 906 1488 910 1491
rect 1122 1488 1126 1491
rect 738 1478 742 1481
rect 774 1472 777 1478
rect 694 1462 697 1468
rect 734 1462 737 1468
rect 758 1462 761 1468
rect 862 1463 865 1468
rect 878 1462 881 1468
rect 990 1462 993 1468
rect 654 1448 662 1451
rect 662 1442 665 1448
rect 558 1362 561 1418
rect 614 1362 617 1418
rect 670 1362 673 1458
rect 758 1452 761 1458
rect 694 1442 697 1448
rect 974 1442 977 1459
rect 1026 1458 1030 1461
rect 1110 1462 1113 1468
rect 1094 1452 1097 1459
rect 794 1418 798 1421
rect 1026 1418 1030 1421
rect 602 1358 606 1361
rect 522 1348 526 1351
rect 546 1348 550 1351
rect 558 1342 561 1358
rect 578 1348 582 1351
rect 610 1348 614 1351
rect 630 1342 633 1358
rect 666 1348 670 1351
rect 686 1342 689 1398
rect 742 1342 745 1408
rect 1134 1402 1137 1528
rect 1158 1472 1161 1478
rect 1174 1392 1177 1518
rect 1206 1472 1209 1538
rect 1254 1532 1257 1538
rect 1290 1478 1294 1481
rect 1222 1472 1225 1478
rect 1242 1468 1246 1471
rect 1190 1463 1193 1468
rect 1182 1392 1185 1438
rect 1206 1392 1209 1468
rect 1238 1452 1241 1458
rect 1226 1448 1230 1451
rect 1250 1448 1254 1451
rect 1278 1442 1281 1478
rect 1302 1472 1305 1478
rect 1310 1462 1313 1468
rect 1294 1452 1297 1458
rect 1310 1442 1313 1448
rect 954 1368 958 1371
rect 970 1368 974 1371
rect 822 1362 825 1368
rect 810 1358 814 1361
rect 750 1342 753 1348
rect 518 1332 521 1338
rect 422 1262 425 1278
rect 430 1272 433 1288
rect 450 1278 454 1281
rect 498 1278 502 1281
rect 510 1272 513 1318
rect 550 1302 553 1338
rect 558 1322 561 1328
rect 582 1302 585 1338
rect 526 1282 529 1298
rect 562 1288 566 1291
rect 490 1268 494 1271
rect 454 1262 457 1268
rect 526 1262 529 1278
rect 590 1272 593 1278
rect 614 1272 617 1318
rect 622 1272 625 1328
rect 638 1292 641 1338
rect 694 1322 697 1338
rect 678 1292 681 1318
rect 702 1272 705 1318
rect 410 1258 414 1261
rect 358 1252 361 1258
rect 398 1242 401 1248
rect 406 1232 409 1248
rect 334 1192 337 1228
rect 344 1203 346 1207
rect 350 1203 353 1207
rect 357 1203 360 1207
rect 438 1182 441 1218
rect 462 1192 465 1258
rect 486 1242 489 1258
rect 302 1142 305 1168
rect 318 1162 321 1178
rect 282 1138 286 1141
rect 230 1132 233 1138
rect 230 1092 233 1128
rect 262 1112 265 1128
rect 270 1122 273 1128
rect 310 1112 313 1148
rect 406 1142 409 1158
rect 414 1152 417 1158
rect 438 1142 441 1158
rect 466 1148 470 1151
rect 486 1142 489 1228
rect 534 1172 537 1218
rect 510 1162 513 1168
rect 494 1142 497 1148
rect 358 1132 361 1138
rect 414 1132 417 1138
rect 542 1132 545 1268
rect 606 1192 609 1238
rect 614 1232 617 1258
rect 622 1192 625 1268
rect 670 1212 673 1268
rect 698 1258 705 1261
rect 702 1252 705 1258
rect 710 1252 713 1318
rect 766 1312 769 1318
rect 814 1292 817 1318
rect 822 1292 825 1338
rect 838 1322 841 1368
rect 846 1352 849 1368
rect 1006 1362 1009 1378
rect 1110 1372 1113 1378
rect 1018 1368 1025 1371
rect 1130 1368 1134 1371
rect 874 1358 881 1361
rect 856 1303 858 1307
rect 862 1303 865 1307
rect 869 1303 872 1307
rect 758 1282 761 1288
rect 766 1272 769 1278
rect 726 1262 729 1268
rect 734 1252 737 1258
rect 742 1252 745 1258
rect 750 1242 753 1268
rect 782 1262 785 1278
rect 830 1272 833 1278
rect 838 1272 841 1278
rect 774 1252 777 1258
rect 790 1251 793 1268
rect 846 1262 849 1278
rect 854 1272 857 1288
rect 802 1258 806 1261
rect 782 1248 793 1251
rect 714 1238 718 1241
rect 710 1192 713 1208
rect 622 1162 625 1178
rect 726 1162 729 1188
rect 762 1168 766 1171
rect 742 1162 745 1168
rect 554 1158 558 1161
rect 550 1142 553 1158
rect 562 1148 566 1151
rect 602 1148 606 1151
rect 646 1142 649 1148
rect 654 1142 657 1158
rect 678 1152 681 1158
rect 714 1148 718 1151
rect 738 1148 742 1151
rect 774 1142 777 1148
rect 566 1132 569 1138
rect 574 1132 577 1138
rect 582 1132 585 1138
rect 426 1128 430 1131
rect 326 1112 329 1128
rect 554 1118 558 1121
rect 374 1092 377 1118
rect 518 1092 521 1098
rect 466 1088 470 1091
rect 170 1078 174 1081
rect 62 1062 65 1068
rect 70 1052 73 1068
rect 142 1062 145 1078
rect 150 1072 153 1078
rect 214 1072 217 1078
rect 270 1072 273 1078
rect 278 1072 281 1088
rect 526 1082 529 1118
rect 122 1058 126 1061
rect 78 1052 81 1058
rect 150 1052 153 1058
rect 174 1052 177 1068
rect 194 1048 198 1051
rect 62 1032 65 1048
rect 102 1042 105 1048
rect 150 992 153 1048
rect 78 952 81 968
rect 22 931 25 948
rect 46 931 49 948
rect 70 931 73 948
rect 18 928 25 931
rect 42 928 49 931
rect 66 928 73 931
rect 110 892 113 928
rect 18 879 25 881
rect 14 878 25 879
rect 42 879 49 881
rect 38 878 49 879
rect 66 879 73 881
rect 62 878 73 879
rect 22 862 25 878
rect 46 862 49 878
rect 62 752 65 868
rect 70 862 73 878
rect 126 863 129 988
rect 138 958 142 961
rect 166 952 169 978
rect 198 962 201 978
rect 178 958 182 961
rect 198 952 201 958
rect 158 942 161 948
rect 194 938 198 941
rect 214 892 217 958
rect 222 952 225 1068
rect 278 1062 281 1068
rect 298 1058 302 1061
rect 242 1038 246 1041
rect 286 992 289 1058
rect 344 1003 346 1007
rect 350 1003 353 1007
rect 357 1003 360 1007
rect 242 968 246 971
rect 278 942 281 948
rect 222 932 225 938
rect 270 922 273 938
rect 302 932 305 978
rect 366 972 369 1068
rect 374 1062 377 1078
rect 390 1062 393 1078
rect 406 1072 409 1078
rect 470 1062 473 1068
rect 478 1062 481 1078
rect 514 1068 521 1071
rect 506 1058 513 1061
rect 382 992 385 998
rect 414 972 417 1058
rect 430 1052 433 1058
rect 446 1042 449 1058
rect 498 1048 502 1051
rect 438 992 441 1008
rect 394 958 398 961
rect 282 928 286 931
rect 202 888 206 891
rect 334 882 337 928
rect 158 862 161 868
rect 262 863 265 878
rect 366 872 369 948
rect 390 932 393 938
rect 390 892 393 918
rect 386 868 390 871
rect 278 862 281 868
rect 294 862 297 868
rect 358 842 361 868
rect 398 852 401 928
rect 406 882 409 948
rect 414 942 417 948
rect 422 932 425 958
rect 438 952 441 958
rect 454 942 457 1038
rect 478 982 481 1018
rect 466 968 470 971
rect 446 922 449 938
rect 438 918 446 921
rect 438 862 441 918
rect 446 892 449 898
rect 454 882 457 938
rect 470 902 473 948
rect 478 911 481 958
rect 494 942 497 1048
rect 510 1032 513 1058
rect 518 1002 521 1068
rect 542 1052 545 1058
rect 534 1022 537 1048
rect 550 1042 553 1108
rect 566 1062 569 1068
rect 562 1048 566 1051
rect 542 1032 545 1038
rect 506 968 510 971
rect 522 968 526 971
rect 502 912 505 928
rect 478 908 486 911
rect 446 872 449 878
rect 470 852 473 898
rect 486 872 489 908
rect 510 892 513 948
rect 526 942 529 968
rect 574 962 577 1118
rect 586 1068 590 1071
rect 582 1052 585 1058
rect 598 1012 601 1138
rect 630 1082 633 1118
rect 646 1082 649 1098
rect 654 1092 657 1138
rect 694 1132 697 1138
rect 702 1132 705 1138
rect 746 1128 750 1131
rect 662 1112 665 1118
rect 662 1072 665 1088
rect 642 1068 646 1071
rect 606 1062 609 1068
rect 622 1052 625 1068
rect 678 1062 681 1108
rect 634 1058 638 1061
rect 694 1052 697 1128
rect 758 1122 761 1128
rect 718 1082 721 1098
rect 702 1072 705 1078
rect 710 1072 713 1078
rect 734 1072 737 1078
rect 774 1072 777 1108
rect 782 1102 785 1248
rect 810 1188 814 1191
rect 810 1168 814 1171
rect 822 1162 825 1168
rect 830 1162 833 1258
rect 862 1252 865 1288
rect 878 1272 881 1358
rect 894 1342 897 1358
rect 918 1352 921 1358
rect 930 1338 934 1341
rect 970 1338 974 1341
rect 898 1328 902 1331
rect 954 1328 958 1331
rect 886 1312 889 1328
rect 886 1292 889 1308
rect 890 1278 894 1281
rect 902 1262 905 1268
rect 926 1212 929 1248
rect 790 1142 793 1158
rect 822 1152 825 1158
rect 830 1152 833 1158
rect 802 1148 806 1151
rect 902 1142 905 1188
rect 934 1182 937 1318
rect 942 1302 945 1328
rect 982 1282 985 1348
rect 990 1322 993 1358
rect 998 1332 1001 1358
rect 1010 1348 1014 1351
rect 1022 1342 1025 1368
rect 1034 1358 1038 1361
rect 1058 1358 1062 1361
rect 1146 1358 1150 1361
rect 1070 1352 1073 1358
rect 1046 1342 1049 1348
rect 1054 1342 1057 1348
rect 1086 1342 1089 1358
rect 1130 1348 1134 1351
rect 1170 1348 1174 1351
rect 1074 1338 1078 1341
rect 1122 1338 1126 1341
rect 1178 1338 1182 1341
rect 1086 1332 1089 1338
rect 1142 1332 1145 1338
rect 1262 1332 1265 1338
rect 954 1278 958 1281
rect 986 1278 990 1281
rect 942 1262 945 1278
rect 966 1272 969 1278
rect 998 1272 1001 1328
rect 1150 1322 1153 1328
rect 1014 1272 1017 1318
rect 1030 1311 1033 1318
rect 1022 1308 1033 1311
rect 1022 1282 1025 1308
rect 1030 1292 1033 1298
rect 1086 1282 1089 1288
rect 1182 1282 1185 1318
rect 1178 1278 1182 1281
rect 998 1262 1001 1268
rect 1022 1262 1025 1278
rect 1062 1272 1065 1278
rect 1050 1268 1054 1271
rect 1090 1268 1094 1271
rect 1118 1262 1121 1268
rect 966 1212 969 1258
rect 990 1202 993 1258
rect 1002 1248 1006 1251
rect 1030 1202 1033 1248
rect 1054 1191 1057 1248
rect 1062 1202 1065 1258
rect 1126 1252 1129 1278
rect 1134 1252 1137 1268
rect 1142 1252 1145 1258
rect 1142 1242 1145 1248
rect 1070 1232 1073 1238
rect 1150 1232 1153 1238
rect 1190 1232 1193 1328
rect 1266 1318 1270 1321
rect 1206 1272 1209 1288
rect 1226 1278 1230 1281
rect 1198 1262 1201 1268
rect 1206 1252 1209 1258
rect 1214 1251 1217 1278
rect 1222 1272 1225 1278
rect 1254 1272 1257 1288
rect 1278 1262 1281 1308
rect 1310 1292 1313 1428
rect 1318 1342 1321 1538
rect 1334 1482 1337 1588
rect 1446 1551 1449 1908
rect 1554 1888 1558 1891
rect 1574 1872 1577 1918
rect 1598 1912 1601 1938
rect 1606 1892 1609 1898
rect 1646 1892 1649 2108
rect 1654 2082 1657 2098
rect 1686 2062 1689 2138
rect 1694 2122 1697 2158
rect 1706 2148 1710 2151
rect 1730 2148 1734 2151
rect 1718 2142 1721 2148
rect 1694 2072 1697 2118
rect 1702 2092 1705 2138
rect 1742 2082 1745 2158
rect 1814 2152 1817 2378
rect 1822 2372 1825 2438
rect 1830 2392 1833 2548
rect 1886 2542 1889 2547
rect 1872 2503 1874 2507
rect 1878 2503 1881 2507
rect 1885 2503 1888 2507
rect 1966 2492 1969 2578
rect 1974 2492 1977 2618
rect 2014 2492 2017 2618
rect 2110 2552 2113 2628
rect 2142 2592 2145 2598
rect 2206 2592 2209 2608
rect 2270 2582 2273 2588
rect 2022 2542 2025 2547
rect 2038 2492 2041 2548
rect 2078 2542 2081 2547
rect 2166 2531 2169 2548
rect 2162 2528 2169 2531
rect 2206 2531 2209 2558
rect 2334 2552 2337 2628
rect 2238 2542 2241 2548
rect 2306 2547 2310 2550
rect 2218 2538 2222 2541
rect 2254 2532 2257 2538
rect 2206 2528 2214 2531
rect 2198 2511 2201 2528
rect 2246 2522 2249 2528
rect 2358 2522 2361 2648
rect 2366 2592 2369 2648
rect 2190 2508 2201 2511
rect 2134 2492 2137 2498
rect 2158 2492 2161 2498
rect 1854 2462 1857 2468
rect 1882 2459 1886 2462
rect 1926 2402 1929 2418
rect 1918 2381 1921 2398
rect 1926 2392 1929 2398
rect 1918 2378 1929 2381
rect 1822 2352 1825 2368
rect 1830 2352 1833 2378
rect 1838 2352 1841 2358
rect 1846 2352 1849 2368
rect 1830 2282 1833 2348
rect 1854 2342 1857 2348
rect 1886 2342 1889 2368
rect 1918 2362 1921 2368
rect 1898 2348 1902 2351
rect 1914 2348 1918 2351
rect 1854 2292 1857 2338
rect 1902 2332 1905 2348
rect 1926 2332 1929 2378
rect 1934 2352 1937 2478
rect 1998 2472 2001 2478
rect 1942 2382 1945 2418
rect 1966 2402 1969 2448
rect 1942 2362 1945 2378
rect 1966 2372 1969 2398
rect 1974 2362 1977 2448
rect 1982 2392 1985 2398
rect 1990 2382 1993 2468
rect 2014 2452 2017 2468
rect 2022 2462 2025 2468
rect 2038 2452 2041 2468
rect 2102 2462 2105 2478
rect 2158 2472 2161 2478
rect 2146 2468 2150 2471
rect 2070 2452 2073 2459
rect 2094 2458 2102 2461
rect 2010 2448 2014 2451
rect 2006 2392 2009 2418
rect 2006 2372 2009 2378
rect 1998 2362 2001 2368
rect 1954 2358 1958 2361
rect 2006 2352 2009 2368
rect 1874 2328 1878 2331
rect 1862 2322 1865 2328
rect 1872 2303 1874 2307
rect 1878 2303 1881 2307
rect 1885 2303 1888 2307
rect 1878 2282 1881 2288
rect 1866 2268 1870 2271
rect 1882 2268 1886 2271
rect 1830 2192 1833 2248
rect 1838 2151 1841 2218
rect 1846 2192 1849 2268
rect 1874 2258 1878 2261
rect 1886 2162 1889 2218
rect 1894 2152 1897 2328
rect 1942 2322 1945 2338
rect 1902 2312 1905 2318
rect 1902 2252 1905 2308
rect 1926 2292 1929 2318
rect 1918 2242 1921 2268
rect 1934 2172 1937 2308
rect 1950 2302 1953 2348
rect 1966 2312 1969 2348
rect 1966 2292 1969 2298
rect 1942 2262 1945 2268
rect 1950 2232 1953 2278
rect 1958 2192 1961 2288
rect 2006 2272 2009 2328
rect 2014 2312 2017 2358
rect 2022 2278 2025 2358
rect 2030 2342 2033 2348
rect 2030 2322 2033 2328
rect 2062 2322 2065 2347
rect 2078 2292 2081 2368
rect 2094 2352 2097 2458
rect 2090 2278 2094 2281
rect 2110 2272 2113 2278
rect 2098 2268 2102 2271
rect 1994 2258 1998 2261
rect 2054 2252 2057 2268
rect 2062 2262 2065 2268
rect 2070 2262 2073 2268
rect 2118 2261 2121 2448
rect 2158 2412 2161 2448
rect 2190 2442 2193 2508
rect 2198 2452 2201 2458
rect 2222 2452 2225 2458
rect 2126 2392 2129 2398
rect 2166 2392 2169 2418
rect 2190 2392 2193 2438
rect 2246 2392 2249 2508
rect 2254 2492 2257 2498
rect 2262 2482 2265 2518
rect 2286 2472 2289 2478
rect 2126 2292 2129 2378
rect 2218 2348 2222 2351
rect 2186 2338 2190 2341
rect 2210 2338 2214 2341
rect 2234 2338 2241 2341
rect 2150 2292 2153 2332
rect 2186 2328 2190 2331
rect 2218 2328 2222 2331
rect 2182 2292 2185 2328
rect 2238 2312 2241 2338
rect 2254 2292 2257 2318
rect 2110 2258 2121 2261
rect 1974 2232 1977 2248
rect 2022 2242 2025 2248
rect 1962 2168 1966 2171
rect 1654 2052 1657 2059
rect 1686 2042 1689 2058
rect 1726 2052 1729 2078
rect 1750 2052 1753 2128
rect 1758 2122 1761 2128
rect 1758 2072 1761 2078
rect 1766 2072 1769 2088
rect 1774 2082 1777 2118
rect 1814 2102 1817 2148
rect 1934 2142 1937 2168
rect 1942 2142 1945 2148
rect 1902 2138 1910 2141
rect 1950 2141 1953 2158
rect 1946 2138 1953 2141
rect 1878 2132 1881 2138
rect 1872 2103 1874 2107
rect 1878 2103 1881 2107
rect 1885 2103 1888 2107
rect 1846 2082 1849 2098
rect 1782 2062 1785 2078
rect 1850 2068 1854 2071
rect 1894 2071 1897 2138
rect 1902 2092 1905 2138
rect 1918 2092 1921 2128
rect 1958 2092 1961 2148
rect 1910 2082 1913 2088
rect 1926 2082 1929 2088
rect 1990 2082 1993 2198
rect 2070 2192 2073 2198
rect 2078 2192 2081 2208
rect 2102 2182 2105 2258
rect 2010 2147 2014 2150
rect 2006 2132 2009 2138
rect 2086 2132 2089 2138
rect 1998 2092 2001 2108
rect 2062 2092 2065 2118
rect 2094 2112 2097 2128
rect 2110 2092 2113 2258
rect 2134 2252 2137 2278
rect 2198 2272 2201 2288
rect 2246 2272 2249 2278
rect 2146 2248 2150 2251
rect 2134 2241 2137 2248
rect 2134 2238 2145 2241
rect 2130 2208 2137 2211
rect 2134 2192 2137 2208
rect 2142 2172 2145 2238
rect 2150 2202 2153 2218
rect 2158 2202 2161 2268
rect 2186 2258 2190 2261
rect 2226 2258 2230 2261
rect 2174 2242 2177 2248
rect 2178 2238 2182 2241
rect 2190 2212 2193 2248
rect 2222 2222 2225 2248
rect 2174 2192 2177 2208
rect 2222 2192 2225 2218
rect 2122 2168 2126 2171
rect 2146 2148 2150 2151
rect 2118 2142 2121 2148
rect 2142 2132 2145 2138
rect 2158 2132 2161 2158
rect 2182 2152 2185 2158
rect 2174 2122 2177 2148
rect 2206 2132 2209 2138
rect 2214 2132 2217 2158
rect 2246 2132 2249 2258
rect 2262 2252 2265 2468
rect 2302 2452 2305 2468
rect 2318 2452 2321 2459
rect 2350 2452 2353 2458
rect 2302 2352 2305 2448
rect 2342 2392 2345 2398
rect 2374 2372 2377 2538
rect 2382 2492 2385 2638
rect 2392 2603 2394 2607
rect 2398 2603 2401 2607
rect 2405 2603 2408 2607
rect 2414 2561 2417 2648
rect 2438 2632 2441 2668
rect 2454 2652 2457 2659
rect 2422 2592 2425 2628
rect 2502 2582 2505 2858
rect 2526 2821 2529 2858
rect 2526 2818 2537 2821
rect 2518 2792 2521 2808
rect 2510 2592 2513 2748
rect 2518 2692 2521 2768
rect 2534 2742 2537 2818
rect 2550 2742 2553 2747
rect 2570 2688 2577 2691
rect 2526 2672 2529 2678
rect 2574 2672 2577 2688
rect 2582 2682 2585 2748
rect 2598 2692 2601 2858
rect 2622 2822 2625 2868
rect 2630 2862 2633 2868
rect 2646 2852 2649 2868
rect 2630 2842 2633 2848
rect 2654 2822 2657 2878
rect 2790 2872 2793 2878
rect 2682 2868 2686 2871
rect 2738 2868 2742 2871
rect 2666 2858 2670 2861
rect 2690 2848 2694 2851
rect 2718 2851 2721 2868
rect 2738 2858 2742 2861
rect 2718 2848 2726 2851
rect 2678 2842 2681 2848
rect 2686 2832 2689 2838
rect 2726 2812 2729 2848
rect 2750 2822 2753 2868
rect 2774 2862 2777 2868
rect 2790 2852 2793 2868
rect 2814 2862 2817 2868
rect 2822 2862 2825 2918
rect 2838 2862 2841 2918
rect 2854 2892 2857 2928
rect 2894 2912 2897 2968
rect 2958 2952 2961 2988
rect 2938 2948 2942 2951
rect 3038 2942 3041 2958
rect 3010 2938 3017 2941
rect 2904 2903 2906 2907
rect 2910 2903 2913 2907
rect 2917 2903 2920 2907
rect 2942 2892 2945 2938
rect 2998 2872 3001 2888
rect 3006 2872 3009 2878
rect 2914 2868 2918 2871
rect 2762 2838 2766 2841
rect 2774 2832 2777 2848
rect 2830 2842 2833 2848
rect 2846 2842 2849 2868
rect 2862 2842 2865 2868
rect 2794 2838 2798 2841
rect 2810 2838 2814 2841
rect 2870 2832 2873 2858
rect 2878 2852 2881 2868
rect 2926 2862 2929 2868
rect 2894 2852 2897 2858
rect 2918 2852 2921 2858
rect 2966 2852 2969 2868
rect 2978 2858 2982 2861
rect 2942 2842 2945 2848
rect 2614 2792 2617 2798
rect 2702 2792 2705 2808
rect 2626 2778 2630 2781
rect 2634 2738 2638 2741
rect 2690 2738 2694 2741
rect 2698 2728 2702 2731
rect 2726 2731 2729 2748
rect 2734 2742 2737 2758
rect 2782 2742 2785 2798
rect 2858 2768 2862 2771
rect 2830 2762 2833 2768
rect 2886 2762 2889 2838
rect 2950 2832 2953 2848
rect 2974 2832 2977 2848
rect 2894 2792 2897 2828
rect 2990 2792 2993 2848
rect 2998 2811 3001 2858
rect 3014 2852 3017 2938
rect 3046 2932 3049 2948
rect 3038 2912 3041 2918
rect 3054 2892 3057 3008
rect 3078 2982 3081 3068
rect 3098 3058 3102 3061
rect 3134 3002 3137 3058
rect 3122 2988 3126 2991
rect 3122 2958 3126 2961
rect 3070 2952 3073 2958
rect 3086 2952 3089 2958
rect 3066 2938 3070 2941
rect 3086 2892 3089 2928
rect 3102 2902 3105 2948
rect 3134 2942 3137 2958
rect 3142 2952 3145 3078
rect 3158 3072 3161 3118
rect 3214 3112 3217 3128
rect 3262 3092 3265 3098
rect 3278 3092 3281 3138
rect 3286 3111 3289 3218
rect 3342 3212 3345 3218
rect 3294 3152 3297 3158
rect 3330 3148 3334 3151
rect 3358 3142 3361 3148
rect 3330 3138 3334 3141
rect 3302 3121 3305 3138
rect 3374 3132 3377 3308
rect 3414 3281 3417 3332
rect 3458 3328 3462 3331
rect 3422 3292 3425 3298
rect 3414 3278 3425 3281
rect 3394 3268 3398 3271
rect 3410 3268 3414 3271
rect 3382 3222 3385 3258
rect 3422 3252 3425 3278
rect 3430 3252 3433 3328
rect 3446 3262 3449 3318
rect 3494 3272 3497 3348
rect 3510 3322 3513 3328
rect 3458 3268 3462 3271
rect 3442 3258 3446 3261
rect 3470 3258 3478 3261
rect 3430 3232 3433 3248
rect 3382 3152 3385 3208
rect 3416 3203 3418 3207
rect 3422 3203 3425 3207
rect 3429 3203 3432 3207
rect 3462 3172 3465 3248
rect 3298 3118 3305 3121
rect 3286 3108 3297 3111
rect 3214 3088 3222 3091
rect 3214 3072 3217 3088
rect 3206 3062 3209 3068
rect 3222 3052 3225 3058
rect 3238 3052 3241 3088
rect 3286 3082 3289 3098
rect 3294 3082 3297 3108
rect 3310 3082 3313 3118
rect 3318 3082 3321 3108
rect 3266 3058 3270 3061
rect 3186 3048 3190 3051
rect 3266 3048 3270 3051
rect 3262 3042 3265 3048
rect 3206 2992 3209 2998
rect 3170 2958 3174 2961
rect 3222 2952 3225 2958
rect 3142 2942 3145 2948
rect 3150 2942 3153 2948
rect 3190 2942 3193 2948
rect 3130 2888 3134 2891
rect 3122 2878 3126 2881
rect 3026 2868 3030 2871
rect 3134 2871 3137 2878
rect 3126 2868 3137 2871
rect 3142 2872 3145 2918
rect 3150 2892 3153 2938
rect 3230 2932 3233 2968
rect 3238 2952 3241 3038
rect 3254 2942 3257 2968
rect 3262 2952 3265 3028
rect 3278 2962 3281 2978
rect 3294 2972 3297 3078
rect 3318 3072 3321 3078
rect 3326 3062 3329 3068
rect 3310 3032 3313 3058
rect 3342 3052 3345 3118
rect 3366 3092 3369 3128
rect 3382 3122 3385 3148
rect 3406 3132 3409 3168
rect 3470 3162 3473 3258
rect 3478 3242 3481 3248
rect 3486 3232 3489 3268
rect 3498 3258 3502 3261
rect 3494 3242 3497 3248
rect 3510 3192 3513 3268
rect 3542 3252 3545 3259
rect 3550 3192 3553 3288
rect 3566 3272 3569 3338
rect 3654 3332 3657 3338
rect 3606 3292 3609 3298
rect 3654 3272 3657 3328
rect 3574 3262 3577 3268
rect 3654 3262 3657 3268
rect 3638 3242 3641 3259
rect 3702 3252 3705 3348
rect 3710 3262 3713 3348
rect 3718 3312 3721 3318
rect 3766 3312 3769 3398
rect 3742 3262 3745 3308
rect 3766 3282 3769 3308
rect 3774 3292 3777 3348
rect 3782 3322 3785 3478
rect 3830 3462 3833 3478
rect 3838 3472 3841 3478
rect 3886 3462 3889 3518
rect 3902 3512 3905 3548
rect 3910 3492 3913 3568
rect 3950 3552 3953 3638
rect 3982 3551 3985 3558
rect 4006 3552 4009 3638
rect 4046 3582 4049 3588
rect 3922 3538 3926 3541
rect 3918 3482 3921 3528
rect 3928 3503 3930 3507
rect 3934 3503 3937 3507
rect 3941 3503 3944 3507
rect 3950 3472 3953 3548
rect 4058 3538 4062 3541
rect 3966 3472 3969 3538
rect 4070 3492 4073 3618
rect 4094 3552 4097 3558
rect 4102 3552 4105 3578
rect 4086 3542 4089 3548
rect 4110 3492 4113 3648
rect 4118 3592 4121 3728
rect 4198 3728 4202 3732
rect 4214 3728 4218 3732
rect 4238 3728 4242 3732
rect 4294 3728 4298 3732
rect 4342 3728 4346 3732
rect 4358 3728 4362 3732
rect 4374 3728 4378 3732
rect 4430 3731 4434 3732
rect 4582 3731 4586 3732
rect 4766 3731 4770 3732
rect 4430 3728 4441 3731
rect 4582 3728 4593 3731
rect 4766 3728 4777 3731
rect 4182 3682 4185 3688
rect 4190 3672 4193 3678
rect 4174 3662 4177 3668
rect 4182 3652 4185 3658
rect 4134 3582 4137 3588
rect 4174 3552 4177 3558
rect 4166 3542 4169 3548
rect 4182 3542 4185 3578
rect 4190 3542 4193 3548
rect 4198 3541 4201 3728
rect 4214 3702 4217 3728
rect 4238 3702 4241 3728
rect 4294 3702 4297 3728
rect 4342 3692 4345 3728
rect 4334 3688 4342 3691
rect 4302 3672 4305 3688
rect 4238 3652 4241 3659
rect 4246 3642 4249 3668
rect 4246 3592 4249 3638
rect 4310 3572 4313 3678
rect 4334 3672 4337 3688
rect 4358 3671 4361 3728
rect 4374 3702 4377 3728
rect 4438 3692 4441 3728
rect 4590 3692 4593 3728
rect 4774 3692 4777 3728
rect 4862 3728 4866 3732
rect 4886 3731 4890 3732
rect 4878 3728 4890 3731
rect 5174 3731 5178 3732
rect 5222 3731 5226 3732
rect 5174 3728 5185 3731
rect 5222 3728 5233 3731
rect 4354 3668 4361 3671
rect 4326 3662 4329 3668
rect 4350 3642 4353 3668
rect 4366 3662 4369 3668
rect 4374 3662 4377 3688
rect 4710 3682 4713 3688
rect 4722 3678 4726 3681
rect 4358 3652 4361 3658
rect 4350 3572 4353 3618
rect 4374 3582 4377 3658
rect 4390 3642 4393 3658
rect 4398 3652 4401 3658
rect 4414 3632 4417 3678
rect 4446 3672 4449 3678
rect 4562 3668 4566 3671
rect 4422 3662 4425 3668
rect 4510 3662 4513 3668
rect 4534 3662 4537 3668
rect 4662 3663 4665 3678
rect 4706 3668 4710 3671
rect 4426 3658 4430 3661
rect 4450 3658 4454 3661
rect 4390 3592 4393 3618
rect 4378 3568 4382 3571
rect 4310 3562 4313 3568
rect 4226 3558 4230 3561
rect 4310 3552 4313 3558
rect 4210 3548 4214 3551
rect 4194 3538 4201 3541
rect 4322 3538 4326 3541
rect 4126 3532 4129 3538
rect 4058 3478 4062 3481
rect 4110 3472 4113 3488
rect 3858 3458 3862 3461
rect 4038 3462 4041 3468
rect 3798 3432 3801 3458
rect 3846 3361 3849 3428
rect 3886 3372 3889 3458
rect 3950 3392 3953 3448
rect 3974 3421 3977 3459
rect 3974 3418 3985 3421
rect 3846 3358 3854 3361
rect 3814 3352 3817 3358
rect 3846 3352 3849 3358
rect 3886 3352 3889 3368
rect 3922 3348 3926 3351
rect 3798 3332 3801 3338
rect 3782 3262 3785 3318
rect 3822 3302 3825 3348
rect 3854 3342 3857 3348
rect 3842 3338 3846 3341
rect 3906 3338 3910 3341
rect 3914 3328 3918 3331
rect 3846 3292 3849 3298
rect 3834 3279 3841 3281
rect 3830 3278 3841 3279
rect 3838 3262 3841 3278
rect 3894 3272 3897 3328
rect 3718 3242 3721 3258
rect 3706 3238 3710 3241
rect 3506 3168 3510 3171
rect 3534 3162 3537 3168
rect 3558 3162 3561 3228
rect 3614 3192 3617 3238
rect 3758 3192 3761 3248
rect 3574 3162 3577 3168
rect 3426 3158 3430 3161
rect 3562 3158 3566 3161
rect 3602 3158 3606 3161
rect 3442 3148 3446 3151
rect 3458 3148 3462 3151
rect 3434 3138 3438 3141
rect 3438 3132 3441 3138
rect 3446 3122 3449 3148
rect 3470 3132 3473 3158
rect 3494 3152 3497 3158
rect 3486 3142 3489 3148
rect 3558 3142 3561 3148
rect 3514 3138 3518 3141
rect 3362 3078 3366 3081
rect 3350 3072 3353 3078
rect 3370 3068 3374 3071
rect 3350 3042 3353 3048
rect 3366 3042 3369 3048
rect 3302 2962 3305 3018
rect 3326 2982 3329 3018
rect 3382 2992 3385 3118
rect 3450 3078 3454 3081
rect 3398 3062 3401 3068
rect 3406 3052 3409 3068
rect 3430 3052 3433 3078
rect 3462 3072 3465 3078
rect 3402 3048 3406 3051
rect 3438 3042 3441 3058
rect 3462 3042 3465 3048
rect 3394 3038 3398 3041
rect 3450 3038 3454 3041
rect 3310 2972 3313 2978
rect 3354 2968 3358 2971
rect 3342 2962 3345 2968
rect 3374 2962 3377 2978
rect 3282 2958 3289 2961
rect 3286 2942 3289 2958
rect 3302 2952 3305 2958
rect 3326 2952 3329 2958
rect 3358 2942 3361 2948
rect 3338 2938 3342 2941
rect 3214 2912 3217 2928
rect 3078 2862 3081 2868
rect 3106 2858 3110 2861
rect 3046 2852 3049 2858
rect 3126 2852 3129 2868
rect 3138 2858 3142 2861
rect 3018 2848 3022 2851
rect 3086 2842 3089 2848
rect 2998 2808 3009 2811
rect 2958 2772 2961 2778
rect 2906 2768 2910 2771
rect 2994 2768 2998 2771
rect 2794 2758 2798 2761
rect 2826 2758 2830 2761
rect 2842 2758 2846 2761
rect 2870 2752 2873 2758
rect 2878 2752 2881 2758
rect 2810 2748 2814 2751
rect 2790 2742 2793 2748
rect 2830 2742 2833 2748
rect 2630 2682 2633 2728
rect 2722 2728 2729 2731
rect 2638 2682 2641 2698
rect 2554 2658 2558 2661
rect 2518 2592 2521 2598
rect 2410 2558 2417 2561
rect 2402 2538 2406 2541
rect 2414 2452 2417 2468
rect 2392 2403 2394 2407
rect 2398 2403 2401 2407
rect 2405 2403 2408 2407
rect 2366 2352 2369 2358
rect 2414 2352 2417 2448
rect 2278 2342 2281 2347
rect 2286 2272 2289 2278
rect 2350 2272 2353 2338
rect 2362 2328 2366 2331
rect 2374 2331 2377 2348
rect 2398 2332 2401 2348
rect 2430 2342 2433 2459
rect 2478 2412 2481 2538
rect 2486 2532 2489 2558
rect 2550 2548 2558 2551
rect 2494 2532 2497 2538
rect 2494 2492 2497 2498
rect 2550 2492 2553 2548
rect 2558 2492 2561 2518
rect 2582 2502 2585 2668
rect 2654 2662 2657 2718
rect 2662 2692 2665 2718
rect 2754 2688 2758 2691
rect 2698 2658 2702 2661
rect 2742 2632 2745 2668
rect 2790 2662 2793 2728
rect 2806 2712 2809 2738
rect 2838 2732 2841 2748
rect 2854 2712 2857 2728
rect 2854 2672 2857 2708
rect 2598 2542 2601 2628
rect 2790 2622 2793 2658
rect 2654 2592 2657 2608
rect 2662 2592 2665 2598
rect 2618 2568 2622 2571
rect 2726 2542 2729 2547
rect 2622 2502 2625 2528
rect 2630 2512 2633 2528
rect 2518 2472 2521 2478
rect 2622 2452 2625 2459
rect 2522 2448 2526 2451
rect 2514 2438 2518 2441
rect 2526 2422 2529 2438
rect 2550 2422 2553 2448
rect 2478 2342 2481 2408
rect 2574 2352 2577 2438
rect 2610 2388 2614 2391
rect 2506 2348 2510 2351
rect 2374 2328 2382 2331
rect 2374 2282 2377 2298
rect 2398 2292 2401 2328
rect 2370 2278 2374 2281
rect 2362 2268 2366 2271
rect 2454 2262 2457 2288
rect 2462 2272 2465 2278
rect 2494 2272 2497 2318
rect 2514 2268 2518 2271
rect 2298 2258 2302 2261
rect 2402 2248 2406 2251
rect 2254 2242 2257 2248
rect 2514 2238 2518 2241
rect 2254 2132 2257 2178
rect 2270 2152 2273 2188
rect 2302 2152 2305 2218
rect 2358 2162 2361 2228
rect 2392 2203 2394 2207
rect 2398 2203 2401 2207
rect 2405 2203 2408 2207
rect 2382 2191 2385 2198
rect 2502 2192 2505 2218
rect 2382 2188 2390 2191
rect 2434 2158 2438 2161
rect 2450 2158 2454 2161
rect 2326 2152 2329 2158
rect 2358 2151 2361 2158
rect 2470 2152 2473 2158
rect 2286 2142 2289 2148
rect 2270 2132 2273 2138
rect 2258 2128 2262 2131
rect 2190 2092 2193 2098
rect 2126 2088 2134 2091
rect 2074 2078 2078 2081
rect 1890 2068 1897 2071
rect 1930 2068 1934 2071
rect 1798 2052 1801 2058
rect 1770 2048 1774 2051
rect 1718 2022 1721 2028
rect 1734 2012 1737 2018
rect 1666 1958 1670 1961
rect 1686 1952 1689 1978
rect 1654 1932 1657 1938
rect 1702 1932 1705 1968
rect 1718 1942 1721 1978
rect 1742 1972 1745 2038
rect 1782 2032 1785 2048
rect 1822 2042 1825 2048
rect 1810 2038 1814 2041
rect 1838 2032 1841 2068
rect 1858 2048 1862 2051
rect 1774 1972 1777 1978
rect 1742 1962 1745 1968
rect 1790 1952 1793 2028
rect 1806 1992 1809 2018
rect 1814 2012 1817 2018
rect 1838 1972 1841 1978
rect 1730 1948 1734 1951
rect 1746 1948 1750 1951
rect 1770 1948 1774 1951
rect 1746 1938 1750 1941
rect 1702 1892 1705 1918
rect 1750 1912 1753 1928
rect 1798 1901 1801 1938
rect 1818 1928 1822 1931
rect 1798 1898 1806 1901
rect 1718 1892 1721 1898
rect 1830 1892 1833 1968
rect 1846 1962 1849 2008
rect 1866 1958 1870 1961
rect 1886 1951 1889 2068
rect 1918 2012 1921 2018
rect 1894 1962 1897 2008
rect 1926 2002 1929 2008
rect 1926 1992 1929 1998
rect 1886 1948 1897 1951
rect 1838 1942 1841 1948
rect 1842 1938 1854 1941
rect 1862 1891 1865 1918
rect 1872 1903 1874 1907
rect 1878 1903 1881 1907
rect 1885 1903 1888 1907
rect 1862 1888 1873 1891
rect 1582 1882 1585 1888
rect 1614 1882 1617 1888
rect 1666 1879 1673 1881
rect 1662 1878 1673 1879
rect 1598 1872 1601 1878
rect 1618 1868 1622 1871
rect 1462 1752 1465 1858
rect 1494 1852 1497 1859
rect 1526 1842 1529 1868
rect 1670 1862 1673 1878
rect 1678 1862 1681 1868
rect 1594 1858 1598 1861
rect 1462 1742 1465 1748
rect 1462 1542 1465 1668
rect 1470 1663 1473 1828
rect 1582 1792 1585 1838
rect 1542 1762 1545 1778
rect 1494 1751 1497 1758
rect 1542 1752 1545 1758
rect 1598 1742 1601 1818
rect 1606 1792 1609 1848
rect 1630 1782 1633 1858
rect 1686 1852 1689 1858
rect 1670 1742 1673 1848
rect 1686 1792 1689 1798
rect 1710 1792 1713 1878
rect 1766 1872 1769 1888
rect 1730 1868 1734 1871
rect 1754 1868 1758 1871
rect 1826 1868 1830 1871
rect 1742 1862 1745 1868
rect 1734 1851 1737 1858
rect 1734 1848 1745 1851
rect 1742 1792 1745 1848
rect 1750 1801 1753 1848
rect 1758 1812 1761 1848
rect 1750 1798 1761 1801
rect 1718 1781 1721 1788
rect 1710 1778 1721 1781
rect 1694 1762 1697 1768
rect 1678 1752 1681 1758
rect 1702 1752 1705 1758
rect 1710 1752 1713 1778
rect 1718 1762 1721 1768
rect 1718 1752 1721 1758
rect 1734 1752 1737 1758
rect 1614 1702 1617 1728
rect 1502 1692 1505 1698
rect 1638 1692 1641 1732
rect 1618 1688 1622 1691
rect 1658 1678 1662 1681
rect 1486 1672 1489 1678
rect 1670 1672 1673 1678
rect 1650 1668 1654 1671
rect 1534 1662 1537 1668
rect 1598 1662 1601 1668
rect 1486 1592 1489 1648
rect 1494 1552 1497 1618
rect 1534 1572 1537 1658
rect 1566 1602 1569 1659
rect 1674 1658 1678 1661
rect 1690 1658 1694 1661
rect 1678 1642 1681 1648
rect 1702 1592 1705 1728
rect 1758 1692 1761 1798
rect 1766 1732 1769 1858
rect 1838 1852 1841 1888
rect 1870 1878 1873 1888
rect 1866 1818 1870 1821
rect 1778 1758 1782 1761
rect 1766 1722 1769 1728
rect 1782 1702 1785 1728
rect 1790 1712 1793 1818
rect 1894 1792 1897 1948
rect 1910 1942 1913 1948
rect 1942 1942 1945 1948
rect 1938 1938 1942 1941
rect 1902 1922 1905 1938
rect 1918 1912 1921 1938
rect 1926 1922 1929 1928
rect 1934 1872 1937 1888
rect 1950 1872 1953 1978
rect 1982 1952 1985 2068
rect 1990 2042 1993 2078
rect 2006 2072 2009 2078
rect 2094 2072 2097 2078
rect 2126 2072 2129 2088
rect 2042 2068 2046 2071
rect 2086 2062 2089 2068
rect 2118 2062 2121 2068
rect 2174 2062 2177 2068
rect 2198 2062 2201 2068
rect 2022 2052 2025 2058
rect 2098 2048 2102 2051
rect 2186 2048 2190 2051
rect 2146 2028 2150 2031
rect 2230 2022 2233 2059
rect 2246 2042 2249 2128
rect 2266 2118 2270 2121
rect 2290 2118 2294 2121
rect 2302 2092 2305 2148
rect 2414 2142 2417 2148
rect 2446 2142 2449 2148
rect 2462 2142 2465 2148
rect 2426 2138 2430 2141
rect 2398 2122 2401 2138
rect 2478 2132 2481 2168
rect 2534 2142 2537 2308
rect 2542 2131 2545 2347
rect 2534 2128 2545 2131
rect 2558 2152 2561 2158
rect 2566 2152 2569 2279
rect 2590 2272 2593 2388
rect 2622 2292 2625 2368
rect 2638 2351 2641 2538
rect 2710 2462 2713 2538
rect 2742 2492 2745 2618
rect 2758 2542 2761 2548
rect 2798 2542 2801 2588
rect 2778 2538 2782 2541
rect 2790 2532 2793 2538
rect 2782 2522 2785 2528
rect 2750 2482 2753 2508
rect 2774 2492 2777 2508
rect 2678 2452 2681 2459
rect 2710 2382 2713 2458
rect 2670 2352 2673 2378
rect 2734 2351 2737 2358
rect 2646 2332 2649 2348
rect 2686 2272 2689 2278
rect 2690 2268 2694 2271
rect 2574 2212 2577 2218
rect 2590 2202 2593 2268
rect 2638 2262 2641 2268
rect 2678 2252 2681 2258
rect 2578 2158 2582 2161
rect 2534 2102 2537 2128
rect 2542 2092 2545 2118
rect 2262 2062 2265 2088
rect 2294 2082 2297 2088
rect 2302 2072 2305 2078
rect 2318 2072 2321 2078
rect 2326 2072 2329 2078
rect 2366 2072 2369 2088
rect 2030 1992 2033 1998
rect 2018 1968 2022 1971
rect 2038 1962 2041 1978
rect 1958 1912 1961 1948
rect 2030 1942 2033 1948
rect 2010 1938 2014 1941
rect 1974 1892 1977 1918
rect 1990 1902 1993 1935
rect 1998 1872 2001 1898
rect 1942 1862 1945 1868
rect 1950 1862 1953 1868
rect 2014 1862 2017 1898
rect 2046 1872 2049 1998
rect 2054 1972 2057 1978
rect 2258 1968 2262 1971
rect 2134 1962 2137 1968
rect 2106 1958 2110 1961
rect 2062 1952 2065 1958
rect 2070 1942 2073 1958
rect 2094 1942 2097 1958
rect 2142 1952 2145 1958
rect 2166 1952 2169 1968
rect 2118 1942 2121 1948
rect 2150 1942 2153 1948
rect 2178 1938 2190 1941
rect 2062 1932 2065 1938
rect 2078 1932 2081 1938
rect 2126 1922 2129 1938
rect 2086 1902 2089 1918
rect 2102 1892 2105 1918
rect 2038 1868 2046 1871
rect 2066 1868 2070 1871
rect 1926 1852 1929 1858
rect 2038 1852 2041 1868
rect 2050 1858 2054 1861
rect 2086 1852 2089 1888
rect 2106 1878 2110 1881
rect 2094 1872 2097 1878
rect 2102 1868 2110 1871
rect 2102 1861 2105 1868
rect 2098 1858 2105 1861
rect 2114 1858 2118 1861
rect 2134 1852 2137 1928
rect 2158 1922 2161 1938
rect 2198 1932 2201 1938
rect 2178 1928 2182 1931
rect 2202 1928 2206 1931
rect 2190 1912 2193 1928
rect 2214 1922 2217 1948
rect 2222 1942 2225 1948
rect 2230 1942 2233 1968
rect 2270 1962 2273 1978
rect 2302 1972 2305 2068
rect 2318 2052 2321 2068
rect 2374 2062 2377 2078
rect 2334 2052 2337 2058
rect 2390 2052 2393 2068
rect 2422 2062 2425 2078
rect 2454 2062 2457 2078
rect 2478 2062 2481 2078
rect 2494 2062 2497 2068
rect 2502 2062 2505 2078
rect 2542 2062 2545 2068
rect 2558 2062 2561 2148
rect 2574 2082 2577 2118
rect 2582 2072 2585 2158
rect 2614 2152 2617 2158
rect 2694 2152 2697 2158
rect 2646 2142 2649 2148
rect 2590 2122 2593 2138
rect 2598 2102 2601 2138
rect 2566 2062 2569 2068
rect 2446 2052 2449 2058
rect 2330 2048 2334 2051
rect 2430 2042 2433 2048
rect 2462 2042 2465 2048
rect 2486 2042 2489 2058
rect 2514 2038 2518 2041
rect 2526 2032 2529 2058
rect 2574 2052 2577 2068
rect 2538 2048 2542 2051
rect 2422 2022 2425 2028
rect 2598 2022 2601 2048
rect 2606 2031 2609 2058
rect 2614 2042 2617 2048
rect 2606 2028 2617 2031
rect 2614 2022 2617 2028
rect 2310 1972 2313 2018
rect 2278 1962 2281 1968
rect 2310 1962 2313 1968
rect 2230 1931 2233 1938
rect 2222 1928 2233 1931
rect 2238 1932 2241 1938
rect 2250 1928 2254 1931
rect 2166 1882 2169 1908
rect 2186 1888 2190 1891
rect 2198 1882 2201 1898
rect 2222 1892 2225 1928
rect 2270 1902 2273 1948
rect 2278 1932 2281 1958
rect 2294 1942 2297 1948
rect 2334 1942 2337 2018
rect 2350 1952 2353 2018
rect 2374 1972 2377 2018
rect 2392 2003 2394 2007
rect 2398 2003 2401 2007
rect 2405 2003 2408 2007
rect 2286 1921 2289 1938
rect 2302 1932 2305 1938
rect 2278 1918 2289 1921
rect 2318 1922 2321 1928
rect 2278 1902 2281 1918
rect 2238 1892 2241 1898
rect 2278 1892 2281 1898
rect 2298 1888 2302 1891
rect 2150 1872 2153 1878
rect 2170 1858 2174 1861
rect 2002 1848 2006 1851
rect 1810 1788 1814 1791
rect 1838 1742 1841 1788
rect 1874 1748 1878 1751
rect 1854 1732 1857 1748
rect 1926 1742 1929 1838
rect 1934 1792 1937 1818
rect 1966 1802 1969 1818
rect 1950 1752 1953 1798
rect 1998 1792 2001 1838
rect 2022 1812 2025 1838
rect 2014 1792 2017 1808
rect 1990 1762 1993 1768
rect 1974 1752 1977 1758
rect 1986 1748 1990 1751
rect 1946 1738 1953 1741
rect 1842 1728 1846 1731
rect 1894 1722 1897 1732
rect 1806 1692 1809 1708
rect 1872 1703 1874 1707
rect 1878 1703 1881 1707
rect 1885 1703 1888 1707
rect 1842 1688 1846 1691
rect 1898 1688 1902 1691
rect 1814 1682 1817 1688
rect 1898 1678 1902 1681
rect 1934 1672 1937 1718
rect 1942 1672 1945 1678
rect 1794 1668 1798 1671
rect 1730 1658 1734 1661
rect 1718 1652 1721 1658
rect 1730 1648 1734 1651
rect 1742 1642 1745 1668
rect 1794 1658 1798 1661
rect 1718 1612 1721 1618
rect 1514 1568 1518 1571
rect 1646 1552 1649 1558
rect 1686 1552 1689 1558
rect 1506 1548 1510 1551
rect 1494 1542 1497 1548
rect 1618 1548 1622 1551
rect 1582 1542 1585 1547
rect 1682 1538 1686 1541
rect 1378 1518 1382 1521
rect 1446 1492 1449 1528
rect 1478 1522 1481 1528
rect 1510 1522 1513 1528
rect 1334 1472 1337 1478
rect 1342 1472 1345 1478
rect 1462 1472 1465 1498
rect 1474 1468 1478 1471
rect 1326 1352 1329 1388
rect 1334 1382 1337 1458
rect 1358 1452 1361 1458
rect 1390 1452 1393 1468
rect 1368 1403 1370 1407
rect 1374 1403 1377 1407
rect 1381 1403 1384 1407
rect 1382 1362 1385 1368
rect 1374 1282 1377 1298
rect 1346 1278 1350 1281
rect 1290 1268 1294 1271
rect 1330 1268 1334 1271
rect 1346 1268 1350 1271
rect 1226 1258 1230 1261
rect 1250 1258 1254 1261
rect 1214 1248 1222 1251
rect 1106 1228 1110 1231
rect 1170 1228 1174 1231
rect 1054 1188 1065 1191
rect 1030 1151 1033 1158
rect 958 1142 961 1148
rect 1018 1138 1022 1141
rect 874 1118 878 1121
rect 910 1121 913 1138
rect 1062 1132 1065 1188
rect 1078 1142 1081 1228
rect 1286 1222 1289 1268
rect 1310 1262 1313 1268
rect 1326 1262 1329 1268
rect 1390 1262 1393 1338
rect 1398 1322 1401 1468
rect 1470 1372 1473 1468
rect 1486 1461 1489 1478
rect 1482 1458 1489 1461
rect 1494 1452 1497 1488
rect 1518 1482 1521 1488
rect 1526 1482 1529 1488
rect 1510 1472 1513 1478
rect 1582 1472 1585 1528
rect 1622 1492 1625 1528
rect 1514 1468 1518 1471
rect 1502 1462 1505 1468
rect 1478 1392 1481 1418
rect 1438 1322 1441 1348
rect 1462 1342 1465 1348
rect 1478 1332 1481 1338
rect 1422 1292 1425 1308
rect 1406 1272 1409 1278
rect 1478 1272 1481 1328
rect 1466 1268 1470 1271
rect 1510 1262 1513 1458
rect 1542 1352 1545 1468
rect 1566 1392 1569 1458
rect 1582 1352 1585 1468
rect 1630 1432 1633 1538
rect 1694 1481 1697 1578
rect 1702 1532 1705 1548
rect 1718 1492 1721 1508
rect 1714 1488 1718 1491
rect 1690 1478 1697 1481
rect 1714 1478 1718 1481
rect 1726 1472 1729 1638
rect 1782 1592 1785 1628
rect 1814 1592 1817 1668
rect 1822 1662 1825 1668
rect 1894 1652 1897 1668
rect 1910 1662 1913 1668
rect 1930 1658 1934 1661
rect 1882 1648 1886 1651
rect 1854 1592 1857 1608
rect 1878 1592 1881 1638
rect 1770 1558 1774 1561
rect 1738 1548 1750 1551
rect 1754 1548 1758 1551
rect 1746 1538 1750 1541
rect 1766 1532 1769 1538
rect 1754 1528 1758 1531
rect 1790 1501 1793 1538
rect 1798 1512 1801 1558
rect 1790 1498 1801 1501
rect 1786 1478 1790 1481
rect 1758 1472 1761 1478
rect 1730 1468 1734 1471
rect 1742 1462 1745 1468
rect 1750 1462 1753 1468
rect 1706 1458 1710 1461
rect 1646 1452 1649 1458
rect 1766 1442 1769 1448
rect 1646 1392 1649 1438
rect 1774 1432 1777 1468
rect 1790 1442 1793 1448
rect 1542 1342 1545 1348
rect 1614 1342 1617 1347
rect 1630 1342 1633 1348
rect 1550 1282 1553 1318
rect 1638 1292 1641 1318
rect 1654 1292 1657 1428
rect 1678 1342 1681 1348
rect 1686 1282 1689 1418
rect 1710 1351 1713 1408
rect 1798 1402 1801 1498
rect 1806 1492 1809 1528
rect 1814 1492 1817 1548
rect 1822 1542 1825 1548
rect 1830 1492 1833 1548
rect 1818 1478 1822 1481
rect 1838 1472 1841 1538
rect 1854 1532 1857 1568
rect 1878 1532 1881 1548
rect 1886 1532 1889 1538
rect 1822 1462 1825 1468
rect 1838 1422 1841 1448
rect 1758 1392 1761 1398
rect 1854 1392 1857 1528
rect 1872 1503 1874 1507
rect 1878 1503 1881 1507
rect 1885 1503 1888 1507
rect 1894 1492 1897 1538
rect 1910 1532 1913 1658
rect 1918 1632 1921 1658
rect 1926 1552 1929 1558
rect 1934 1552 1937 1568
rect 1950 1562 1953 1738
rect 1982 1692 1985 1728
rect 2006 1692 2009 1758
rect 2014 1752 2017 1778
rect 2030 1772 2033 1818
rect 1958 1682 1961 1688
rect 1974 1682 1977 1688
rect 1966 1672 1969 1678
rect 1966 1652 1969 1668
rect 1990 1652 1993 1668
rect 2002 1658 2006 1661
rect 1974 1592 1977 1628
rect 2006 1592 2009 1648
rect 2014 1592 2017 1748
rect 2038 1732 2041 1788
rect 2054 1771 2057 1818
rect 2046 1768 2057 1771
rect 2046 1742 2049 1768
rect 2094 1742 2097 1808
rect 2102 1792 2105 1848
rect 2122 1818 2126 1821
rect 2142 1802 2145 1858
rect 2134 1792 2137 1798
rect 2038 1692 2041 1728
rect 2046 1692 2049 1708
rect 2022 1662 2025 1668
rect 2030 1612 2033 1668
rect 2078 1582 2081 1718
rect 2110 1702 2113 1768
rect 2118 1742 2121 1748
rect 2106 1688 2110 1691
rect 2086 1672 2089 1678
rect 2134 1672 2137 1748
rect 2142 1732 2145 1778
rect 2150 1752 2153 1758
rect 2158 1742 2161 1768
rect 2166 1762 2169 1818
rect 2182 1762 2185 1818
rect 2190 1772 2193 1878
rect 2246 1872 2249 1888
rect 2326 1872 2329 1918
rect 2342 1882 2345 1908
rect 2350 1902 2353 1938
rect 2358 1932 2361 1968
rect 2370 1938 2374 1941
rect 2370 1918 2374 1921
rect 2422 1872 2425 1998
rect 2454 1972 2457 2018
rect 2430 1932 2433 1958
rect 2446 1942 2449 1958
rect 2454 1952 2457 1968
rect 2462 1952 2465 1978
rect 2470 1962 2473 2018
rect 2510 2002 2513 2018
rect 2606 2002 2609 2018
rect 2622 1982 2625 2108
rect 2670 2092 2673 2148
rect 2678 2112 2681 2138
rect 2630 2052 2633 2078
rect 2646 2042 2649 2068
rect 2686 2062 2689 2118
rect 2658 2058 2662 2061
rect 2674 2058 2678 2061
rect 2666 2048 2670 2051
rect 2694 2042 2697 2138
rect 2702 2102 2705 2318
rect 2758 2302 2761 2468
rect 2782 2412 2785 2468
rect 2766 2352 2769 2378
rect 2750 2222 2753 2228
rect 2762 2158 2766 2161
rect 2718 2142 2721 2148
rect 2782 2142 2785 2398
rect 2790 2272 2793 2478
rect 2798 2402 2801 2538
rect 2806 2512 2809 2658
rect 2838 2632 2841 2668
rect 2862 2662 2865 2748
rect 2886 2672 2889 2758
rect 2894 2752 2897 2768
rect 2918 2762 2921 2768
rect 2894 2672 2897 2748
rect 2904 2703 2906 2707
rect 2910 2703 2913 2707
rect 2917 2703 2920 2707
rect 2926 2692 2929 2768
rect 2902 2672 2905 2678
rect 2934 2662 2937 2758
rect 2946 2748 2950 2751
rect 2970 2748 2974 2751
rect 2970 2728 2974 2731
rect 2982 2722 2985 2758
rect 3006 2751 3009 2808
rect 3022 2792 3025 2798
rect 3150 2792 3153 2808
rect 3166 2802 3169 2858
rect 3182 2842 3185 2908
rect 3246 2902 3249 2918
rect 3262 2892 3265 2938
rect 3302 2932 3305 2938
rect 3318 2932 3321 2938
rect 3278 2922 3281 2928
rect 3366 2922 3369 2948
rect 3382 2942 3385 2958
rect 3390 2952 3393 3028
rect 3398 3022 3401 3028
rect 3416 3003 3418 3007
rect 3422 3003 3425 3007
rect 3429 3003 3432 3007
rect 3406 2942 3409 2958
rect 3414 2931 3417 2958
rect 3422 2952 3425 2968
rect 3470 2962 3473 3128
rect 3582 3122 3585 3148
rect 3594 3128 3598 3131
rect 3630 3122 3633 3158
rect 3658 3148 3662 3151
rect 3694 3151 3697 3158
rect 3894 3152 3897 3268
rect 3910 3263 3913 3318
rect 3918 3312 3921 3328
rect 3926 3322 3929 3348
rect 3928 3303 3930 3307
rect 3934 3303 3937 3307
rect 3941 3303 3944 3307
rect 3950 3262 3953 3388
rect 3962 3368 3966 3371
rect 3974 3292 3977 3328
rect 3982 3252 3985 3418
rect 4014 3382 4017 3418
rect 4054 3362 4057 3468
rect 4118 3462 4121 3508
rect 4126 3472 4129 3528
rect 4142 3482 4145 3488
rect 4086 3372 4089 3458
rect 4094 3422 4097 3458
rect 4078 3352 4081 3368
rect 4086 3352 4089 3358
rect 3998 3292 4001 3308
rect 4022 3292 4025 3348
rect 4030 3312 4033 3348
rect 4038 3322 4041 3328
rect 4038 3262 4041 3308
rect 4050 3288 4054 3291
rect 4078 3272 4081 3328
rect 4094 3312 4097 3418
rect 4118 3392 4121 3458
rect 4114 3368 4118 3371
rect 4110 3352 4113 3358
rect 4102 3332 4105 3348
rect 4126 3292 4129 3468
rect 4150 3442 4153 3538
rect 4302 3532 4305 3538
rect 4334 3532 4337 3568
rect 4402 3558 4406 3561
rect 4342 3542 4345 3558
rect 4158 3441 4161 3518
rect 4190 3492 4193 3518
rect 4174 3482 4177 3488
rect 4230 3481 4233 3528
rect 4230 3478 4241 3481
rect 4186 3468 4190 3471
rect 4210 3468 4214 3471
rect 4230 3462 4233 3468
rect 4238 3462 4241 3478
rect 4178 3458 4182 3461
rect 4194 3458 4198 3461
rect 4206 3452 4209 3458
rect 4186 3448 4190 3451
rect 4158 3438 4166 3441
rect 4174 3352 4177 3378
rect 4214 3342 4217 3438
rect 4222 3392 4225 3458
rect 4238 3402 4241 3458
rect 4246 3442 4249 3468
rect 4270 3462 4273 3468
rect 4278 3462 4281 3488
rect 4294 3462 4297 3478
rect 4326 3472 4329 3518
rect 4342 3472 4345 3538
rect 4350 3472 4353 3548
rect 4358 3542 4361 3558
rect 4378 3548 4382 3551
rect 4398 3542 4401 3548
rect 4414 3542 4417 3628
rect 4440 3603 4442 3607
rect 4446 3603 4449 3607
rect 4453 3603 4456 3607
rect 4426 3538 4430 3541
rect 4358 3482 4361 3488
rect 4374 3472 4377 3538
rect 4306 3468 4310 3471
rect 4354 3468 4361 3471
rect 4298 3458 4302 3461
rect 4326 3452 4329 3458
rect 4334 3452 4337 3458
rect 4290 3448 4294 3451
rect 4254 3442 4257 3448
rect 4270 3442 4273 3448
rect 4342 3442 4345 3448
rect 4358 3441 4361 3468
rect 4382 3462 4385 3518
rect 4406 3482 4409 3488
rect 4414 3472 4417 3538
rect 4422 3482 4425 3488
rect 4390 3462 4393 3468
rect 4406 3462 4409 3468
rect 4370 3448 4374 3451
rect 4358 3438 4369 3441
rect 4238 3362 4241 3368
rect 4278 3342 4281 3347
rect 4350 3342 4353 3348
rect 4366 3342 4369 3438
rect 4390 3362 4393 3428
rect 4390 3352 4393 3358
rect 4398 3342 4401 3438
rect 4110 3252 4113 3259
rect 4198 3262 4201 3338
rect 4214 3282 4217 3338
rect 4246 3322 4249 3328
rect 4230 3292 4233 3298
rect 4262 3282 4265 3338
rect 4358 3332 4361 3338
rect 4326 3292 4329 3328
rect 4390 3312 4393 3318
rect 4414 3302 4417 3468
rect 4438 3462 4441 3588
rect 4446 3542 4449 3578
rect 4462 3572 4465 3638
rect 4462 3542 4465 3568
rect 4446 3532 4449 3538
rect 4470 3522 4473 3558
rect 4494 3552 4497 3658
rect 4502 3642 4505 3658
rect 4510 3561 4513 3658
rect 4526 3642 4529 3658
rect 4574 3652 4577 3658
rect 4598 3642 4601 3648
rect 4678 3632 4681 3668
rect 4718 3652 4721 3658
rect 4518 3582 4521 3618
rect 4502 3558 4513 3561
rect 4486 3542 4489 3548
rect 4502 3542 4505 3558
rect 4510 3542 4513 3548
rect 4518 3542 4521 3568
rect 4526 3552 4529 3558
rect 4558 3552 4561 3578
rect 4542 3542 4545 3548
rect 4582 3542 4585 3558
rect 4590 3552 4593 3568
rect 4666 3558 4670 3561
rect 4614 3552 4617 3558
rect 4666 3548 4670 3551
rect 4630 3542 4633 3548
rect 4638 3542 4641 3548
rect 4646 3542 4649 3548
rect 4562 3538 4566 3541
rect 4610 3538 4614 3541
rect 4470 3492 4473 3518
rect 4494 3502 4497 3518
rect 4474 3478 4478 3481
rect 4486 3472 4489 3488
rect 4494 3482 4497 3488
rect 4462 3462 4465 3468
rect 4494 3462 4497 3468
rect 4502 3461 4505 3538
rect 4510 3471 4513 3538
rect 4566 3528 4569 3538
rect 4526 3492 4529 3518
rect 4522 3478 4526 3481
rect 4510 3468 4518 3471
rect 4542 3462 4545 3488
rect 4502 3458 4510 3461
rect 4478 3442 4481 3448
rect 4458 3438 4462 3441
rect 4440 3403 4442 3407
rect 4446 3403 4449 3407
rect 4453 3403 4456 3407
rect 4502 3392 4505 3458
rect 4550 3452 4553 3498
rect 4574 3491 4577 3518
rect 4566 3488 4577 3491
rect 4566 3472 4569 3488
rect 4574 3472 4577 3478
rect 4610 3468 4614 3471
rect 4630 3462 4633 3538
rect 4670 3532 4673 3538
rect 4678 3532 4681 3628
rect 4694 3562 4697 3578
rect 4718 3562 4721 3648
rect 4734 3622 4737 3678
rect 4762 3658 4766 3661
rect 4734 3592 4737 3618
rect 4766 3572 4769 3638
rect 4782 3622 4785 3658
rect 4814 3632 4817 3658
rect 4766 3562 4769 3568
rect 4706 3558 4710 3561
rect 4706 3538 4710 3541
rect 4666 3528 4670 3531
rect 4646 3472 4649 3478
rect 4442 3358 4446 3361
rect 4542 3352 4545 3418
rect 4462 3342 4465 3348
rect 4434 3328 4438 3331
rect 4470 3302 4473 3338
rect 4478 3302 4481 3348
rect 4362 3288 4366 3291
rect 4326 3272 4329 3288
rect 4486 3282 4489 3338
rect 4494 3292 4497 3298
rect 4502 3282 4505 3308
rect 4382 3272 4385 3278
rect 4406 3275 4410 3278
rect 4486 3272 4489 3278
rect 4510 3272 4513 3278
rect 4534 3272 4537 3308
rect 4542 3292 4545 3338
rect 4558 3322 4561 3348
rect 4566 3291 4569 3438
rect 4590 3412 4593 3458
rect 4626 3448 4630 3451
rect 4598 3361 4601 3418
rect 4654 3402 4657 3468
rect 4598 3358 4609 3361
rect 4598 3342 4601 3348
rect 4582 3312 4585 3338
rect 4606 3322 4609 3358
rect 4614 3342 4617 3358
rect 4662 3351 4665 3518
rect 4710 3492 4713 3528
rect 4718 3512 4721 3548
rect 4718 3442 4721 3508
rect 4734 3492 4737 3558
rect 4782 3552 4785 3618
rect 4830 3592 4833 3668
rect 4846 3663 4849 3678
rect 4846 3552 4849 3558
rect 4862 3552 4865 3728
rect 4878 3552 4881 3728
rect 4952 3703 4954 3707
rect 4958 3703 4961 3707
rect 4965 3703 4968 3707
rect 5182 3692 5185 3728
rect 5154 3688 5158 3691
rect 4894 3682 4897 3688
rect 4886 3622 4889 3678
rect 4998 3672 5001 3678
rect 4894 3662 4897 3668
rect 4982 3662 4985 3668
rect 4902 3652 4905 3658
rect 4990 3652 4993 3658
rect 4990 3552 4993 3648
rect 5006 3622 5009 3678
rect 5038 3672 5041 3678
rect 5062 3662 5065 3688
rect 5190 3679 5198 3681
rect 5190 3678 5201 3679
rect 4882 3548 4886 3551
rect 4750 3522 4753 3548
rect 4774 3532 4777 3548
rect 4806 3542 4809 3548
rect 4766 3492 4769 3498
rect 4774 3482 4777 3488
rect 4798 3472 4801 3488
rect 4758 3462 4761 3468
rect 4822 3462 4825 3538
rect 4838 3532 4841 3548
rect 4862 3542 4865 3548
rect 4918 3542 4921 3548
rect 4854 3522 4857 3538
rect 4894 3532 4897 3538
rect 4918 3532 4921 3538
rect 4854 3502 4857 3518
rect 4830 3472 4833 3498
rect 4878 3482 4881 3518
rect 4898 3488 4902 3491
rect 4918 3491 4921 3518
rect 4910 3488 4921 3491
rect 4750 3422 4753 3458
rect 4778 3448 4782 3451
rect 4674 3358 4678 3361
rect 4658 3348 4665 3351
rect 4694 3352 4697 3378
rect 4710 3342 4713 3418
rect 4626 3338 4633 3341
rect 4642 3338 4646 3341
rect 4630 3332 4633 3338
rect 4618 3328 4622 3331
rect 4566 3288 4577 3291
rect 4550 3282 4553 3288
rect 4574 3282 4577 3288
rect 4562 3278 4566 3281
rect 4606 3272 4609 3308
rect 4330 3268 4334 3271
rect 4038 3192 4041 3248
rect 4150 3192 4153 3258
rect 4166 3252 4169 3259
rect 4198 3212 4201 3258
rect 4246 3212 4249 3268
rect 4390 3262 4393 3268
rect 4466 3258 4470 3261
rect 4554 3258 4558 3261
rect 4270 3252 4273 3258
rect 4462 3242 4465 3248
rect 4418 3238 4422 3241
rect 4214 3192 4217 3208
rect 3930 3188 3934 3191
rect 4158 3152 4161 3168
rect 3770 3148 3774 3151
rect 3946 3148 3950 3151
rect 3726 3142 3729 3148
rect 3870 3142 3873 3148
rect 3894 3142 3897 3148
rect 4014 3142 4017 3148
rect 4010 3138 4014 3141
rect 3646 3132 3649 3138
rect 3830 3132 3833 3138
rect 3990 3132 3993 3138
rect 3502 3072 3505 3108
rect 3928 3103 3930 3107
rect 3934 3103 3937 3107
rect 3941 3103 3944 3107
rect 3878 3092 3881 3098
rect 3990 3092 3993 3128
rect 3818 3088 3822 3091
rect 4022 3091 4025 3138
rect 4018 3088 4025 3091
rect 4070 3092 4073 3138
rect 4078 3131 4081 3148
rect 4102 3131 4105 3148
rect 4158 3142 4161 3148
rect 4078 3128 4086 3131
rect 4102 3128 4110 3131
rect 3538 3078 3542 3081
rect 3586 3078 3590 3081
rect 3642 3078 3646 3081
rect 3518 3072 3521 3078
rect 3534 3062 3537 3068
rect 3490 3058 3494 3061
rect 3494 3042 3497 3048
rect 3502 3031 3505 3058
rect 3550 3052 3553 3078
rect 3558 3062 3561 3068
rect 3494 3028 3505 3031
rect 3494 2982 3497 3028
rect 3506 2978 3510 2981
rect 3406 2928 3417 2931
rect 3278 2892 3281 2908
rect 3274 2878 3278 2881
rect 3206 2872 3209 2878
rect 3242 2868 3249 2871
rect 3194 2858 3198 2861
rect 3194 2848 3198 2851
rect 3006 2748 3014 2751
rect 2990 2742 2993 2748
rect 2878 2652 2881 2658
rect 2910 2592 2913 2628
rect 2942 2622 2945 2678
rect 2958 2632 2961 2668
rect 2974 2652 2977 2659
rect 2982 2622 2985 2718
rect 3006 2682 3009 2748
rect 3030 2742 3033 2768
rect 3038 2742 3041 2748
rect 3118 2742 3121 2788
rect 3194 2778 3198 2781
rect 3054 2732 3057 2738
rect 3034 2728 3038 2731
rect 3062 2722 3065 2728
rect 3070 2721 3073 2738
rect 3126 2722 3129 2748
rect 3134 2742 3137 2748
rect 3070 2718 3078 2721
rect 3102 2702 3105 2718
rect 3038 2692 3041 2698
rect 3134 2692 3137 2738
rect 3150 2732 3153 2778
rect 3174 2772 3177 2778
rect 3158 2722 3161 2758
rect 3166 2742 3169 2748
rect 3206 2742 3209 2848
rect 3222 2832 3225 2858
rect 3230 2812 3233 2868
rect 3238 2862 3241 2868
rect 3222 2792 3225 2798
rect 3246 2752 3249 2868
rect 3254 2862 3257 2868
rect 3294 2862 3297 2878
rect 3302 2872 3305 2898
rect 3406 2892 3409 2928
rect 3430 2922 3433 2958
rect 3446 2932 3449 2938
rect 3454 2922 3457 2948
rect 3470 2932 3473 2938
rect 3486 2932 3489 2948
rect 3494 2942 3497 2978
rect 3518 2972 3521 2978
rect 3526 2972 3529 2978
rect 3534 2962 3537 2968
rect 3522 2948 3526 2951
rect 3534 2941 3537 2958
rect 3558 2952 3561 3018
rect 3546 2948 3550 2951
rect 3566 2942 3569 3048
rect 3598 3042 3601 3068
rect 3606 3052 3609 3058
rect 3614 3052 3617 3078
rect 3782 3072 3785 3078
rect 3950 3072 3953 3078
rect 3626 3068 3630 3071
rect 3690 3068 3694 3071
rect 3714 3068 3721 3071
rect 3666 3058 3670 3061
rect 3690 3058 3694 3061
rect 3622 3052 3625 3058
rect 3706 3048 3710 3051
rect 3598 3032 3601 3038
rect 3582 2962 3585 2968
rect 3574 2952 3577 2958
rect 3606 2952 3609 3018
rect 3614 2962 3617 3048
rect 3670 3042 3673 3048
rect 3678 2992 3681 3048
rect 3718 3042 3721 3068
rect 4014 3070 4017 3088
rect 3630 2962 3633 2988
rect 3702 2962 3705 2968
rect 3630 2952 3633 2958
rect 3642 2948 3646 2951
rect 3534 2938 3542 2941
rect 3562 2938 3566 2941
rect 3562 2918 3566 2921
rect 3254 2842 3257 2848
rect 3270 2832 3273 2848
rect 3270 2792 3273 2828
rect 3294 2792 3297 2858
rect 3310 2782 3313 2878
rect 3326 2862 3329 2888
rect 3422 2872 3425 2908
rect 3438 2902 3441 2918
rect 3462 2912 3465 2918
rect 3494 2892 3497 2918
rect 3466 2888 3470 2891
rect 3570 2888 3574 2891
rect 3442 2878 3446 2881
rect 3370 2868 3374 2871
rect 3590 2871 3593 2938
rect 3598 2912 3601 2948
rect 3670 2942 3673 2958
rect 3686 2952 3689 2958
rect 3682 2948 3686 2951
rect 3718 2951 3721 3018
rect 3726 2992 3729 3068
rect 3754 3058 3758 3061
rect 3790 3032 3793 3068
rect 3838 3062 3841 3068
rect 3846 3052 3849 3068
rect 3838 2992 3841 3038
rect 3870 2992 3873 3048
rect 3894 3042 3897 3068
rect 3902 3062 3905 3068
rect 4006 3062 4009 3068
rect 4030 3062 4033 3068
rect 4038 3062 4041 3078
rect 4086 3062 4089 3108
rect 4126 3072 4129 3138
rect 4134 3132 4137 3140
rect 4142 3072 4145 3128
rect 4166 3082 4169 3088
rect 4182 3082 4185 3148
rect 4234 3138 4238 3141
rect 4222 3092 4225 3138
rect 4254 3132 4257 3138
rect 4230 3092 4233 3118
rect 4262 3112 4265 3158
rect 4286 3152 4289 3158
rect 4270 3142 4273 3148
rect 4334 3142 4337 3208
rect 4350 3151 4353 3158
rect 4318 3132 4321 3138
rect 4094 3062 4097 3068
rect 4166 3062 4169 3068
rect 3922 3058 3926 3061
rect 4066 3058 4070 3061
rect 4154 3058 4158 3061
rect 3974 3052 3977 3058
rect 4054 3052 4057 3058
rect 4086 3052 4089 3058
rect 4042 3048 4046 3051
rect 4114 3048 4118 3051
rect 4074 3038 4078 3041
rect 4106 3038 4110 3041
rect 4154 3038 4158 3041
rect 3734 2962 3737 2978
rect 3718 2948 3729 2951
rect 3738 2948 3742 2951
rect 3610 2938 3614 2941
rect 3658 2938 3662 2941
rect 3630 2932 3633 2938
rect 3638 2922 3641 2928
rect 3654 2922 3657 2928
rect 3694 2922 3697 2948
rect 3714 2938 3718 2941
rect 3622 2882 3625 2908
rect 3638 2872 3641 2898
rect 3654 2892 3657 2918
rect 3710 2882 3713 2918
rect 3726 2892 3729 2948
rect 3750 2942 3753 2978
rect 3766 2972 3769 2978
rect 4094 2971 4097 3018
rect 4110 2992 4113 3018
rect 4158 2992 4161 3028
rect 4182 2992 4185 3078
rect 4238 3072 4241 3108
rect 4270 3092 4273 3118
rect 4398 3092 4401 3228
rect 4440 3203 4442 3207
rect 4446 3203 4449 3207
rect 4453 3203 4456 3207
rect 4470 3192 4473 3238
rect 4418 3178 4422 3181
rect 4550 3142 4553 3168
rect 4438 3092 4441 3138
rect 4462 3112 4465 3132
rect 4462 3092 4465 3108
rect 4494 3102 4497 3138
rect 4510 3082 4513 3118
rect 4362 3078 4366 3081
rect 4298 3068 4302 3071
rect 4190 3032 4193 3068
rect 4246 3032 4249 3068
rect 4334 3062 4337 3068
rect 4342 3062 4345 3078
rect 4438 3072 4441 3078
rect 4510 3072 4513 3078
rect 4490 3068 4494 3071
rect 4366 3062 4369 3068
rect 4406 3062 4409 3068
rect 4526 3062 4529 3068
rect 4534 3062 4537 3088
rect 4542 3072 4545 3138
rect 4550 3092 4553 3138
rect 4574 3092 4577 3258
rect 4606 3192 4609 3268
rect 4630 3262 4633 3318
rect 4654 3282 4657 3338
rect 4674 3328 4678 3331
rect 4670 3301 4673 3318
rect 4670 3298 4681 3301
rect 4666 3288 4670 3291
rect 4678 3272 4681 3298
rect 4686 3282 4689 3318
rect 4698 3278 4702 3281
rect 4710 3262 4713 3318
rect 4726 3302 4729 3418
rect 4790 3381 4793 3458
rect 4798 3452 4801 3458
rect 4810 3448 4814 3451
rect 4798 3392 4801 3408
rect 4790 3378 4801 3381
rect 4734 3342 4737 3348
rect 4790 3342 4793 3368
rect 4798 3312 4801 3378
rect 4810 3368 4814 3371
rect 4814 3302 4817 3348
rect 4822 3322 4825 3358
rect 4830 3332 4833 3448
rect 4838 3362 4841 3368
rect 4846 3352 4849 3478
rect 4910 3472 4913 3488
rect 4926 3481 4929 3528
rect 4918 3478 4929 3481
rect 4918 3472 4921 3478
rect 4942 3472 4945 3538
rect 4950 3522 4953 3548
rect 5014 3542 5017 3648
rect 5022 3562 5025 3658
rect 5030 3652 5033 3658
rect 5078 3632 5081 3668
rect 5190 3662 5193 3678
rect 5094 3652 5097 3659
rect 5022 3552 5025 3558
rect 5062 3552 5065 3568
rect 4952 3503 4954 3507
rect 4958 3503 4961 3507
rect 4965 3503 4968 3507
rect 4998 3492 5001 3518
rect 5014 3481 5017 3538
rect 5010 3478 5017 3481
rect 5022 3472 5025 3548
rect 4858 3468 4862 3471
rect 4882 3468 4886 3471
rect 4930 3468 4934 3471
rect 4854 3372 4857 3458
rect 4854 3342 4857 3368
rect 4862 3352 4865 3468
rect 4998 3462 5001 3468
rect 5006 3462 5009 3468
rect 4890 3458 4894 3461
rect 4890 3448 4894 3451
rect 4878 3442 4881 3448
rect 4910 3362 4913 3368
rect 4898 3358 4902 3361
rect 4926 3352 4929 3418
rect 4882 3348 4886 3351
rect 4834 3328 4838 3331
rect 4726 3292 4729 3298
rect 4758 3282 4761 3288
rect 4738 3278 4742 3281
rect 4674 3258 4678 3261
rect 4614 3252 4617 3258
rect 4726 3192 4729 3248
rect 4626 3148 4630 3151
rect 4662 3151 4665 3158
rect 4734 3152 4737 3268
rect 4742 3262 4745 3268
rect 4774 3262 4777 3298
rect 4838 3292 4841 3298
rect 4854 3292 4857 3318
rect 4862 3292 4865 3348
rect 4934 3342 4937 3458
rect 5014 3452 5017 3458
rect 5030 3432 5033 3548
rect 5070 3532 5073 3618
rect 5126 3552 5129 3558
rect 5090 3548 5094 3551
rect 5070 3482 5073 3528
rect 5062 3462 5065 3478
rect 5078 3462 5081 3548
rect 5142 3542 5145 3638
rect 5218 3618 5222 3621
rect 5218 3568 5222 3571
rect 5158 3551 5161 3558
rect 4982 3372 4985 3418
rect 5010 3358 5014 3361
rect 4982 3352 4985 3358
rect 4990 3352 4993 3358
rect 5022 3352 5025 3358
rect 4882 3338 4886 3341
rect 4898 3338 4902 3341
rect 4870 3332 4873 3338
rect 4934 3332 4937 3338
rect 4966 3332 4969 3338
rect 5006 3332 5009 3348
rect 5042 3338 5046 3341
rect 5054 3338 5062 3341
rect 5038 3328 5046 3331
rect 4850 3278 4854 3281
rect 4806 3252 4809 3278
rect 4870 3270 4873 3298
rect 4894 3292 4897 3308
rect 4952 3303 4954 3307
rect 4958 3303 4961 3307
rect 4965 3303 4968 3307
rect 4930 3288 4934 3291
rect 4890 3278 4894 3281
rect 4902 3272 4905 3288
rect 5038 3282 5041 3328
rect 5054 3292 5057 3338
rect 5070 3292 5073 3348
rect 5078 3342 5081 3368
rect 5094 3362 5097 3488
rect 5142 3482 5145 3538
rect 5230 3492 5233 3728
rect 5238 3728 5242 3732
rect 5238 3702 5241 3728
rect 5250 3658 5254 3661
rect 5278 3652 5281 3659
rect 5246 3592 5249 3648
rect 5298 3568 5302 3571
rect 5290 3558 5294 3561
rect 5250 3548 5254 3551
rect 5282 3548 5286 3551
rect 5266 3528 5270 3531
rect 5206 3482 5209 3488
rect 5254 3462 5257 3508
rect 5262 3472 5265 3518
rect 5110 3452 5113 3458
rect 5142 3452 5145 3459
rect 5270 3452 5273 3458
rect 5262 3442 5265 3448
rect 5110 3372 5113 3378
rect 5122 3368 5126 3371
rect 5138 3368 5142 3371
rect 5102 3362 5105 3368
rect 5094 3352 5097 3358
rect 5106 3348 5110 3351
rect 5182 3351 5185 3358
rect 5134 3342 5137 3348
rect 5190 3342 5193 3438
rect 5278 3432 5281 3438
rect 5242 3388 5246 3391
rect 5270 3372 5273 3418
rect 5286 3362 5289 3518
rect 5274 3358 5278 3361
rect 5090 3338 5094 3341
rect 5250 3338 5254 3341
rect 5102 3292 5105 3338
rect 5150 3322 5153 3328
rect 5190 3292 5193 3328
rect 4954 3278 4958 3281
rect 4994 3278 4998 3281
rect 5146 3278 5150 3281
rect 4918 3272 4921 3278
rect 4942 3272 4945 3278
rect 5022 3272 5025 3278
rect 5062 3272 5065 3278
rect 4830 3262 4833 3268
rect 4890 3268 4894 3271
rect 4910 3262 4913 3268
rect 4934 3252 4937 3268
rect 4958 3262 4961 3268
rect 4982 3252 4985 3268
rect 4998 3262 5001 3268
rect 5046 3262 5049 3268
rect 5046 3252 5049 3258
rect 4758 3162 4761 3218
rect 4790 3152 4793 3218
rect 4858 3188 4862 3191
rect 4842 3168 4846 3171
rect 4862 3152 4865 3158
rect 4870 3152 4873 3158
rect 4774 3142 4777 3148
rect 4798 3141 4801 3148
rect 4790 3138 4801 3141
rect 4622 3122 4625 3128
rect 4590 3072 4593 3078
rect 4606 3072 4609 3118
rect 4394 3058 4398 3061
rect 4278 2992 4281 3038
rect 4318 3032 4321 3058
rect 4302 3011 4305 3018
rect 4294 3008 4305 3011
rect 4086 2968 4097 2971
rect 3798 2962 3801 2968
rect 4086 2962 4089 2968
rect 3806 2952 3809 2958
rect 3910 2952 3913 2958
rect 4006 2952 4009 2958
rect 4086 2952 4089 2958
rect 3834 2948 3838 2951
rect 3762 2928 3766 2931
rect 3774 2931 3777 2948
rect 3850 2938 3854 2941
rect 3774 2928 3782 2931
rect 3822 2922 3825 2938
rect 3902 2932 3905 2938
rect 3846 2922 3849 2928
rect 3742 2892 3745 2898
rect 3798 2882 3801 2918
rect 3658 2878 3662 2881
rect 3590 2868 3598 2871
rect 3450 2858 3454 2861
rect 3474 2858 3478 2861
rect 3334 2812 3337 2858
rect 3494 2852 3497 2868
rect 3510 2862 3513 2868
rect 3494 2812 3497 2848
rect 3534 2822 3537 2858
rect 3542 2852 3545 2868
rect 3666 2858 3670 2861
rect 3682 2858 3686 2861
rect 3638 2852 3641 2858
rect 3650 2848 3654 2851
rect 3674 2848 3678 2851
rect 3614 2842 3617 2848
rect 3694 2842 3697 2868
rect 3686 2832 3689 2838
rect 3416 2803 3418 2807
rect 3422 2803 3425 2807
rect 3429 2803 3432 2807
rect 3470 2792 3473 2808
rect 3694 2792 3697 2828
rect 3710 2792 3713 2868
rect 3782 2862 3785 2878
rect 3802 2868 3806 2871
rect 3814 2862 3817 2868
rect 3830 2862 3833 2908
rect 3928 2903 3930 2907
rect 3934 2903 3937 2907
rect 3941 2903 3944 2907
rect 3846 2882 3849 2888
rect 3898 2868 3902 2871
rect 3734 2792 3737 2858
rect 3862 2852 3865 2868
rect 3870 2862 3873 2868
rect 3766 2792 3769 2838
rect 3878 2832 3881 2858
rect 3310 2772 3313 2778
rect 3258 2768 3262 2771
rect 3294 2758 3302 2761
rect 3274 2748 3278 2751
rect 3178 2738 3182 2741
rect 3206 2732 3209 2738
rect 3194 2728 3198 2731
rect 3046 2688 3054 2691
rect 3046 2672 3049 2688
rect 3094 2672 3097 2678
rect 3118 2662 3121 2678
rect 3062 2622 3065 2628
rect 3030 2592 3033 2598
rect 3054 2592 3057 2618
rect 2850 2548 2854 2551
rect 2834 2538 2838 2541
rect 2858 2538 2862 2541
rect 2814 2522 2817 2528
rect 2822 2392 2825 2448
rect 2830 2442 2833 2498
rect 2886 2492 2889 2548
rect 2966 2542 2969 2547
rect 3038 2542 3041 2558
rect 3062 2552 3065 2618
rect 3126 2602 3129 2668
rect 3142 2652 3145 2668
rect 3110 2562 3113 2598
rect 3122 2568 3126 2571
rect 3074 2558 3078 2561
rect 3106 2558 3110 2561
rect 3142 2561 3145 2648
rect 3150 2632 3153 2658
rect 3158 2592 3161 2708
rect 3166 2682 3169 2698
rect 3174 2692 3177 2728
rect 3150 2572 3153 2578
rect 3138 2558 3145 2561
rect 3166 2562 3169 2658
rect 3174 2652 3177 2668
rect 3190 2662 3193 2698
rect 3198 2672 3201 2708
rect 3230 2682 3233 2698
rect 3238 2692 3241 2738
rect 3246 2712 3249 2748
rect 3286 2742 3289 2758
rect 3294 2752 3297 2758
rect 3454 2752 3457 2788
rect 3774 2772 3777 2778
rect 3762 2768 3766 2771
rect 3602 2758 3606 2761
rect 3634 2758 3638 2761
rect 3666 2758 3670 2761
rect 3410 2748 3414 2751
rect 3286 2732 3289 2738
rect 3294 2692 3297 2748
rect 3310 2702 3313 2718
rect 3326 2712 3329 2748
rect 3342 2742 3345 2748
rect 3334 2702 3337 2738
rect 3390 2721 3393 2738
rect 3386 2718 3393 2721
rect 3374 2702 3377 2718
rect 3462 2712 3465 2748
rect 3486 2742 3489 2758
rect 3602 2748 3606 2751
rect 3634 2748 3641 2751
rect 3542 2742 3545 2748
rect 3478 2712 3481 2728
rect 3514 2718 3518 2721
rect 3534 2721 3537 2738
rect 3530 2718 3537 2721
rect 3570 2718 3574 2721
rect 3590 2721 3593 2738
rect 3586 2718 3593 2721
rect 3622 2721 3625 2738
rect 3618 2718 3625 2721
rect 3210 2668 3214 2671
rect 3226 2668 3230 2671
rect 3242 2668 3246 2671
rect 3214 2652 3217 2668
rect 3254 2662 3257 2668
rect 3262 2652 3265 2678
rect 3334 2672 3337 2698
rect 3350 2682 3353 2698
rect 3582 2692 3585 2708
rect 3450 2688 3454 2691
rect 3466 2688 3470 2691
rect 3566 2688 3574 2691
rect 3566 2672 3569 2688
rect 3622 2682 3625 2698
rect 3614 2672 3617 2678
rect 3630 2672 3633 2728
rect 3638 2722 3641 2748
rect 3294 2662 3297 2668
rect 3314 2658 3318 2661
rect 3278 2652 3281 2658
rect 3174 2642 3177 2648
rect 3222 2632 3225 2648
rect 3294 2632 3297 2648
rect 3302 2642 3305 2648
rect 3262 2592 3265 2618
rect 3090 2548 3094 2551
rect 3114 2548 3118 2551
rect 3154 2548 3158 2551
rect 3198 2551 3201 2558
rect 3326 2552 3329 2648
rect 3338 2638 3342 2641
rect 3382 2612 3385 2659
rect 3506 2658 3510 2661
rect 3522 2658 3526 2661
rect 3414 2652 3417 2658
rect 3416 2603 3418 2607
rect 3422 2603 3425 2607
rect 3429 2603 3432 2607
rect 3114 2538 3118 2541
rect 2846 2472 2849 2478
rect 2894 2472 2897 2538
rect 2904 2503 2906 2507
rect 2910 2503 2913 2507
rect 2917 2503 2920 2507
rect 2950 2492 2953 2538
rect 2974 2472 2977 2478
rect 3022 2472 3025 2478
rect 2854 2442 2857 2468
rect 2810 2368 2814 2371
rect 2798 2362 2801 2368
rect 2830 2362 2833 2438
rect 2870 2402 2873 2448
rect 2894 2412 2897 2468
rect 3038 2462 3041 2538
rect 3062 2521 3065 2538
rect 3070 2532 3073 2538
rect 3058 2518 3065 2521
rect 3086 2521 3089 2538
rect 3086 2518 3094 2521
rect 3054 2492 3057 2498
rect 3150 2492 3153 2518
rect 3070 2462 3073 2468
rect 3086 2463 3089 2478
rect 3198 2472 3201 2528
rect 3246 2492 3249 2498
rect 3294 2492 3297 2547
rect 3374 2532 3377 2538
rect 3326 2488 3334 2491
rect 3266 2479 3273 2481
rect 3262 2478 3273 2479
rect 2990 2442 2993 2459
rect 3166 2462 3169 2468
rect 3270 2462 3273 2478
rect 3326 2472 3329 2488
rect 3334 2472 3337 2488
rect 3278 2462 3281 2468
rect 3182 2452 3185 2459
rect 3338 2458 3342 2461
rect 3310 2452 3313 2458
rect 3350 2452 3353 2478
rect 3358 2462 3361 2518
rect 3366 2462 3369 2468
rect 3346 2448 3350 2451
rect 3390 2442 3393 2448
rect 3378 2438 3382 2441
rect 2950 2382 2953 2418
rect 2990 2382 2993 2388
rect 2906 2368 2910 2371
rect 2966 2362 2969 2368
rect 2874 2358 2878 2361
rect 2822 2342 2825 2348
rect 2794 2258 2798 2261
rect 2810 2148 2814 2151
rect 2726 2122 2729 2128
rect 2814 2122 2817 2138
rect 2822 2132 2825 2198
rect 2830 2152 2833 2358
rect 2886 2352 2889 2358
rect 2870 2348 2878 2351
rect 2850 2338 2854 2341
rect 2846 2292 2849 2298
rect 2854 2272 2857 2288
rect 2862 2261 2865 2338
rect 2870 2332 2873 2348
rect 2918 2332 2921 2348
rect 2926 2342 2929 2348
rect 2942 2342 2945 2348
rect 2950 2332 2953 2358
rect 2978 2340 2982 2343
rect 2998 2342 3001 2348
rect 3014 2342 3017 2378
rect 3042 2358 3046 2361
rect 3054 2352 3057 2378
rect 3138 2358 3142 2361
rect 3030 2342 3033 2348
rect 2870 2292 2873 2328
rect 2878 2282 2881 2318
rect 2904 2303 2906 2307
rect 2910 2303 2913 2307
rect 2917 2303 2920 2307
rect 2966 2302 2969 2338
rect 2886 2282 2889 2288
rect 2922 2278 2926 2281
rect 2970 2278 2974 2281
rect 2898 2268 2902 2271
rect 2966 2262 2969 2268
rect 2982 2262 2985 2268
rect 2862 2258 2873 2261
rect 2870 2252 2873 2258
rect 2954 2258 2958 2261
rect 2986 2258 2990 2261
rect 2902 2222 2905 2258
rect 2966 2242 2969 2258
rect 2862 2192 2865 2198
rect 2870 2181 2873 2198
rect 2862 2178 2873 2181
rect 2854 2162 2857 2178
rect 2850 2158 2854 2161
rect 2862 2152 2865 2178
rect 2870 2162 2873 2168
rect 2850 2148 2857 2151
rect 2806 2118 2814 2121
rect 2706 2058 2710 2061
rect 2682 2038 2686 2041
rect 2698 2038 2702 2041
rect 2670 2032 2673 2038
rect 2694 2022 2697 2028
rect 2630 2012 2633 2018
rect 2610 1978 2614 1981
rect 2458 1938 2462 1941
rect 2478 1932 2481 1938
rect 2534 1932 2537 1938
rect 2438 1912 2441 1918
rect 2462 1892 2465 1928
rect 2478 1912 2481 1928
rect 2506 1918 2510 1921
rect 2434 1888 2438 1891
rect 2470 1882 2473 1898
rect 2566 1882 2569 1938
rect 2210 1868 2214 1871
rect 2230 1852 2233 1868
rect 2246 1862 2249 1868
rect 2266 1866 2270 1869
rect 2290 1868 2294 1871
rect 2326 1862 2329 1868
rect 2374 1862 2377 1868
rect 2302 1842 2305 1848
rect 2198 1762 2201 1798
rect 2270 1772 2273 1818
rect 2310 1762 2313 1818
rect 2326 1812 2329 1818
rect 2318 1762 2321 1768
rect 2290 1758 2294 1761
rect 2198 1742 2201 1758
rect 2342 1752 2345 1858
rect 2366 1852 2369 1858
rect 2382 1852 2385 1868
rect 2414 1862 2417 1868
rect 2366 1762 2369 1848
rect 2394 1818 2398 1821
rect 2392 1803 2394 1807
rect 2398 1803 2401 1807
rect 2405 1803 2408 1807
rect 2414 1772 2417 1858
rect 2422 1852 2425 1868
rect 2438 1852 2441 1868
rect 2446 1852 2449 1858
rect 2350 1752 2353 1758
rect 2258 1738 2262 1741
rect 2206 1732 2209 1738
rect 2278 1732 2281 1748
rect 2318 1742 2321 1748
rect 2294 1732 2297 1738
rect 2142 1682 2145 1728
rect 2158 1672 2161 1708
rect 2166 1692 2169 1718
rect 2166 1672 2169 1678
rect 2138 1668 2145 1671
rect 1946 1548 1950 1551
rect 1962 1548 1966 1551
rect 1990 1542 1993 1548
rect 2038 1542 2041 1548
rect 1966 1532 1969 1538
rect 2046 1532 2049 1548
rect 2054 1542 2057 1548
rect 2086 1542 2089 1658
rect 2142 1652 2145 1668
rect 2174 1662 2177 1728
rect 2226 1718 2230 1721
rect 2182 1702 2185 1718
rect 2182 1672 2185 1698
rect 2206 1671 2209 1688
rect 2218 1678 2222 1681
rect 2206 1668 2214 1671
rect 2238 1671 2241 1718
rect 2254 1682 2257 1688
rect 2262 1682 2265 1688
rect 2230 1668 2241 1671
rect 2194 1648 2198 1651
rect 2126 1592 2129 1628
rect 2102 1552 2105 1558
rect 2066 1538 2070 1541
rect 1914 1528 1918 1531
rect 1986 1528 1990 1531
rect 2074 1528 2078 1531
rect 1990 1492 1993 1518
rect 2022 1492 2025 1508
rect 2070 1492 2073 1498
rect 1922 1488 1926 1491
rect 1898 1478 1902 1481
rect 2034 1478 2057 1481
rect 1862 1462 1865 1468
rect 1802 1388 1806 1391
rect 1834 1378 1838 1381
rect 1862 1372 1865 1458
rect 1870 1422 1873 1478
rect 1910 1472 1913 1478
rect 1974 1472 1977 1478
rect 1934 1462 1937 1468
rect 1962 1458 1966 1461
rect 1882 1348 1886 1351
rect 1894 1342 1897 1438
rect 1910 1432 1913 1458
rect 1922 1448 1926 1451
rect 1950 1392 1953 1408
rect 1974 1392 1977 1468
rect 1982 1452 1985 1478
rect 2054 1472 2057 1478
rect 2002 1468 2006 1471
rect 2018 1468 2022 1471
rect 2086 1470 2089 1538
rect 2094 1502 2097 1548
rect 2102 1532 2105 1538
rect 2110 1512 2113 1558
rect 2134 1542 2137 1548
rect 2142 1532 2145 1598
rect 2166 1592 2169 1618
rect 2206 1552 2209 1618
rect 2158 1542 2161 1548
rect 2182 1532 2185 1538
rect 2110 1492 2113 1498
rect 2142 1492 2145 1528
rect 2190 1491 2193 1528
rect 2186 1488 2193 1491
rect 2102 1482 2105 1488
rect 2106 1478 2113 1481
rect 2030 1462 2033 1468
rect 2038 1462 2041 1468
rect 2098 1468 2102 1471
rect 2006 1452 2009 1458
rect 1982 1392 1985 1438
rect 2022 1392 2025 1448
rect 2062 1422 2065 1448
rect 1930 1388 1934 1391
rect 1914 1378 1918 1381
rect 1918 1352 1921 1358
rect 1926 1352 1929 1378
rect 1934 1342 1937 1368
rect 1794 1338 1798 1341
rect 1874 1338 1878 1341
rect 1898 1338 1902 1341
rect 1718 1292 1721 1298
rect 1734 1292 1737 1318
rect 1538 1278 1542 1281
rect 1674 1278 1678 1281
rect 1730 1278 1734 1281
rect 1518 1272 1521 1278
rect 1298 1258 1302 1261
rect 1394 1258 1398 1261
rect 1334 1252 1337 1258
rect 1518 1252 1521 1258
rect 1550 1252 1553 1278
rect 1590 1272 1593 1278
rect 1618 1268 1622 1271
rect 1658 1268 1662 1271
rect 1674 1268 1678 1271
rect 1558 1262 1561 1268
rect 1578 1258 1582 1261
rect 1314 1248 1318 1251
rect 1482 1248 1486 1251
rect 1538 1248 1542 1251
rect 1590 1242 1593 1268
rect 1606 1262 1609 1268
rect 1602 1248 1606 1251
rect 1474 1218 1478 1221
rect 1086 1152 1089 1198
rect 1142 1172 1145 1218
rect 1198 1202 1201 1218
rect 1294 1191 1297 1218
rect 1368 1203 1370 1207
rect 1374 1203 1377 1207
rect 1381 1203 1384 1207
rect 1286 1188 1297 1191
rect 1266 1168 1270 1171
rect 910 1118 918 1121
rect 970 1118 974 1121
rect 830 1092 833 1118
rect 856 1103 858 1107
rect 862 1103 865 1107
rect 869 1103 872 1107
rect 910 1092 913 1098
rect 850 1088 857 1091
rect 854 1072 857 1088
rect 878 1088 886 1091
rect 878 1072 881 1088
rect 826 1068 830 1071
rect 926 1062 929 1118
rect 934 1082 937 1098
rect 942 1072 945 1098
rect 1062 1092 1065 1128
rect 1070 1122 1073 1128
rect 1094 1102 1097 1158
rect 1238 1151 1241 1158
rect 1286 1152 1289 1188
rect 1494 1162 1497 1218
rect 1398 1152 1401 1158
rect 1110 1122 1113 1138
rect 1102 1082 1105 1118
rect 1118 1112 1121 1128
rect 1126 1112 1129 1118
rect 1134 1102 1137 1148
rect 1126 1082 1129 1088
rect 1134 1082 1137 1088
rect 934 1062 937 1068
rect 966 1062 969 1078
rect 738 1058 742 1061
rect 762 1058 766 1061
rect 726 1052 729 1058
rect 626 1048 630 1051
rect 746 1048 750 1051
rect 830 1042 833 1048
rect 614 962 617 968
rect 546 958 550 961
rect 574 952 577 958
rect 582 952 585 958
rect 538 948 542 951
rect 566 942 569 948
rect 622 942 625 1038
rect 846 1022 849 1058
rect 990 1052 993 1078
rect 1014 1062 1017 1078
rect 1046 1062 1049 1078
rect 1026 1048 1030 1051
rect 958 1042 961 1048
rect 1002 1038 1006 1041
rect 1034 1038 1038 1041
rect 1014 1032 1017 1038
rect 1046 1032 1049 1038
rect 682 1018 686 1021
rect 630 972 633 978
rect 650 968 654 971
rect 678 962 681 968
rect 638 952 641 958
rect 662 942 665 948
rect 550 932 553 938
rect 534 922 537 928
rect 558 922 561 928
rect 534 882 537 918
rect 614 892 617 898
rect 550 882 553 888
rect 558 882 561 888
rect 502 872 505 878
rect 542 871 545 878
rect 606 872 609 878
rect 638 872 641 938
rect 670 912 673 958
rect 710 952 713 1018
rect 722 948 726 951
rect 678 942 681 948
rect 710 922 713 938
rect 670 892 673 908
rect 650 878 654 881
rect 686 872 689 888
rect 702 882 705 898
rect 726 892 729 928
rect 734 902 737 918
rect 714 888 718 891
rect 730 888 737 891
rect 542 868 550 871
rect 494 862 497 868
rect 534 862 537 868
rect 586 858 590 861
rect 650 858 654 861
rect 690 858 694 861
rect 710 852 713 878
rect 734 872 737 888
rect 766 872 769 948
rect 730 858 734 861
rect 594 848 598 851
rect 618 848 622 851
rect 686 842 689 848
rect 194 818 201 821
rect 34 747 38 750
rect 130 748 134 751
rect 142 748 150 751
rect 178 748 182 751
rect 18 679 25 681
rect 14 678 25 679
rect 22 662 25 678
rect 46 671 49 738
rect 94 712 97 718
rect 102 702 105 738
rect 38 668 49 671
rect 54 679 62 681
rect 78 679 86 681
rect 54 678 65 679
rect 78 678 89 679
rect 22 531 25 548
rect 18 528 25 531
rect 38 542 41 668
rect 54 662 57 678
rect 78 662 81 678
rect 110 652 113 748
rect 126 661 129 718
rect 142 692 145 748
rect 150 742 153 748
rect 178 738 182 741
rect 134 662 137 668
rect 150 662 153 678
rect 158 672 161 738
rect 174 712 177 728
rect 190 712 193 748
rect 166 672 169 678
rect 198 672 201 818
rect 344 803 346 807
rect 350 803 353 807
rect 357 803 360 807
rect 638 792 641 818
rect 298 778 302 781
rect 346 768 353 771
rect 242 758 246 761
rect 206 742 209 758
rect 270 752 273 758
rect 218 748 222 751
rect 218 738 222 741
rect 238 722 241 728
rect 206 682 209 718
rect 230 702 233 718
rect 262 702 265 738
rect 318 732 321 738
rect 206 672 209 678
rect 214 672 217 688
rect 238 682 241 698
rect 278 692 281 708
rect 266 678 270 681
rect 186 668 190 671
rect 126 658 134 661
rect 194 658 198 661
rect 218 658 222 661
rect 230 652 233 668
rect 226 648 230 651
rect 62 572 65 588
rect 62 552 65 568
rect 38 512 41 538
rect 110 492 113 648
rect 222 592 225 628
rect 210 568 214 571
rect 182 562 185 568
rect 194 558 198 561
rect 118 512 121 518
rect 18 479 25 481
rect 14 478 25 479
rect 22 462 25 478
rect 54 479 62 481
rect 54 478 65 479
rect 54 462 57 478
rect 134 472 137 508
rect 142 502 145 548
rect 158 542 161 558
rect 238 552 241 668
rect 278 662 281 688
rect 262 652 265 658
rect 286 652 289 668
rect 294 662 297 668
rect 302 652 305 678
rect 326 672 329 758
rect 338 748 342 751
rect 350 742 353 768
rect 450 768 454 771
rect 474 768 478 771
rect 490 768 494 771
rect 690 768 694 771
rect 374 742 377 748
rect 334 732 337 738
rect 378 728 382 731
rect 334 712 337 728
rect 358 692 361 698
rect 390 682 393 758
rect 414 752 417 768
rect 438 742 441 748
rect 442 728 446 731
rect 398 692 401 728
rect 438 722 441 728
rect 446 702 449 718
rect 454 692 457 738
rect 482 728 489 731
rect 486 692 489 728
rect 398 672 401 688
rect 446 682 449 688
rect 494 682 497 768
rect 514 758 518 761
rect 502 752 505 758
rect 550 752 553 758
rect 514 748 518 751
rect 586 748 590 751
rect 502 732 505 738
rect 526 732 529 738
rect 554 728 558 731
rect 534 722 537 728
rect 542 692 545 728
rect 566 722 569 738
rect 590 732 593 738
rect 598 722 601 758
rect 766 752 769 868
rect 774 862 777 888
rect 790 862 793 1018
rect 846 972 849 978
rect 974 972 977 978
rect 990 972 993 1018
rect 1030 972 1033 978
rect 946 968 950 971
rect 962 968 966 971
rect 834 958 838 961
rect 798 951 801 958
rect 830 892 833 958
rect 850 938 854 941
rect 838 892 841 938
rect 856 903 858 907
rect 862 903 865 907
rect 869 903 872 907
rect 886 882 889 948
rect 902 942 905 948
rect 918 932 921 958
rect 930 948 937 951
rect 934 942 937 948
rect 942 892 945 948
rect 914 878 918 881
rect 862 872 865 878
rect 958 872 961 968
rect 978 958 982 961
rect 970 948 974 951
rect 982 881 985 958
rect 990 942 993 958
rect 998 952 1001 968
rect 1014 962 1017 968
rect 1046 962 1049 968
rect 1054 952 1057 1068
rect 1070 1062 1073 1078
rect 1142 1072 1145 1118
rect 1150 1072 1153 1108
rect 1158 1102 1161 1140
rect 1166 1122 1169 1138
rect 1234 1128 1238 1131
rect 1182 1122 1185 1128
rect 1094 1062 1097 1068
rect 1070 1052 1073 1058
rect 1102 1051 1105 1058
rect 1098 1048 1105 1051
rect 1110 1052 1113 1068
rect 1094 972 1097 1048
rect 1118 1032 1121 1068
rect 1142 1052 1145 1068
rect 1150 1062 1153 1068
rect 1174 1061 1177 1118
rect 1234 1078 1238 1081
rect 1198 1072 1201 1078
rect 1262 1072 1265 1098
rect 1286 1092 1289 1138
rect 1302 1132 1305 1148
rect 1334 1142 1337 1147
rect 1394 1128 1398 1131
rect 1366 1102 1369 1118
rect 1390 1092 1393 1118
rect 1274 1078 1278 1081
rect 1170 1058 1177 1061
rect 1166 1052 1169 1058
rect 1182 1042 1185 1068
rect 1310 1062 1313 1068
rect 1326 1062 1329 1078
rect 1398 1072 1401 1128
rect 1338 1068 1342 1071
rect 1202 1058 1206 1061
rect 1218 1058 1222 1061
rect 1346 1058 1350 1061
rect 1270 1052 1273 1058
rect 1302 1052 1305 1058
rect 1214 1042 1217 1048
rect 1230 982 1233 1018
rect 1206 962 1209 968
rect 1090 958 1094 961
rect 1034 948 1038 951
rect 1058 948 1062 951
rect 1094 942 1097 958
rect 1230 952 1233 958
rect 1246 952 1249 1018
rect 1110 942 1113 948
rect 1134 942 1137 948
rect 1174 942 1177 948
rect 1286 942 1289 1048
rect 1358 1032 1361 1048
rect 1368 1003 1370 1007
rect 1374 1003 1377 1007
rect 1381 1003 1384 1007
rect 1406 992 1409 1138
rect 1422 1122 1425 1138
rect 1438 1122 1441 1148
rect 1446 1142 1449 1148
rect 1454 1132 1457 1158
rect 1510 1142 1513 1148
rect 1566 1142 1569 1218
rect 1614 1192 1617 1268
rect 1638 1262 1641 1268
rect 1654 1262 1657 1268
rect 1626 1258 1630 1261
rect 1662 1252 1665 1258
rect 1642 1248 1646 1251
rect 1598 1172 1601 1178
rect 1610 1168 1614 1171
rect 1622 1142 1625 1148
rect 1586 1138 1590 1141
rect 1422 1052 1425 1058
rect 1430 1052 1433 1088
rect 1442 1068 1446 1071
rect 1454 1061 1457 1108
rect 1462 1092 1465 1138
rect 1450 1058 1457 1061
rect 1470 1052 1473 1058
rect 1414 1042 1417 1048
rect 1430 1042 1433 1048
rect 1414 1002 1417 1038
rect 1302 962 1305 988
rect 1430 972 1433 978
rect 1314 968 1318 971
rect 1446 971 1449 1018
rect 1462 1002 1465 1048
rect 1446 968 1457 971
rect 1454 962 1457 968
rect 1374 951 1377 958
rect 1414 942 1417 948
rect 1438 942 1441 948
rect 1446 942 1449 958
rect 994 938 1001 941
rect 982 878 990 881
rect 966 872 969 878
rect 854 852 857 858
rect 886 852 889 858
rect 918 852 921 868
rect 942 862 945 868
rect 946 848 950 851
rect 714 748 718 751
rect 798 751 801 758
rect 830 752 833 778
rect 814 742 817 748
rect 926 741 929 758
rect 922 738 929 741
rect 654 732 657 738
rect 662 722 665 738
rect 474 678 478 681
rect 310 662 313 668
rect 318 642 321 648
rect 270 592 273 638
rect 326 632 329 668
rect 358 662 361 668
rect 390 662 393 668
rect 406 652 409 678
rect 482 668 489 671
rect 426 658 430 661
rect 338 648 342 651
rect 362 648 366 651
rect 402 648 406 651
rect 434 648 438 651
rect 344 603 346 607
rect 350 603 353 607
rect 357 603 360 607
rect 322 548 326 551
rect 198 542 201 548
rect 222 542 225 548
rect 150 512 153 528
rect 158 492 161 538
rect 182 522 185 538
rect 238 532 241 548
rect 186 518 193 521
rect 190 472 193 518
rect 198 470 201 488
rect 66 348 70 351
rect 22 331 25 348
rect 18 328 25 331
rect 38 332 41 338
rect 78 322 81 468
rect 182 441 185 468
rect 222 462 225 488
rect 238 482 241 498
rect 246 482 249 518
rect 270 472 273 548
rect 278 462 281 538
rect 294 502 297 538
rect 390 492 393 638
rect 414 632 417 648
rect 414 592 417 618
rect 438 592 441 628
rect 470 622 473 658
rect 486 592 489 668
rect 522 668 526 671
rect 494 642 497 668
rect 526 662 529 668
rect 534 662 537 668
rect 550 662 553 708
rect 614 675 617 708
rect 630 692 633 718
rect 654 672 657 678
rect 702 672 705 678
rect 710 672 713 738
rect 870 732 873 738
rect 782 672 785 698
rect 790 692 793 728
rect 856 703 858 707
rect 862 703 865 707
rect 869 703 872 707
rect 902 702 905 718
rect 918 712 921 738
rect 930 718 934 721
rect 562 668 566 671
rect 586 668 590 671
rect 502 632 505 658
rect 590 652 593 658
rect 514 648 518 651
rect 530 648 534 651
rect 550 642 553 648
rect 518 592 521 638
rect 598 592 601 668
rect 806 652 809 698
rect 926 692 929 718
rect 934 692 937 708
rect 942 692 945 738
rect 950 712 953 738
rect 838 662 841 668
rect 818 658 822 661
rect 794 648 798 651
rect 646 592 649 638
rect 678 582 681 618
rect 566 572 569 578
rect 522 568 526 571
rect 634 568 638 571
rect 402 558 406 561
rect 414 492 417 548
rect 298 488 302 491
rect 350 488 358 491
rect 350 472 353 488
rect 422 482 425 498
rect 430 492 433 538
rect 462 532 465 558
rect 454 472 457 518
rect 462 482 465 498
rect 486 492 489 568
rect 506 558 510 561
rect 494 492 497 548
rect 510 532 513 558
rect 538 548 542 551
rect 518 542 521 548
rect 550 542 553 568
rect 642 548 646 551
rect 562 528 566 531
rect 462 472 465 478
rect 510 472 513 488
rect 526 472 529 498
rect 310 462 313 468
rect 398 462 401 468
rect 210 458 214 461
rect 266 458 270 461
rect 174 438 185 441
rect 310 442 313 458
rect 406 452 409 458
rect 446 452 449 458
rect 470 452 473 468
rect 554 458 558 461
rect 378 448 382 451
rect 490 448 494 451
rect 174 392 177 438
rect 344 403 346 407
rect 350 403 353 407
rect 357 403 360 407
rect 342 362 345 368
rect 134 342 137 348
rect 198 342 201 348
rect 214 342 217 358
rect 398 352 401 368
rect 242 348 246 351
rect 242 338 246 341
rect 22 262 25 318
rect 142 302 145 338
rect 174 332 178 335
rect 78 292 81 298
rect 66 268 70 271
rect 46 262 49 268
rect 130 258 134 261
rect 22 202 25 258
rect 38 242 41 248
rect 46 232 49 258
rect 102 252 105 258
rect 110 252 113 258
rect 166 252 169 258
rect 58 248 62 251
rect 82 248 86 251
rect 146 248 150 251
rect 90 218 94 221
rect 46 201 49 218
rect 46 198 57 201
rect 6 141 9 148
rect 6 138 14 141
rect 14 131 17 138
rect 30 132 33 148
rect 54 142 57 198
rect 102 192 105 248
rect 118 242 121 248
rect 190 242 193 338
rect 254 332 257 348
rect 310 342 313 348
rect 358 342 361 348
rect 498 347 502 350
rect 518 342 521 408
rect 574 372 577 538
rect 622 521 625 538
rect 618 518 625 521
rect 630 492 633 548
rect 606 482 609 488
rect 638 468 646 471
rect 626 458 630 461
rect 606 392 609 448
rect 566 362 569 368
rect 534 342 537 358
rect 542 342 545 348
rect 574 342 577 368
rect 598 362 601 368
rect 622 362 625 438
rect 630 362 633 448
rect 638 442 641 468
rect 582 352 585 358
rect 598 342 601 348
rect 294 332 297 340
rect 434 338 438 341
rect 562 338 566 341
rect 218 328 222 331
rect 230 312 233 318
rect 214 262 217 278
rect 226 268 230 271
rect 226 258 230 261
rect 238 261 241 278
rect 262 272 265 318
rect 270 312 273 328
rect 270 272 273 278
rect 278 271 281 318
rect 302 301 305 338
rect 298 298 305 301
rect 286 282 289 288
rect 274 268 281 271
rect 294 272 297 298
rect 310 272 313 328
rect 406 302 409 332
rect 350 282 353 298
rect 322 278 326 281
rect 262 262 265 268
rect 238 258 246 261
rect 274 258 278 261
rect 298 258 302 261
rect 246 252 249 258
rect 310 252 313 268
rect 338 258 342 261
rect 350 252 353 278
rect 414 272 417 288
rect 422 282 425 298
rect 422 272 425 278
rect 78 172 81 178
rect 118 172 121 238
rect 134 212 137 238
rect 90 168 94 171
rect 118 158 126 161
rect 118 152 121 158
rect 142 152 145 218
rect 150 192 153 228
rect 318 222 321 248
rect 358 242 361 268
rect 370 258 374 261
rect 398 242 401 248
rect 386 238 390 241
rect 166 182 169 218
rect 190 162 193 218
rect 214 192 217 208
rect 270 192 273 198
rect 230 162 233 178
rect 54 112 57 128
rect 30 79 38 81
rect 30 78 41 79
rect 30 62 33 78
rect 62 62 65 138
rect 70 62 73 108
rect 94 92 97 148
rect 118 132 121 148
rect 158 142 161 158
rect 182 152 185 158
rect 150 138 158 141
rect 126 122 129 128
rect 150 92 153 138
rect 166 92 169 138
rect 238 131 241 188
rect 230 128 241 131
rect 246 142 249 148
rect 254 142 257 148
rect 310 142 313 218
rect 318 182 321 218
rect 334 162 337 208
rect 344 203 346 207
rect 350 203 353 207
rect 357 203 360 207
rect 334 152 337 158
rect 366 152 369 178
rect 390 172 393 218
rect 430 171 433 308
rect 438 302 441 318
rect 446 292 449 338
rect 478 272 481 278
rect 518 272 521 338
rect 534 332 537 338
rect 582 332 585 338
rect 598 292 601 338
rect 606 332 609 348
rect 630 332 633 358
rect 646 332 649 458
rect 654 422 657 558
rect 678 552 681 578
rect 686 542 689 548
rect 686 512 689 538
rect 694 532 697 538
rect 702 531 705 618
rect 766 612 769 618
rect 798 592 801 628
rect 838 621 841 658
rect 846 632 849 668
rect 870 662 873 678
rect 954 668 958 671
rect 886 662 889 668
rect 858 658 862 661
rect 886 622 889 658
rect 902 652 905 668
rect 966 662 969 868
rect 974 862 977 868
rect 990 862 993 868
rect 998 852 1001 938
rect 1266 938 1270 941
rect 1038 932 1041 938
rect 1078 932 1081 938
rect 1094 902 1097 918
rect 1102 892 1105 918
rect 1134 912 1137 928
rect 1134 882 1137 898
rect 1142 882 1145 938
rect 1150 912 1153 928
rect 1166 912 1169 928
rect 1150 892 1153 898
rect 1078 872 1081 878
rect 1050 858 1054 861
rect 1006 832 1009 858
rect 1022 842 1025 848
rect 1038 842 1041 858
rect 1062 852 1065 868
rect 1078 852 1081 858
rect 1006 752 1009 808
rect 1014 802 1017 838
rect 1046 832 1049 848
rect 1054 762 1057 768
rect 1062 752 1065 848
rect 1078 832 1081 848
rect 1086 842 1089 868
rect 1102 852 1105 868
rect 1158 862 1161 868
rect 1166 862 1169 868
rect 1174 862 1177 878
rect 1198 872 1201 908
rect 1206 872 1209 932
rect 1222 902 1225 938
rect 1246 922 1249 938
rect 1238 912 1241 918
rect 1234 878 1238 881
rect 1198 862 1201 868
rect 1214 862 1217 878
rect 1246 872 1249 918
rect 1098 848 1102 851
rect 1110 842 1113 858
rect 1230 852 1233 858
rect 1238 852 1241 868
rect 1254 862 1257 938
rect 1270 922 1273 928
rect 1278 912 1281 928
rect 1278 872 1281 878
rect 1266 868 1270 871
rect 1286 852 1289 938
rect 1302 902 1305 918
rect 1302 882 1305 898
rect 1318 872 1321 878
rect 1326 862 1329 908
rect 1390 892 1393 938
rect 1454 922 1457 948
rect 1470 942 1473 1038
rect 1478 1032 1481 1058
rect 1486 1032 1489 1038
rect 1478 992 1481 1028
rect 1494 1021 1497 1118
rect 1518 1102 1521 1138
rect 1502 1052 1505 1078
rect 1526 1072 1529 1098
rect 1510 1052 1513 1058
rect 1534 1022 1537 1118
rect 1574 1112 1577 1128
rect 1550 1082 1553 1088
rect 1550 1062 1553 1068
rect 1558 1062 1561 1098
rect 1598 1082 1601 1098
rect 1570 1068 1574 1071
rect 1586 1058 1590 1061
rect 1606 1042 1609 1118
rect 1614 1062 1617 1138
rect 1630 1092 1633 1158
rect 1638 1142 1641 1148
rect 1646 1142 1649 1168
rect 1686 1162 1689 1278
rect 1742 1272 1745 1338
rect 1814 1332 1817 1338
rect 1914 1328 1918 1331
rect 1806 1322 1809 1328
rect 1872 1303 1874 1307
rect 1878 1303 1881 1307
rect 1885 1303 1888 1307
rect 1846 1282 1849 1298
rect 1762 1278 1766 1281
rect 1790 1272 1793 1278
rect 1838 1272 1841 1278
rect 1746 1268 1750 1271
rect 1694 1232 1697 1268
rect 1774 1262 1777 1268
rect 1782 1262 1785 1268
rect 1706 1258 1710 1261
rect 1754 1258 1758 1261
rect 1846 1261 1849 1278
rect 1854 1272 1857 1278
rect 1894 1272 1897 1318
rect 1918 1292 1921 1318
rect 1926 1292 1929 1328
rect 1942 1301 1945 1388
rect 2030 1362 2033 1368
rect 2038 1352 2041 1398
rect 2110 1382 2113 1478
rect 2118 1472 2121 1488
rect 2130 1468 2134 1471
rect 2162 1468 2166 1471
rect 2134 1442 2137 1448
rect 2150 1432 2153 1468
rect 2174 1432 2177 1468
rect 2182 1452 2185 1478
rect 2198 1462 2201 1538
rect 2214 1482 2217 1628
rect 2222 1592 2225 1668
rect 2230 1662 2233 1668
rect 2270 1662 2273 1678
rect 2278 1672 2281 1718
rect 2302 1712 2305 1738
rect 2310 1702 2313 1738
rect 2342 1732 2345 1738
rect 2358 1722 2361 1738
rect 2374 1732 2377 1758
rect 2378 1728 2382 1731
rect 2294 1682 2297 1688
rect 2366 1672 2369 1718
rect 2390 1692 2393 1768
rect 2422 1742 2425 1748
rect 2430 1742 2433 1818
rect 2438 1772 2441 1848
rect 2470 1812 2473 1878
rect 2574 1862 2577 1918
rect 2498 1858 2502 1861
rect 2530 1858 2534 1861
rect 2562 1858 2566 1861
rect 2582 1861 2585 1958
rect 2642 1948 2646 1951
rect 2718 1942 2721 2118
rect 2726 2082 2729 2098
rect 2726 2052 2729 2078
rect 2790 2072 2793 2118
rect 2806 2082 2809 2118
rect 2838 2092 2841 2138
rect 2854 2092 2857 2148
rect 2870 2082 2873 2158
rect 2886 2142 2889 2178
rect 2898 2158 2902 2161
rect 2926 2152 2929 2218
rect 2942 2192 2945 2198
rect 2998 2192 3001 2338
rect 3054 2332 3057 2338
rect 3062 2332 3065 2358
rect 3074 2338 3078 2341
rect 3014 2312 3017 2328
rect 3102 2322 3105 2338
rect 3118 2322 3121 2338
rect 3150 2332 3153 2358
rect 3174 2352 3177 2388
rect 3214 2372 3217 2388
rect 3234 2368 3238 2371
rect 3198 2362 3201 2368
rect 3206 2352 3209 2358
rect 3246 2352 3249 2368
rect 3254 2362 3257 2368
rect 3262 2362 3265 2378
rect 3278 2362 3281 2368
rect 3326 2362 3329 2368
rect 3358 2362 3361 2378
rect 3370 2368 3377 2371
rect 3314 2358 3318 2361
rect 3346 2358 3350 2361
rect 3362 2358 3366 2361
rect 3274 2348 3278 2351
rect 3322 2348 3326 2351
rect 3362 2348 3366 2351
rect 3166 2342 3169 2348
rect 3190 2342 3193 2348
rect 3374 2342 3377 2368
rect 3382 2362 3385 2418
rect 3398 2352 3401 2558
rect 3542 2551 3545 2558
rect 3406 2502 3409 2538
rect 3430 2512 3433 2528
rect 3434 2508 3441 2511
rect 3414 2482 3417 2498
rect 3406 2472 3409 2478
rect 3438 2472 3441 2508
rect 3446 2482 3449 2548
rect 3458 2528 3462 2531
rect 3470 2512 3473 2518
rect 3478 2502 3481 2548
rect 3550 2542 3553 2668
rect 3630 2622 3633 2668
rect 3638 2662 3641 2718
rect 3646 2702 3649 2738
rect 3654 2722 3657 2748
rect 3662 2721 3665 2758
rect 3678 2751 3681 2758
rect 3674 2748 3681 2751
rect 3686 2741 3689 2768
rect 3706 2758 3710 2761
rect 3694 2752 3697 2758
rect 3706 2748 3710 2751
rect 3678 2738 3689 2741
rect 3662 2718 3673 2721
rect 3662 2692 3665 2708
rect 3646 2672 3649 2678
rect 3670 2672 3673 2718
rect 3678 2712 3681 2738
rect 3718 2732 3721 2738
rect 3734 2732 3737 2768
rect 3782 2762 3785 2818
rect 3886 2792 3889 2868
rect 3918 2842 3921 2878
rect 3950 2872 3953 2918
rect 3958 2871 3961 2948
rect 4134 2942 4137 2958
rect 4218 2948 4222 2951
rect 4082 2938 4086 2941
rect 3966 2882 3969 2938
rect 3974 2922 3977 2928
rect 3982 2892 3985 2938
rect 4038 2912 4041 2938
rect 4046 2932 4049 2938
rect 4074 2928 4078 2931
rect 4046 2892 4049 2928
rect 4054 2892 4057 2908
rect 4014 2872 4017 2878
rect 4078 2872 4081 2918
rect 4142 2912 4145 2928
rect 4158 2922 4161 2938
rect 4086 2882 4089 2888
rect 4094 2882 4097 2888
rect 3958 2868 3966 2871
rect 3958 2862 3961 2868
rect 3970 2858 3974 2861
rect 3942 2842 3945 2848
rect 3974 2842 3977 2848
rect 3990 2832 3993 2868
rect 3998 2842 4001 2868
rect 4038 2862 4041 2868
rect 3998 2822 4001 2838
rect 4014 2832 4017 2848
rect 4022 2842 4025 2848
rect 4030 2832 4033 2858
rect 4042 2838 4046 2841
rect 3798 2772 3801 2778
rect 3850 2758 3854 2761
rect 3742 2752 3745 2758
rect 3750 2732 3753 2748
rect 3782 2732 3785 2758
rect 3814 2752 3817 2758
rect 3842 2748 3846 2751
rect 3798 2742 3801 2748
rect 3822 2742 3825 2748
rect 3686 2692 3689 2728
rect 3782 2722 3785 2728
rect 3790 2721 3793 2738
rect 3846 2732 3849 2738
rect 3790 2718 3798 2721
rect 3726 2672 3729 2708
rect 3790 2688 3798 2691
rect 3782 2682 3785 2688
rect 3790 2672 3793 2688
rect 3658 2648 3662 2651
rect 3682 2648 3686 2651
rect 3646 2642 3649 2648
rect 3606 2592 3609 2598
rect 3702 2592 3705 2668
rect 3718 2652 3721 2659
rect 3714 2588 3718 2591
rect 3574 2552 3577 2558
rect 3670 2552 3673 2558
rect 3726 2552 3729 2668
rect 3806 2661 3809 2698
rect 3814 2692 3817 2728
rect 3838 2712 3841 2728
rect 3854 2692 3857 2738
rect 3862 2692 3865 2748
rect 3870 2732 3873 2738
rect 3886 2732 3889 2768
rect 3894 2742 3897 2748
rect 3942 2742 3945 2748
rect 3928 2703 3930 2707
rect 3934 2703 3937 2707
rect 3941 2703 3944 2707
rect 3802 2658 3809 2661
rect 3822 2672 3825 2678
rect 3834 2668 3838 2671
rect 3822 2652 3825 2668
rect 3878 2662 3881 2698
rect 3894 2672 3897 2688
rect 3910 2682 3913 2698
rect 3950 2692 3953 2808
rect 4014 2792 4017 2818
rect 4030 2812 4033 2828
rect 4078 2812 4081 2868
rect 4086 2862 4089 2878
rect 4110 2862 4113 2868
rect 4110 2832 4113 2848
rect 4118 2842 4121 2888
rect 4134 2862 4137 2868
rect 4142 2861 4145 2878
rect 4150 2872 4153 2878
rect 4166 2872 4169 2948
rect 4214 2942 4217 2948
rect 4246 2942 4249 2948
rect 4294 2942 4297 3008
rect 4318 3002 4321 3028
rect 4302 2952 4305 2998
rect 4326 2952 4329 3048
rect 4334 3042 4337 3058
rect 4342 3052 4345 3058
rect 4414 3052 4417 3058
rect 4430 3052 4433 3058
rect 4382 2992 4385 3038
rect 4326 2942 4329 2948
rect 4350 2942 4353 2948
rect 4142 2858 4150 2861
rect 4038 2792 4041 2808
rect 4090 2788 4094 2791
rect 4134 2782 4137 2858
rect 4174 2852 4177 2858
rect 4142 2842 4145 2848
rect 4166 2792 4169 2848
rect 4190 2822 4193 2858
rect 4198 2852 4201 2868
rect 3970 2768 3974 2771
rect 4026 2768 4030 2771
rect 4046 2762 4049 2778
rect 4062 2762 4065 2768
rect 4098 2758 4102 2761
rect 3966 2742 3969 2758
rect 3982 2752 3985 2758
rect 3998 2752 4001 2758
rect 4042 2748 4046 2751
rect 3982 2742 3985 2748
rect 4054 2742 4057 2748
rect 4094 2742 4097 2748
rect 4102 2742 4105 2758
rect 4142 2751 4145 2758
rect 4206 2752 4209 2918
rect 4326 2892 4329 2938
rect 4406 2901 4409 2938
rect 4414 2932 4417 2940
rect 4406 2898 4414 2901
rect 4226 2888 4230 2891
rect 4218 2868 4222 2871
rect 4270 2822 4273 2868
rect 4278 2862 4281 2868
rect 4290 2848 4294 2851
rect 4310 2812 4313 2858
rect 4342 2772 4345 2868
rect 4358 2802 4361 2858
rect 4430 2792 4433 3048
rect 4478 3042 4481 3058
rect 4494 3042 4497 3058
rect 4542 3052 4545 3068
rect 4590 3062 4593 3068
rect 4622 3063 4625 3068
rect 4440 3003 4442 3007
rect 4446 3003 4449 3007
rect 4453 3003 4456 3007
rect 4506 2968 4510 2971
rect 4546 2968 4553 2971
rect 4542 2962 4545 2968
rect 4442 2958 4446 2961
rect 4494 2952 4497 2958
rect 4458 2938 4462 2941
rect 4470 2932 4473 2948
rect 4518 2942 4521 2958
rect 4526 2942 4529 2948
rect 4438 2892 4441 2918
rect 4454 2892 4457 2928
rect 4470 2892 4473 2928
rect 4478 2922 4481 2938
rect 4550 2932 4553 2968
rect 4574 2952 4577 2958
rect 4562 2938 4566 2941
rect 4502 2922 4505 2928
rect 4446 2888 4454 2891
rect 4446 2872 4449 2888
rect 4494 2882 4497 2918
rect 4542 2892 4545 2918
rect 4550 2882 4553 2898
rect 4542 2878 4550 2881
rect 4494 2832 4497 2868
rect 4542 2862 4545 2878
rect 4558 2872 4561 2928
rect 4590 2872 4593 2918
rect 4598 2862 4601 2878
rect 4440 2803 4442 2807
rect 4446 2803 4449 2807
rect 4453 2803 4456 2807
rect 4518 2792 4521 2858
rect 4606 2852 4609 2918
rect 4614 2892 4617 2948
rect 4638 2942 4641 3088
rect 4646 3072 4649 3138
rect 4694 3132 4697 3138
rect 4750 3122 4753 3128
rect 4686 3092 4689 3098
rect 4694 3082 4697 3098
rect 4790 3092 4793 3138
rect 4742 3072 4745 3088
rect 4830 3072 4833 3088
rect 4846 3072 4849 3078
rect 4854 3072 4857 3088
rect 4714 3068 4718 3071
rect 4846 3062 4849 3068
rect 4862 3062 4865 3148
rect 4730 3058 4734 3061
rect 4830 3052 4833 3058
rect 4870 3052 4873 3108
rect 4910 3092 4913 3218
rect 4982 3182 4985 3248
rect 5014 3242 5017 3248
rect 5062 3232 5065 3268
rect 5086 3262 5089 3268
rect 5070 3242 5073 3248
rect 5094 3242 5097 3268
rect 5110 3262 5113 3278
rect 5206 3272 5209 3278
rect 5130 3268 5134 3271
rect 5154 3268 5166 3271
rect 5106 3258 5110 3261
rect 5170 3258 5174 3261
rect 5182 3258 5190 3261
rect 4918 3152 4921 3158
rect 4938 3148 4942 3151
rect 4918 3132 4921 3138
rect 4934 3052 4937 3148
rect 4946 3138 4950 3141
rect 4942 3122 4945 3128
rect 4950 3122 4953 3128
rect 4942 3072 4945 3108
rect 4952 3103 4954 3107
rect 4958 3103 4961 3107
rect 4965 3103 4968 3107
rect 4950 3062 4953 3078
rect 4958 3062 4961 3088
rect 4946 3058 4950 3061
rect 4818 3048 4822 3051
rect 4750 2952 4753 3048
rect 4850 2988 4854 2991
rect 4738 2948 4742 2951
rect 4782 2951 4785 2958
rect 4702 2942 4705 2948
rect 4710 2922 4713 2948
rect 4886 2942 4889 2948
rect 4766 2932 4769 2938
rect 4638 2882 4641 2918
rect 4726 2912 4729 2928
rect 4614 2862 4617 2878
rect 4622 2852 4625 2868
rect 4638 2862 4641 2868
rect 4574 2842 4577 2848
rect 4662 2842 4665 2858
rect 4670 2852 4673 2888
rect 4698 2868 4702 2871
rect 4730 2868 4734 2871
rect 4750 2862 4753 2888
rect 4854 2882 4857 2918
rect 4774 2862 4777 2878
rect 4790 2872 4793 2878
rect 4854 2872 4857 2878
rect 4790 2862 4793 2868
rect 4690 2858 4694 2861
rect 4722 2858 4726 2861
rect 4814 2852 4817 2868
rect 4830 2852 4833 2868
rect 4870 2862 4873 2940
rect 4886 2922 4889 2938
rect 4878 2882 4881 2898
rect 4886 2872 4889 2878
rect 4902 2862 4905 2958
rect 4934 2951 4937 3048
rect 4950 2952 4953 3058
rect 4934 2948 4942 2951
rect 4954 2938 4958 2941
rect 4974 2932 4977 3118
rect 4986 3068 4990 3071
rect 4998 2992 5001 3228
rect 5022 3132 5025 3148
rect 5030 3142 5033 3168
rect 5006 3062 5009 3088
rect 5038 3082 5041 3118
rect 5070 3072 5073 3168
rect 5078 3162 5081 3168
rect 5094 3152 5097 3178
rect 5086 3082 5089 3148
rect 5034 3068 5038 3071
rect 5022 3062 5025 3068
rect 5030 3052 5033 3058
rect 5086 3052 5089 3059
rect 5030 2992 5033 3048
rect 4998 2952 5001 2988
rect 5054 2972 5057 2978
rect 5102 2952 5105 3258
rect 5118 3232 5121 3258
rect 5182 3251 5185 3258
rect 5162 3248 5185 3251
rect 5198 3252 5201 3268
rect 5214 3262 5217 3268
rect 5238 3262 5241 3308
rect 5262 3292 5265 3318
rect 5258 3279 5265 3281
rect 5254 3278 5265 3279
rect 5262 3262 5265 3278
rect 5270 3252 5273 3258
rect 5278 3231 5281 3318
rect 5286 3282 5289 3298
rect 5294 3262 5297 3348
rect 5310 3312 5313 3338
rect 5278 3228 5286 3231
rect 5246 3172 5249 3178
rect 5198 3152 5201 3158
rect 5270 3151 5273 3188
rect 5278 3182 5281 3218
rect 5290 3158 5294 3161
rect 5270 3148 5278 3151
rect 5126 3142 5129 3148
rect 4986 2948 4990 2951
rect 5058 2948 5062 2951
rect 5074 2948 5078 2951
rect 5006 2932 5009 2938
rect 4954 2918 4958 2921
rect 4910 2882 4913 2918
rect 4952 2903 4954 2907
rect 4958 2903 4961 2907
rect 4965 2903 4968 2907
rect 5038 2892 5041 2948
rect 5118 2932 5121 3118
rect 5134 2992 5137 3148
rect 5214 3142 5217 3148
rect 5142 3122 5145 3128
rect 5146 3088 5150 3091
rect 5182 3063 5185 3118
rect 5238 3102 5241 3148
rect 5262 3142 5265 3148
rect 5246 3092 5249 3138
rect 5270 3131 5273 3138
rect 5262 3128 5273 3131
rect 5134 2952 5137 2988
rect 5166 2952 5169 2958
rect 5198 2951 5201 2958
rect 5070 2882 5073 2898
rect 5078 2892 5081 2898
rect 4918 2872 4921 2878
rect 4942 2862 4945 2878
rect 4866 2858 4870 2861
rect 4854 2851 4857 2858
rect 4854 2848 4865 2851
rect 4586 2838 4590 2841
rect 4650 2838 4654 2841
rect 4598 2832 4601 2838
rect 4566 2792 4569 2828
rect 4390 2772 4393 2778
rect 4414 2772 4417 2778
rect 4402 2768 4406 2771
rect 4358 2762 4361 2768
rect 4598 2762 4601 2768
rect 4450 2758 4454 2761
rect 4506 2758 4510 2761
rect 4430 2752 4433 2758
rect 4142 2748 4150 2751
rect 4058 2738 4065 2741
rect 3958 2722 3961 2738
rect 4054 2672 4057 2708
rect 3918 2662 3921 2668
rect 4062 2662 4065 2738
rect 4138 2738 4142 2741
rect 4070 2712 4073 2728
rect 4078 2692 4081 2738
rect 4126 2681 4129 2728
rect 4118 2678 4129 2681
rect 4086 2672 4089 2678
rect 4094 2662 4097 2668
rect 3838 2652 3841 2658
rect 3862 2652 3865 2658
rect 3930 2648 3934 2651
rect 3854 2642 3857 2648
rect 3902 2642 3905 2648
rect 3982 2632 3985 2659
rect 4014 2642 4017 2658
rect 4074 2648 4078 2651
rect 3642 2547 3646 2550
rect 3462 2492 3465 2498
rect 3470 2482 3473 2498
rect 3446 2462 3449 2478
rect 3550 2472 3553 2488
rect 3482 2468 3486 2471
rect 3534 2462 3537 2468
rect 3522 2458 3526 2461
rect 3538 2448 3542 2451
rect 3494 2442 3497 2448
rect 3526 2442 3529 2448
rect 3558 2442 3561 2478
rect 3574 2472 3577 2508
rect 3598 2482 3601 2488
rect 3654 2482 3657 2498
rect 3630 2472 3633 2478
rect 3566 2462 3569 2468
rect 3626 2458 3630 2461
rect 3650 2458 3654 2461
rect 3582 2452 3585 2458
rect 3606 2452 3609 2458
rect 3638 2452 3641 2458
rect 3662 2451 3665 2538
rect 3742 2532 3745 2538
rect 3774 2502 3777 2548
rect 3814 2531 3817 2548
rect 3838 2542 3841 2578
rect 3858 2558 3862 2561
rect 3810 2528 3817 2531
rect 3822 2522 3825 2528
rect 3670 2472 3673 2478
rect 3686 2462 3689 2478
rect 3734 2462 3737 2478
rect 3782 2472 3785 2518
rect 3822 2472 3825 2478
rect 3798 2462 3801 2468
rect 3654 2448 3665 2451
rect 3718 2452 3721 2458
rect 3506 2438 3510 2441
rect 3398 2342 3401 2348
rect 3282 2338 3286 2341
rect 3314 2338 3318 2341
rect 3158 2332 3161 2338
rect 3246 2332 3249 2338
rect 3294 2332 3297 2338
rect 3186 2328 3190 2331
rect 3006 2292 3009 2308
rect 3006 2282 3009 2288
rect 3070 2282 3073 2318
rect 3014 2252 3017 2268
rect 3062 2241 3065 2268
rect 3070 2252 3073 2278
rect 3086 2262 3089 2288
rect 3102 2282 3105 2318
rect 3134 2272 3137 2318
rect 3142 2312 3145 2328
rect 3206 2322 3209 2328
rect 3098 2268 3102 2271
rect 3098 2258 3102 2261
rect 3118 2251 3121 2268
rect 3142 2262 3145 2288
rect 3130 2258 3134 2261
rect 3150 2251 3153 2318
rect 3166 2272 3169 2278
rect 3214 2272 3217 2318
rect 3222 2272 3225 2288
rect 3274 2268 3278 2271
rect 3294 2262 3297 2268
rect 3302 2261 3305 2318
rect 3310 2282 3313 2328
rect 3358 2292 3361 2338
rect 3386 2328 3390 2331
rect 3366 2292 3369 2318
rect 3382 2292 3385 2318
rect 3406 2292 3409 2428
rect 3526 2422 3529 2438
rect 3416 2403 3418 2407
rect 3422 2403 3425 2407
rect 3429 2403 3432 2407
rect 3454 2392 3457 2398
rect 3518 2372 3521 2418
rect 3478 2362 3481 2368
rect 3494 2352 3497 2358
rect 3494 2342 3497 2348
rect 3418 2338 3422 2341
rect 3470 2332 3473 2338
rect 3510 2322 3513 2368
rect 3518 2362 3521 2368
rect 3522 2348 3526 2351
rect 3582 2342 3585 2388
rect 3622 2362 3625 2418
rect 3618 2348 3622 2351
rect 3590 2342 3593 2348
rect 3638 2342 3641 2428
rect 3646 2352 3649 2358
rect 3530 2338 3534 2341
rect 3518 2332 3521 2338
rect 3610 2318 3614 2321
rect 3478 2282 3481 2318
rect 3526 2292 3529 2308
rect 3550 2302 3553 2318
rect 3534 2288 3542 2291
rect 3554 2288 3558 2291
rect 3418 2278 3422 2281
rect 3534 2272 3537 2288
rect 3582 2272 3585 2278
rect 3590 2272 3593 2278
rect 3638 2272 3641 2298
rect 3298 2258 3305 2261
rect 3370 2268 3374 2271
rect 3642 2268 3649 2271
rect 3326 2252 3329 2268
rect 3118 2248 3129 2251
rect 3150 2248 3158 2251
rect 3062 2238 3073 2241
rect 3046 2182 3049 2218
rect 3070 2192 3073 2238
rect 3126 2192 3129 2248
rect 3286 2242 3289 2248
rect 3334 2232 3337 2258
rect 3382 2252 3385 2268
rect 3390 2262 3393 2268
rect 3362 2248 3366 2251
rect 3186 2218 3190 2221
rect 3142 2202 3145 2218
rect 3182 2168 3198 2171
rect 3202 2168 3217 2171
rect 3066 2158 3070 2161
rect 3042 2148 3046 2151
rect 2894 2092 2897 2148
rect 3054 2142 3057 2158
rect 3078 2152 3081 2168
rect 3134 2152 3137 2168
rect 3182 2161 3185 2168
rect 3214 2162 3217 2168
rect 3154 2158 3185 2161
rect 3202 2158 3206 2161
rect 3234 2158 3238 2161
rect 3066 2148 3070 2151
rect 3146 2148 3158 2151
rect 2926 2132 2929 2138
rect 2974 2132 2977 2138
rect 2982 2132 2985 2138
rect 2922 2118 2929 2121
rect 2904 2103 2906 2107
rect 2910 2103 2913 2107
rect 2917 2103 2920 2107
rect 2926 2082 2929 2118
rect 3030 2102 3033 2138
rect 3038 2122 3041 2138
rect 3054 2092 3057 2138
rect 3070 2132 3073 2148
rect 3118 2142 3121 2148
rect 3098 2138 3102 2141
rect 3142 2132 3145 2148
rect 3162 2138 3166 2141
rect 3190 2132 3193 2158
rect 3210 2148 3214 2151
rect 3226 2148 3230 2151
rect 3246 2142 3249 2208
rect 3254 2162 3257 2218
rect 3270 2161 3273 2168
rect 3262 2158 3273 2161
rect 3262 2152 3265 2158
rect 3274 2148 3278 2151
rect 3286 2142 3289 2148
rect 3294 2142 3297 2218
rect 3366 2172 3369 2198
rect 3382 2162 3385 2238
rect 3390 2152 3393 2258
rect 3398 2222 3401 2268
rect 3474 2258 3478 2261
rect 3416 2203 3418 2207
rect 3422 2203 3425 2207
rect 3429 2203 3432 2207
rect 3406 2162 3409 2198
rect 3306 2148 3310 2151
rect 3322 2148 3326 2151
rect 3378 2148 3385 2151
rect 3334 2142 3337 2148
rect 3234 2138 3238 2141
rect 3266 2138 3270 2141
rect 3094 2112 3097 2128
rect 3046 2082 3049 2088
rect 2770 2068 2774 2071
rect 2794 2068 2798 2071
rect 2742 2062 2745 2068
rect 2822 2062 2825 2068
rect 2830 2062 2833 2068
rect 2762 2058 2766 2061
rect 2794 2058 2798 2061
rect 2770 2048 2774 2051
rect 2782 2042 2785 2058
rect 2854 2052 2857 2078
rect 2926 2072 2929 2078
rect 2842 2048 2846 2051
rect 2726 1951 2729 1998
rect 2798 1992 2801 2048
rect 2838 2002 2841 2048
rect 2854 2041 2857 2048
rect 2846 2038 2857 2041
rect 2782 1952 2785 1958
rect 2590 1921 2593 1938
rect 2590 1918 2598 1921
rect 2602 1878 2606 1881
rect 2590 1862 2593 1868
rect 2582 1858 2590 1861
rect 2506 1848 2510 1851
rect 2522 1838 2526 1841
rect 2534 1822 2537 1848
rect 2566 1842 2569 1848
rect 2554 1838 2558 1841
rect 2446 1742 2449 1768
rect 2462 1762 2465 1768
rect 2478 1752 2481 1818
rect 2558 1781 2561 1818
rect 2558 1778 2569 1781
rect 2542 1768 2550 1771
rect 2554 1768 2558 1771
rect 2458 1748 2462 1751
rect 2478 1742 2481 1748
rect 2502 1742 2505 1748
rect 2430 1732 2433 1738
rect 2422 1721 2425 1728
rect 2438 1721 2441 1738
rect 2486 1732 2489 1738
rect 2510 1732 2513 1738
rect 2518 1732 2521 1758
rect 2542 1752 2545 1768
rect 2566 1762 2569 1778
rect 2582 1762 2585 1768
rect 2550 1752 2553 1758
rect 2566 1752 2569 1758
rect 2574 1752 2577 1758
rect 2598 1752 2601 1868
rect 2606 1822 2609 1848
rect 2614 1792 2617 1918
rect 2630 1872 2633 1898
rect 2638 1892 2641 1938
rect 2718 1902 2721 1938
rect 2662 1872 2665 1898
rect 2694 1892 2697 1898
rect 2690 1878 2694 1881
rect 2718 1872 2721 1878
rect 2622 1862 2625 1868
rect 2654 1862 2657 1868
rect 2670 1862 2673 1868
rect 2706 1866 2710 1869
rect 2658 1858 2665 1861
rect 2630 1852 2633 1858
rect 2642 1848 2646 1851
rect 2662 1851 2665 1858
rect 2726 1852 2729 1898
rect 2734 1872 2737 1908
rect 2758 1892 2761 1948
rect 2798 1932 2801 1948
rect 2806 1942 2809 1948
rect 2814 1942 2817 1948
rect 2830 1942 2833 1948
rect 2818 1928 2822 1931
rect 2830 1922 2833 1928
rect 2766 1892 2769 1898
rect 2798 1882 2801 1908
rect 2806 1882 2809 1908
rect 2814 1892 2817 1898
rect 2738 1858 2742 1861
rect 2750 1852 2753 1868
rect 2662 1848 2673 1851
rect 2670 1842 2673 1848
rect 2758 1841 2761 1878
rect 2774 1862 2777 1868
rect 2782 1852 2785 1858
rect 2750 1838 2761 1841
rect 2638 1792 2641 1818
rect 2646 1762 2649 1768
rect 2634 1758 2638 1761
rect 2674 1748 2678 1751
rect 2538 1738 2542 1741
rect 2530 1728 2534 1731
rect 2422 1718 2441 1721
rect 2414 1682 2417 1718
rect 2462 1712 2465 1718
rect 2446 1692 2449 1698
rect 2558 1692 2561 1728
rect 2566 1722 2569 1748
rect 2582 1742 2585 1748
rect 2598 1742 2601 1748
rect 2606 1742 2609 1748
rect 2614 1731 2617 1748
rect 2606 1728 2617 1731
rect 2686 1741 2689 1838
rect 2718 1762 2721 1828
rect 2678 1738 2689 1741
rect 2718 1741 2721 1758
rect 2714 1738 2721 1741
rect 2742 1751 2745 1818
rect 2734 1748 2745 1751
rect 2750 1752 2753 1838
rect 2726 1742 2729 1748
rect 2646 1732 2649 1738
rect 2658 1728 2662 1731
rect 2574 1692 2577 1698
rect 2606 1692 2609 1728
rect 2534 1682 2537 1688
rect 2598 1682 2601 1688
rect 2398 1678 2406 1681
rect 2506 1678 2510 1681
rect 2554 1678 2558 1681
rect 2374 1672 2377 1678
rect 2398 1672 2401 1678
rect 2678 1672 2681 1738
rect 2734 1732 2737 1748
rect 2706 1728 2710 1731
rect 2694 1692 2697 1728
rect 2742 1722 2745 1738
rect 2750 1732 2753 1748
rect 2346 1668 2350 1671
rect 2474 1668 2478 1671
rect 2522 1668 2526 1671
rect 2246 1612 2249 1658
rect 2270 1652 2273 1658
rect 2326 1652 2329 1658
rect 2342 1652 2345 1658
rect 2306 1648 2310 1651
rect 2386 1648 2390 1651
rect 2258 1588 2262 1591
rect 2294 1582 2297 1618
rect 2314 1588 2318 1591
rect 2226 1548 2230 1551
rect 2246 1532 2249 1578
rect 2350 1572 2353 1608
rect 2298 1568 2302 1571
rect 2366 1562 2369 1648
rect 2382 1602 2385 1648
rect 2398 1622 2401 1668
rect 2406 1652 2409 1668
rect 2454 1662 2457 1668
rect 2470 1652 2473 1658
rect 2458 1648 2462 1651
rect 2392 1603 2394 1607
rect 2398 1603 2401 1607
rect 2405 1603 2408 1607
rect 2282 1558 2286 1561
rect 2322 1558 2326 1561
rect 2362 1548 2366 1551
rect 2238 1522 2241 1528
rect 2270 1482 2273 1538
rect 2278 1502 2281 1528
rect 2294 1492 2297 1548
rect 2374 1532 2377 1548
rect 2318 1512 2321 1518
rect 2342 1492 2345 1528
rect 2382 1502 2385 1598
rect 2406 1542 2409 1578
rect 2414 1562 2417 1568
rect 2446 1532 2449 1548
rect 2454 1542 2457 1648
rect 2510 1592 2513 1668
rect 2574 1652 2577 1658
rect 2590 1652 2593 1668
rect 2614 1662 2617 1668
rect 2622 1652 2625 1658
rect 2522 1648 2526 1651
rect 2646 1642 2649 1648
rect 2502 1542 2505 1568
rect 2478 1492 2481 1508
rect 2534 1502 2537 1618
rect 2542 1572 2545 1628
rect 2694 1612 2697 1658
rect 2702 1642 2705 1658
rect 2742 1642 2745 1659
rect 2626 1588 2630 1591
rect 2738 1568 2742 1571
rect 2582 1542 2585 1548
rect 2278 1482 2281 1488
rect 2490 1478 2494 1481
rect 2302 1472 2305 1478
rect 2366 1472 2369 1478
rect 2510 1472 2513 1478
rect 2474 1468 2478 1471
rect 2218 1459 2222 1462
rect 2074 1378 2078 1381
rect 2114 1358 2118 1361
rect 2014 1342 2017 1348
rect 1958 1312 1961 1328
rect 1966 1322 1969 1338
rect 1934 1298 1945 1301
rect 2046 1302 2049 1358
rect 2142 1352 2145 1398
rect 2174 1392 2177 1408
rect 2222 1392 2225 1398
rect 2278 1392 2281 1458
rect 2286 1442 2289 1468
rect 2306 1448 2310 1451
rect 2302 1392 2305 1438
rect 2334 1392 2337 1448
rect 2438 1432 2441 1448
rect 2454 1442 2457 1468
rect 2486 1462 2489 1468
rect 2494 1462 2497 1468
rect 2462 1452 2465 1458
rect 2518 1452 2521 1498
rect 2526 1488 2534 1491
rect 2526 1472 2529 1488
rect 2574 1472 2577 1518
rect 2590 1491 2593 1558
rect 2750 1552 2753 1728
rect 2766 1722 2769 1748
rect 2774 1742 2777 1848
rect 2798 1752 2801 1878
rect 2830 1872 2833 1918
rect 2838 1892 2841 1948
rect 2846 1902 2849 2038
rect 2870 1992 2873 2068
rect 2878 1942 2881 2068
rect 2982 2062 2985 2068
rect 3006 2062 3009 2078
rect 3078 2072 3081 2108
rect 3174 2102 3177 2118
rect 3202 2078 3206 2081
rect 3094 2072 3097 2078
rect 3102 2072 3105 2078
rect 3134 2072 3137 2078
rect 3074 2068 3078 2071
rect 2894 1992 2897 2038
rect 2946 2018 2950 2021
rect 2886 1952 2889 1958
rect 2854 1932 2857 1940
rect 2862 1922 2865 1938
rect 2866 1868 2870 1871
rect 2826 1858 2830 1861
rect 2838 1852 2841 1868
rect 2830 1848 2838 1851
rect 2830 1792 2833 1848
rect 2822 1742 2825 1748
rect 2846 1742 2849 1868
rect 2854 1862 2857 1868
rect 2854 1822 2857 1858
rect 2870 1852 2873 1858
rect 2878 1842 2881 1928
rect 2904 1903 2906 1907
rect 2910 1903 2913 1907
rect 2917 1903 2920 1907
rect 2926 1882 2929 2008
rect 2990 1942 2993 1948
rect 3022 1942 3025 1947
rect 3030 1942 3033 2068
rect 3066 2058 3070 2061
rect 2942 1932 2945 1938
rect 2934 1922 2937 1928
rect 2958 1912 2961 1918
rect 2958 1892 2961 1898
rect 2998 1892 3001 1918
rect 2910 1872 2913 1878
rect 2886 1868 2905 1871
rect 2886 1862 2889 1868
rect 2902 1862 2905 1868
rect 2918 1862 2921 1868
rect 2870 1792 2873 1818
rect 2894 1762 2897 1858
rect 2862 1752 2865 1758
rect 2862 1742 2865 1748
rect 2874 1738 2878 1741
rect 2758 1662 2761 1718
rect 2774 1712 2777 1738
rect 2854 1732 2857 1738
rect 2918 1722 2921 1748
rect 2926 1742 2929 1878
rect 2962 1868 2966 1871
rect 2990 1862 2993 1868
rect 3030 1862 3033 1938
rect 2938 1858 2942 1861
rect 2970 1858 2974 1861
rect 2958 1762 2961 1848
rect 2990 1792 2993 1848
rect 3022 1792 3025 1818
rect 2990 1772 2993 1788
rect 3030 1781 3033 1858
rect 3022 1778 3033 1781
rect 3046 1781 3049 1858
rect 3054 1792 3057 2018
rect 3078 2002 3081 2058
rect 3094 1932 3097 2068
rect 3158 2062 3161 2068
rect 3106 2058 3110 2061
rect 3138 2058 3142 2061
rect 3174 2052 3177 2078
rect 3234 2068 3238 2071
rect 3218 2058 3222 2061
rect 3130 2048 3134 2051
rect 3110 2032 3113 2038
rect 3102 1942 3105 1998
rect 3150 1992 3153 2028
rect 3118 1942 3121 1948
rect 3086 1922 3089 1928
rect 3094 1872 3097 1928
rect 3046 1778 3057 1781
rect 2938 1758 2942 1761
rect 2994 1758 2998 1761
rect 2934 1742 2937 1748
rect 2942 1742 2945 1758
rect 2926 1732 2929 1738
rect 2946 1728 2950 1731
rect 2794 1718 2798 1721
rect 2846 1692 2849 1708
rect 2810 1688 2814 1691
rect 2878 1672 2881 1708
rect 2904 1703 2906 1707
rect 2910 1703 2913 1707
rect 2917 1703 2920 1707
rect 2958 1692 2961 1758
rect 2970 1748 2974 1751
rect 2982 1732 2985 1758
rect 3014 1752 3017 1768
rect 3006 1742 3009 1748
rect 2974 1692 2977 1698
rect 2982 1692 2985 1718
rect 2774 1662 2777 1668
rect 2814 1662 2817 1668
rect 2942 1662 2945 1668
rect 3022 1662 3025 1778
rect 3030 1762 3033 1768
rect 3046 1752 3049 1768
rect 3038 1742 3041 1748
rect 3054 1702 3057 1778
rect 3062 1742 3065 1858
rect 3094 1752 3097 1868
rect 3102 1852 3105 1938
rect 3114 1888 3118 1891
rect 3126 1872 3129 1958
rect 3142 1952 3145 1968
rect 3158 1952 3161 1998
rect 3134 1872 3137 1948
rect 3114 1868 3118 1871
rect 3134 1852 3137 1868
rect 3142 1862 3145 1928
rect 3158 1892 3161 1948
rect 3174 1942 3177 2038
rect 3170 1938 3174 1941
rect 3182 1932 3185 2048
rect 3190 2002 3193 2058
rect 3246 2052 3249 2138
rect 3286 2112 3289 2128
rect 3326 2122 3329 2138
rect 3254 2062 3257 2078
rect 3318 2062 3321 2068
rect 3290 2058 3294 2061
rect 3210 2048 3214 2051
rect 3298 2048 3302 2051
rect 3326 2042 3329 2098
rect 3342 2081 3345 2118
rect 3350 2102 3353 2128
rect 3334 2078 3345 2081
rect 3374 2081 3377 2118
rect 3382 2092 3385 2148
rect 3406 2142 3409 2148
rect 3478 2142 3481 2218
rect 3494 2212 3497 2258
rect 3646 2252 3649 2268
rect 3566 2172 3569 2248
rect 3614 2202 3617 2218
rect 3570 2168 3574 2171
rect 3602 2148 3606 2151
rect 3622 2142 3625 2228
rect 3654 2192 3657 2448
rect 3726 2442 3729 2448
rect 3694 2362 3697 2378
rect 3726 2362 3729 2408
rect 3734 2392 3737 2458
rect 3758 2452 3761 2458
rect 3742 2432 3745 2438
rect 3750 2362 3753 2418
rect 3758 2372 3761 2448
rect 3766 2382 3769 2458
rect 3810 2448 3814 2451
rect 3806 2392 3809 2428
rect 3830 2392 3833 2518
rect 3870 2462 3873 2568
rect 3890 2548 3894 2551
rect 3914 2548 3918 2551
rect 3878 2532 3881 2538
rect 3886 2512 3889 2528
rect 3902 2492 3905 2548
rect 3910 2532 3913 2538
rect 3942 2532 3945 2558
rect 3958 2522 3961 2588
rect 3982 2572 3985 2578
rect 3990 2562 3993 2568
rect 4014 2562 4017 2568
rect 4046 2562 4049 2618
rect 4070 2602 4073 2648
rect 4102 2572 4105 2658
rect 4118 2652 4121 2678
rect 4142 2672 4145 2678
rect 4154 2668 4158 2671
rect 4126 2662 4129 2668
rect 4162 2658 4166 2661
rect 4182 2651 4185 2738
rect 4206 2692 4209 2748
rect 4278 2742 4281 2748
rect 4298 2747 4302 2750
rect 4506 2748 4510 2751
rect 4378 2738 4382 2741
rect 4230 2732 4233 2738
rect 4266 2718 4270 2721
rect 4366 2712 4369 2728
rect 4278 2682 4281 2698
rect 4194 2678 4198 2681
rect 4174 2648 4185 2651
rect 4174 2642 4177 2648
rect 4174 2572 4177 2638
rect 4182 2592 4185 2618
rect 3928 2503 3930 2507
rect 3934 2503 3937 2507
rect 3941 2503 3944 2507
rect 3858 2458 3862 2461
rect 3870 2452 3873 2458
rect 3878 2452 3881 2478
rect 3918 2462 3921 2468
rect 3934 2462 3937 2468
rect 3890 2458 3894 2461
rect 3910 2452 3913 2458
rect 3886 2442 3889 2448
rect 3942 2442 3945 2478
rect 3950 2462 3953 2518
rect 3958 2462 3961 2518
rect 3974 2482 3977 2528
rect 3982 2522 3985 2558
rect 4014 2552 4017 2558
rect 4022 2552 4025 2558
rect 3982 2492 3985 2508
rect 3990 2502 3993 2548
rect 4030 2522 4033 2558
rect 4054 2542 4057 2548
rect 4038 2522 4041 2528
rect 4062 2522 4065 2548
rect 4130 2547 4134 2550
rect 4078 2538 4086 2541
rect 4006 2498 4014 2501
rect 3974 2472 3977 2478
rect 3998 2462 4001 2488
rect 4006 2472 4009 2498
rect 4014 2482 4017 2488
rect 4022 2471 4025 2518
rect 4046 2472 4049 2518
rect 4062 2502 4065 2518
rect 4022 2468 4030 2471
rect 4034 2458 4038 2461
rect 3998 2452 4001 2458
rect 4046 2452 4049 2458
rect 4006 2442 4009 2448
rect 4054 2441 4057 2458
rect 4078 2452 4081 2538
rect 4086 2492 4089 2518
rect 4094 2512 4097 2528
rect 4158 2522 4161 2548
rect 4190 2532 4193 2648
rect 4214 2642 4217 2668
rect 4222 2652 4225 2658
rect 4230 2652 4233 2678
rect 4238 2662 4241 2678
rect 4262 2672 4265 2678
rect 4286 2672 4289 2678
rect 4302 2672 4305 2688
rect 4350 2672 4353 2688
rect 4366 2682 4369 2708
rect 4374 2672 4377 2718
rect 4414 2692 4417 2748
rect 4430 2732 4433 2748
rect 4462 2742 4465 2748
rect 4494 2742 4497 2748
rect 4390 2679 4398 2681
rect 4390 2678 4401 2679
rect 4382 2672 4385 2678
rect 4334 2662 4337 2668
rect 4238 2652 4241 2658
rect 4262 2652 4265 2658
rect 4302 2652 4305 2658
rect 4326 2652 4329 2658
rect 4358 2652 4361 2668
rect 4390 2662 4393 2678
rect 4430 2672 4433 2688
rect 4454 2672 4457 2718
rect 4462 2662 4465 2738
rect 4486 2732 4489 2738
rect 4526 2732 4529 2758
rect 4534 2742 4537 2748
rect 4542 2732 4545 2748
rect 4578 2738 4582 2741
rect 4614 2732 4617 2768
rect 4630 2762 4633 2768
rect 4662 2752 4665 2818
rect 4678 2772 4681 2848
rect 4710 2832 4713 2848
rect 4742 2842 4745 2848
rect 4862 2842 4865 2848
rect 4694 2782 4697 2818
rect 4710 2762 4713 2768
rect 4718 2762 4721 2778
rect 4726 2762 4729 2818
rect 4742 2762 4745 2838
rect 4758 2832 4761 2838
rect 4738 2748 4742 2751
rect 4622 2742 4625 2748
rect 4694 2742 4697 2748
rect 4750 2741 4753 2818
rect 4758 2752 4761 2828
rect 4746 2738 4753 2741
rect 4782 2741 4785 2818
rect 4798 2752 4801 2818
rect 4846 2742 4849 2748
rect 4778 2738 4785 2741
rect 4810 2738 4814 2741
rect 4826 2738 4830 2741
rect 4638 2732 4641 2738
rect 4478 2712 4481 2728
rect 4486 2701 4489 2728
rect 4478 2698 4489 2701
rect 4478 2692 4481 2698
rect 4486 2688 4494 2691
rect 4486 2672 4489 2688
rect 4574 2678 4577 2718
rect 4598 2682 4601 2718
rect 4614 2692 4617 2728
rect 4686 2722 4689 2738
rect 4750 2732 4753 2738
rect 4798 2732 4801 2738
rect 4862 2732 4865 2758
rect 4878 2742 4881 2768
rect 4894 2762 4897 2818
rect 4894 2751 4897 2758
rect 4890 2748 4897 2751
rect 4926 2752 4929 2758
rect 4926 2742 4929 2748
rect 4898 2738 4902 2741
rect 4818 2728 4822 2731
rect 4758 2722 4761 2728
rect 4790 2722 4793 2728
rect 4622 2692 4625 2718
rect 4646 2682 4649 2718
rect 4670 2702 4673 2718
rect 4642 2678 4646 2681
rect 4594 2668 4598 2671
rect 4650 2668 4654 2671
rect 4506 2658 4510 2661
rect 4282 2648 4286 2651
rect 4250 2638 4254 2641
rect 4198 2552 4201 2628
rect 4198 2542 4201 2548
rect 4190 2512 4193 2518
rect 4238 2492 4241 2618
rect 4262 2592 4265 2648
rect 4338 2638 4342 2641
rect 4414 2622 4417 2648
rect 4462 2622 4465 2658
rect 4534 2632 4537 2668
rect 4542 2662 4545 2668
rect 4614 2652 4617 2668
rect 4622 2662 4625 2668
rect 4610 2648 4614 2651
rect 4574 2642 4577 2648
rect 4686 2642 4689 2658
rect 4702 2652 4705 2668
rect 4710 2661 4713 2718
rect 4726 2682 4729 2718
rect 4750 2702 4753 2718
rect 4782 2702 4785 2718
rect 4790 2672 4793 2688
rect 4738 2668 4742 2671
rect 4718 2662 4721 2668
rect 4710 2658 4718 2661
rect 4798 2652 4801 2728
rect 4814 2722 4817 2728
rect 4870 2722 4873 2728
rect 4822 2712 4825 2718
rect 4814 2662 4817 2688
rect 4822 2672 4825 2678
rect 4846 2651 4849 2698
rect 4854 2682 4857 2718
rect 4894 2711 4897 2728
rect 4922 2718 4926 2721
rect 4886 2708 4897 2711
rect 4878 2672 4881 2678
rect 4878 2652 4881 2668
rect 4846 2648 4854 2651
rect 4710 2642 4713 2648
rect 4862 2642 4865 2648
rect 4730 2638 4734 2641
rect 4646 2632 4649 2638
rect 4334 2592 4337 2618
rect 4534 2612 4537 2628
rect 4440 2603 4442 2607
rect 4446 2603 4449 2607
rect 4453 2603 4456 2607
rect 4478 2572 4481 2578
rect 4426 2568 4430 2571
rect 4466 2568 4470 2571
rect 4498 2568 4502 2571
rect 4390 2562 4393 2568
rect 4622 2562 4625 2568
rect 4418 2558 4422 2561
rect 4562 2558 4566 2561
rect 4586 2558 4590 2561
rect 4406 2552 4409 2558
rect 4366 2542 4369 2548
rect 4422 2542 4425 2548
rect 4478 2542 4481 2548
rect 4386 2538 4390 2541
rect 4402 2538 4406 2541
rect 4246 2532 4249 2538
rect 4302 2521 4305 2538
rect 4302 2518 4310 2521
rect 4102 2488 4110 2491
rect 4094 2472 4097 2488
rect 4102 2472 4105 2488
rect 4234 2478 4238 2481
rect 4246 2472 4249 2518
rect 4270 2472 4273 2478
rect 4186 2468 4190 2471
rect 4218 2468 4222 2471
rect 4082 2448 4086 2451
rect 4046 2438 4057 2441
rect 4066 2438 4070 2441
rect 3662 2342 3665 2348
rect 3678 2342 3681 2348
rect 3710 2342 3713 2348
rect 3774 2342 3777 2358
rect 3782 2352 3785 2358
rect 3798 2352 3801 2388
rect 3822 2352 3825 2358
rect 3754 2338 3758 2341
rect 3786 2338 3790 2341
rect 3670 2272 3673 2278
rect 3662 2262 3665 2268
rect 3678 2262 3681 2328
rect 3718 2271 3721 2338
rect 3710 2268 3721 2271
rect 3694 2232 3697 2248
rect 3710 2242 3713 2268
rect 3718 2252 3721 2258
rect 3726 2252 3729 2308
rect 3734 2282 3737 2318
rect 3750 2312 3753 2338
rect 3830 2332 3833 2378
rect 3854 2342 3857 2348
rect 3870 2332 3873 2348
rect 3886 2332 3889 2418
rect 3934 2412 3937 2418
rect 3942 2382 3945 2438
rect 3914 2358 3918 2361
rect 3930 2358 3934 2361
rect 3898 2340 3902 2343
rect 3910 2342 3913 2358
rect 3874 2328 3878 2331
rect 3758 2322 3761 2328
rect 3770 2318 3774 2321
rect 3878 2302 3881 2318
rect 3882 2288 3886 2291
rect 3734 2272 3737 2278
rect 3742 2262 3745 2288
rect 3766 2282 3769 2288
rect 3854 2282 3857 2288
rect 3894 2282 3897 2340
rect 3950 2341 3953 2378
rect 3962 2368 3966 2371
rect 3974 2362 3977 2408
rect 4046 2392 4049 2438
rect 4054 2382 4057 2418
rect 4002 2368 4006 2371
rect 4058 2368 4062 2371
rect 3970 2348 3974 2351
rect 3946 2338 3953 2341
rect 3982 2342 3985 2348
rect 3998 2342 4001 2348
rect 4006 2341 4009 2358
rect 4030 2342 4033 2368
rect 4070 2362 4073 2378
rect 4094 2362 4097 2458
rect 4118 2452 4121 2458
rect 4134 2382 4137 2388
rect 4106 2368 4110 2371
rect 4078 2352 4081 2358
rect 4042 2348 4046 2351
rect 4066 2348 4070 2351
rect 4118 2342 4121 2358
rect 4006 2338 4014 2341
rect 4014 2332 4017 2338
rect 4078 2332 4081 2338
rect 4126 2332 4129 2368
rect 4142 2342 4145 2428
rect 4150 2422 4153 2468
rect 4238 2462 4241 2468
rect 4218 2458 4222 2461
rect 4174 2452 4177 2458
rect 4206 2452 4209 2458
rect 4158 2392 4161 2448
rect 4190 2432 4193 2448
rect 4222 2442 4225 2448
rect 4206 2432 4209 2438
rect 4166 2352 4169 2418
rect 4174 2412 4177 2418
rect 4246 2372 4249 2468
rect 4246 2358 4254 2361
rect 4166 2342 4169 2348
rect 4142 2332 4145 2338
rect 3910 2312 3913 2318
rect 3928 2303 3930 2307
rect 3934 2303 3937 2307
rect 3941 2303 3944 2307
rect 3882 2278 3886 2281
rect 3670 2142 3673 2168
rect 3678 2152 3681 2218
rect 3694 2192 3697 2218
rect 3718 2202 3721 2218
rect 3742 2192 3745 2208
rect 3750 2142 3753 2258
rect 3758 2252 3761 2278
rect 3794 2268 3798 2271
rect 3766 2262 3769 2268
rect 3782 2252 3785 2268
rect 3790 2242 3793 2258
rect 3802 2248 3806 2251
rect 3814 2242 3817 2268
rect 3854 2262 3857 2268
rect 3842 2258 3846 2261
rect 3842 2228 3846 2231
rect 3830 2152 3833 2218
rect 3846 2172 3849 2228
rect 3870 2222 3873 2278
rect 3898 2268 3902 2271
rect 3902 2242 3905 2258
rect 3910 2162 3913 2218
rect 3918 2152 3921 2278
rect 3926 2272 3929 2288
rect 3938 2278 3942 2281
rect 3934 2272 3937 2278
rect 3926 2242 3929 2268
rect 3946 2248 3950 2251
rect 3930 2158 3934 2161
rect 3802 2148 3806 2151
rect 3902 2142 3905 2148
rect 3958 2142 3961 2318
rect 4022 2292 4025 2318
rect 4182 2292 4185 2348
rect 4206 2342 4209 2348
rect 4198 2312 4201 2328
rect 4246 2292 4249 2358
rect 4262 2352 4265 2458
rect 4270 2451 4273 2468
rect 4310 2462 4313 2468
rect 4278 2452 4281 2458
rect 4270 2448 4278 2451
rect 4270 2372 4273 2448
rect 4326 2392 4329 2459
rect 4350 2402 4353 2538
rect 4390 2512 4393 2538
rect 4494 2532 4497 2558
rect 4530 2548 4542 2551
rect 4562 2548 4566 2551
rect 4578 2548 4582 2551
rect 4510 2532 4513 2548
rect 4526 2542 4529 2548
rect 4622 2542 4625 2548
rect 4402 2468 4406 2471
rect 4422 2452 4425 2478
rect 4430 2472 4433 2518
rect 4534 2512 4537 2538
rect 4590 2532 4593 2538
rect 4558 2512 4561 2528
rect 4630 2512 4633 2548
rect 4638 2501 4641 2618
rect 4630 2498 4641 2501
rect 4486 2472 4489 2478
rect 4466 2468 4470 2471
rect 4394 2448 4398 2451
rect 4458 2448 4462 2451
rect 4482 2448 4486 2451
rect 4494 2451 4497 2478
rect 4510 2472 4513 2478
rect 4534 2462 4537 2468
rect 4490 2448 4497 2451
rect 4510 2452 4513 2458
rect 4522 2448 4526 2451
rect 4274 2358 4278 2361
rect 4306 2358 4310 2361
rect 4310 2348 4326 2351
rect 4302 2342 4305 2348
rect 4270 2332 4273 2338
rect 3966 2242 3969 2288
rect 4134 2282 4137 2288
rect 3990 2272 3993 2278
rect 4078 2272 4081 2278
rect 4110 2272 4113 2278
rect 4166 2272 4169 2278
rect 4010 2268 4014 2271
rect 4098 2268 4102 2271
rect 3974 2242 3977 2258
rect 3982 2252 3985 2268
rect 4030 2262 4033 2268
rect 4050 2258 4054 2261
rect 4090 2258 4094 2261
rect 4106 2258 4110 2261
rect 4130 2258 4134 2261
rect 4014 2252 4017 2258
rect 4050 2248 4054 2251
rect 3990 2182 3993 2248
rect 4022 2232 4025 2238
rect 4030 2222 4033 2238
rect 3982 2152 3985 2158
rect 3990 2152 3993 2168
rect 3998 2142 4001 2198
rect 4062 2192 4065 2228
rect 4026 2158 4030 2161
rect 3850 2138 3854 2141
rect 3374 2078 3385 2081
rect 3202 2038 3206 2041
rect 3218 2038 3222 2041
rect 3258 2038 3262 2041
rect 3286 2022 3289 2038
rect 3294 2032 3297 2038
rect 3254 1962 3257 2018
rect 3310 1962 3313 2018
rect 3218 1948 3222 1951
rect 3198 1942 3201 1948
rect 3214 1932 3217 1938
rect 3190 1922 3193 1928
rect 3230 1922 3233 1938
rect 3214 1892 3217 1908
rect 3238 1882 3241 1958
rect 3246 1931 3249 1948
rect 3254 1942 3257 1958
rect 3262 1942 3265 1948
rect 3286 1932 3289 1958
rect 3310 1952 3313 1958
rect 3318 1942 3321 1968
rect 3334 1961 3337 2078
rect 3358 2072 3361 2078
rect 3346 2068 3350 2071
rect 3366 2062 3369 2068
rect 3374 2062 3377 2068
rect 3342 2052 3345 2058
rect 3358 2052 3361 2058
rect 3358 2032 3361 2048
rect 3366 2042 3369 2058
rect 3366 1992 3369 2028
rect 3326 1958 3337 1961
rect 3354 1958 3358 1961
rect 3326 1942 3329 1958
rect 3370 1948 3374 1951
rect 3334 1942 3337 1948
rect 3358 1942 3361 1948
rect 3382 1942 3385 2078
rect 3390 2072 3393 2078
rect 3398 1952 3401 2048
rect 3406 2032 3409 2138
rect 3450 2118 3454 2121
rect 3414 2062 3417 2098
rect 3422 2082 3425 2118
rect 3486 2112 3489 2138
rect 3534 2121 3537 2138
rect 3530 2118 3537 2121
rect 3558 2102 3561 2135
rect 3694 2102 3697 2132
rect 3502 2092 3505 2098
rect 3726 2092 3729 2138
rect 3650 2088 3654 2091
rect 3714 2088 3718 2091
rect 3494 2078 3513 2081
rect 3422 2072 3425 2078
rect 3494 2072 3497 2078
rect 3434 2068 3438 2071
rect 3510 2071 3513 2078
rect 3754 2078 3758 2081
rect 3566 2072 3569 2078
rect 3622 2072 3625 2078
rect 3630 2072 3633 2078
rect 3798 2072 3801 2138
rect 3826 2128 3830 2131
rect 3850 2128 3854 2131
rect 3838 2122 3841 2128
rect 3870 2112 3873 2118
rect 3910 2092 3913 2138
rect 4030 2132 4033 2138
rect 4018 2128 4022 2131
rect 4006 2122 4009 2128
rect 4038 2122 4041 2158
rect 4062 2142 4065 2168
rect 4078 2132 4081 2158
rect 4094 2142 4097 2168
rect 4102 2162 4105 2248
rect 4150 2192 4153 2258
rect 4090 2128 4094 2131
rect 4142 2122 4145 2128
rect 3928 2103 3930 2107
rect 3934 2103 3937 2107
rect 3941 2103 3944 2107
rect 3822 2072 3825 2078
rect 3510 2068 3518 2071
rect 3802 2068 3806 2071
rect 3438 2062 3441 2068
rect 3442 2048 3446 2051
rect 3414 2032 3417 2038
rect 3416 2003 3418 2007
rect 3422 2003 3425 2007
rect 3429 2003 3432 2007
rect 3406 1962 3409 1968
rect 3454 1952 3457 2028
rect 3462 2022 3465 2068
rect 3470 2052 3473 2068
rect 3502 2062 3505 2068
rect 3574 2062 3577 2068
rect 3554 2058 3558 2061
rect 3478 2022 3481 2058
rect 3590 2052 3593 2058
rect 3534 2032 3537 2038
rect 3534 1972 3537 2028
rect 3542 2022 3545 2048
rect 3558 2042 3561 2048
rect 3606 1992 3609 2048
rect 3506 1948 3510 1951
rect 3298 1938 3302 1941
rect 3246 1928 3254 1931
rect 3282 1928 3286 1931
rect 3350 1892 3353 1918
rect 3390 1892 3393 1918
rect 3398 1912 3401 1928
rect 3478 1892 3481 1928
rect 3486 1922 3489 1938
rect 3534 1932 3537 1938
rect 3514 1918 3518 1921
rect 3542 1912 3545 1938
rect 3566 1922 3569 1932
rect 3578 1918 3582 1921
rect 3486 1892 3489 1908
rect 3598 1892 3601 1918
rect 3606 1892 3609 1988
rect 3654 1952 3657 2018
rect 3678 1992 3681 2068
rect 3686 2032 3689 2068
rect 3734 2042 3737 2068
rect 3838 2052 3841 2059
rect 3750 2022 3753 2028
rect 3750 1992 3753 1998
rect 3902 1952 3905 1958
rect 3934 1952 3937 2018
rect 3746 1948 3750 1951
rect 3158 1862 3161 1868
rect 3106 1848 3110 1851
rect 3154 1848 3158 1851
rect 3166 1851 3169 1878
rect 3254 1872 3257 1878
rect 3162 1848 3169 1851
rect 3194 1868 3198 1871
rect 3134 1822 3137 1848
rect 3174 1822 3177 1868
rect 3198 1852 3201 1858
rect 3214 1852 3217 1858
rect 3210 1848 3214 1851
rect 3190 1782 3193 1818
rect 3270 1792 3273 1808
rect 3166 1742 3169 1758
rect 3110 1722 3113 1738
rect 3078 1712 3081 1718
rect 3078 1692 3081 1698
rect 3046 1663 3049 1678
rect 2910 1652 2913 1659
rect 2790 1592 2793 1608
rect 2674 1548 2678 1551
rect 2606 1542 2609 1548
rect 2702 1542 2705 1548
rect 2766 1542 2769 1568
rect 2918 1552 2921 1618
rect 2822 1542 2825 1548
rect 2718 1532 2721 1538
rect 2582 1488 2593 1491
rect 2610 1488 2614 1491
rect 2582 1472 2585 1488
rect 2630 1452 2633 1468
rect 2654 1462 2657 1488
rect 2670 1482 2673 1488
rect 2714 1478 2718 1481
rect 2706 1468 2710 1471
rect 2758 1462 2761 1468
rect 2774 1462 2777 1538
rect 2830 1521 2833 1538
rect 2878 1532 2881 1538
rect 2918 1522 2921 1548
rect 2974 1542 2977 1588
rect 2998 1562 3001 1568
rect 3078 1552 3081 1658
rect 3094 1612 3097 1658
rect 3086 1552 3089 1558
rect 3034 1548 3038 1551
rect 3034 1538 3038 1541
rect 2830 1518 2838 1521
rect 2846 1502 2849 1518
rect 2904 1503 2906 1507
rect 2910 1503 2913 1507
rect 2917 1503 2920 1507
rect 2926 1492 2929 1538
rect 2982 1522 2985 1538
rect 2954 1518 2958 1521
rect 2898 1488 2902 1491
rect 2862 1472 2865 1478
rect 2926 1472 2929 1478
rect 2974 1472 2977 1498
rect 3006 1492 3009 1518
rect 2998 1472 3001 1478
rect 3014 1472 3017 1478
rect 3022 1472 3025 1478
rect 3042 1468 3046 1471
rect 3086 1462 3089 1488
rect 3094 1462 3097 1608
rect 2690 1448 2694 1451
rect 2714 1448 2718 1451
rect 2746 1448 2750 1451
rect 2650 1438 2654 1441
rect 2638 1432 2641 1438
rect 2530 1418 2537 1421
rect 2546 1418 2550 1421
rect 2234 1378 2238 1381
rect 2246 1372 2249 1378
rect 2342 1372 2345 1378
rect 2246 1362 2249 1368
rect 2382 1362 2385 1418
rect 2392 1403 2394 1407
rect 2398 1403 2401 1407
rect 2405 1403 2408 1407
rect 2534 1392 2537 1418
rect 2194 1358 2198 1361
rect 2266 1358 2270 1361
rect 2322 1358 2326 1361
rect 2178 1348 2182 1351
rect 2194 1348 2198 1351
rect 2250 1348 2254 1351
rect 2106 1338 2110 1341
rect 1934 1282 1937 1298
rect 1942 1272 1945 1288
rect 2054 1282 2057 1338
rect 2086 1281 2089 1332
rect 2118 1282 2121 1338
rect 2126 1292 2129 1328
rect 2086 1278 2094 1281
rect 1862 1261 1865 1268
rect 1838 1258 1849 1261
rect 1854 1258 1865 1261
rect 1874 1258 1878 1261
rect 1822 1252 1825 1258
rect 1762 1248 1766 1251
rect 1758 1192 1761 1228
rect 1782 1192 1785 1248
rect 1838 1192 1841 1258
rect 1854 1192 1857 1258
rect 1894 1212 1897 1268
rect 2002 1259 2006 1262
rect 1902 1182 1905 1258
rect 1910 1192 1913 1258
rect 1670 1152 1673 1158
rect 1706 1148 1710 1151
rect 1666 1138 1670 1141
rect 1654 1112 1657 1118
rect 1662 1092 1665 1128
rect 1686 1122 1689 1138
rect 1726 1121 1729 1148
rect 1774 1142 1777 1148
rect 1726 1118 1734 1121
rect 1694 1102 1697 1118
rect 1658 1088 1662 1091
rect 1622 1082 1625 1088
rect 1630 1082 1633 1088
rect 1742 1082 1745 1132
rect 1782 1092 1785 1178
rect 1830 1162 1833 1168
rect 1902 1162 1905 1168
rect 1926 1162 1929 1218
rect 1958 1192 1961 1208
rect 2022 1192 2025 1268
rect 2054 1262 2057 1268
rect 2070 1262 2073 1278
rect 2110 1272 2113 1278
rect 2134 1272 2137 1348
rect 2214 1342 2217 1348
rect 2286 1342 2289 1358
rect 2350 1352 2353 1358
rect 2398 1352 2401 1358
rect 2410 1348 2414 1351
rect 2234 1338 2238 1341
rect 2142 1272 2145 1338
rect 2162 1328 2166 1331
rect 2190 1328 2198 1331
rect 2266 1328 2270 1331
rect 2182 1292 2185 1328
rect 2154 1278 2158 1281
rect 2178 1278 2182 1281
rect 2190 1272 2193 1328
rect 2286 1282 2289 1338
rect 2310 1322 2313 1338
rect 2318 1332 2321 1348
rect 2422 1342 2425 1348
rect 2470 1342 2473 1378
rect 2662 1362 2665 1448
rect 2846 1442 2849 1459
rect 2958 1452 2961 1459
rect 2994 1458 2998 1461
rect 3034 1458 3038 1461
rect 3102 1452 3105 1668
rect 3118 1622 3121 1738
rect 3138 1718 3142 1721
rect 3182 1672 3185 1768
rect 3190 1762 3193 1778
rect 3238 1732 3241 1747
rect 3254 1742 3257 1748
rect 3254 1682 3257 1738
rect 3286 1692 3289 1859
rect 3302 1752 3305 1868
rect 3326 1842 3329 1888
rect 3342 1878 3350 1881
rect 3334 1872 3337 1878
rect 3342 1862 3345 1878
rect 3354 1858 3358 1861
rect 3334 1852 3337 1858
rect 3342 1852 3345 1858
rect 3366 1852 3369 1878
rect 3406 1872 3409 1888
rect 3426 1868 3430 1871
rect 3394 1858 3398 1861
rect 3398 1842 3401 1848
rect 3302 1742 3305 1748
rect 3334 1742 3337 1747
rect 3390 1712 3393 1747
rect 3406 1742 3409 1858
rect 3442 1848 3446 1851
rect 3416 1803 3418 1807
rect 3422 1803 3425 1807
rect 3429 1803 3432 1807
rect 3502 1752 3505 1868
rect 3566 1862 3569 1868
rect 3622 1862 3625 1928
rect 3630 1922 3633 1948
rect 3694 1942 3697 1948
rect 3742 1932 3745 1938
rect 3690 1918 3694 1921
rect 3686 1872 3689 1878
rect 3702 1872 3705 1918
rect 3790 1912 3793 1948
rect 3874 1947 3878 1950
rect 3742 1892 3745 1908
rect 3928 1903 3930 1907
rect 3934 1903 3937 1907
rect 3941 1903 3944 1907
rect 3950 1902 3953 1948
rect 3842 1888 3846 1891
rect 3550 1792 3553 1858
rect 3494 1742 3497 1748
rect 3518 1742 3521 1748
rect 3534 1742 3537 1748
rect 3558 1742 3561 1748
rect 3566 1742 3569 1748
rect 3590 1742 3593 1748
rect 3462 1732 3465 1738
rect 3482 1728 3486 1731
rect 3458 1718 3462 1721
rect 3342 1692 3345 1708
rect 3334 1682 3337 1688
rect 3374 1682 3377 1688
rect 3318 1672 3321 1678
rect 3306 1668 3310 1671
rect 3134 1662 3137 1668
rect 3250 1659 3254 1662
rect 3134 1592 3137 1658
rect 3190 1642 3193 1648
rect 3150 1572 3153 1618
rect 3254 1592 3257 1608
rect 3294 1562 3297 1668
rect 3302 1652 3305 1658
rect 3318 1642 3321 1658
rect 3134 1552 3137 1558
rect 3190 1551 3193 1558
rect 3150 1544 3153 1548
rect 3258 1548 3262 1551
rect 3110 1462 3113 1498
rect 3150 1491 3153 1540
rect 3146 1488 3153 1491
rect 3158 1492 3161 1538
rect 3222 1502 3225 1548
rect 3266 1538 3270 1541
rect 3230 1492 3233 1508
rect 3246 1492 3249 1538
rect 3278 1492 3281 1518
rect 3194 1478 3198 1481
rect 3182 1471 3185 1478
rect 3182 1468 3193 1471
rect 3210 1468 3214 1471
rect 3242 1468 3246 1471
rect 3046 1442 3049 1448
rect 3158 1442 3161 1448
rect 2678 1412 2681 1418
rect 2726 1402 2729 1418
rect 2790 1392 2793 1438
rect 2682 1378 2686 1381
rect 2550 1342 2553 1348
rect 2606 1342 2609 1358
rect 2530 1338 2534 1341
rect 2714 1338 2718 1341
rect 2374 1332 2377 1338
rect 2390 1332 2393 1338
rect 2294 1292 2297 1308
rect 2306 1278 2310 1281
rect 2198 1272 2201 1278
rect 2082 1268 2086 1271
rect 2098 1268 2102 1271
rect 2130 1268 2134 1271
rect 2250 1268 2254 1271
rect 2290 1268 2294 1271
rect 2042 1258 2046 1261
rect 2086 1252 2089 1258
rect 2042 1248 2046 1251
rect 2070 1162 2073 1178
rect 1802 1158 1806 1161
rect 1850 1158 1854 1161
rect 1798 1132 1801 1138
rect 1814 1132 1817 1138
rect 1790 1122 1793 1128
rect 1830 1122 1833 1158
rect 1842 1148 1846 1151
rect 1866 1138 1870 1141
rect 1886 1132 1889 1158
rect 1814 1092 1817 1118
rect 1872 1103 1874 1107
rect 1878 1103 1881 1107
rect 1885 1103 1888 1107
rect 1902 1092 1905 1158
rect 1990 1152 1993 1158
rect 2054 1152 2057 1158
rect 2086 1152 2089 1228
rect 2094 1162 2097 1168
rect 1942 1142 1945 1148
rect 1914 1138 1918 1141
rect 1970 1138 1974 1141
rect 1934 1132 1937 1138
rect 1950 1112 1953 1138
rect 1982 1132 1985 1148
rect 2038 1142 2041 1148
rect 2094 1142 2097 1158
rect 2110 1152 2113 1268
rect 2134 1192 2137 1248
rect 2138 1148 2142 1151
rect 2050 1138 2054 1141
rect 2106 1138 2110 1141
rect 2130 1138 2134 1141
rect 1958 1122 1961 1128
rect 1990 1082 1993 1138
rect 2006 1092 2009 1135
rect 1970 1078 1974 1081
rect 1758 1072 1761 1078
rect 1846 1072 1849 1078
rect 1810 1068 1814 1071
rect 1850 1068 1854 1071
rect 1494 1018 1505 1021
rect 1494 992 1497 1008
rect 1494 952 1497 958
rect 1474 928 1478 931
rect 1414 872 1417 878
rect 1422 872 1425 918
rect 1454 872 1457 918
rect 1486 892 1489 918
rect 1502 881 1505 1018
rect 1590 992 1593 998
rect 1534 982 1537 988
rect 1598 981 1601 1028
rect 1590 978 1601 981
rect 1542 962 1545 968
rect 1530 958 1534 961
rect 1566 952 1569 968
rect 1510 932 1513 938
rect 1550 892 1553 948
rect 1566 932 1569 948
rect 1582 932 1585 938
rect 1502 878 1510 881
rect 1346 868 1350 871
rect 1502 862 1505 868
rect 1510 862 1513 878
rect 1534 872 1537 888
rect 1542 868 1550 871
rect 1294 852 1297 858
rect 1382 852 1385 858
rect 1134 842 1137 848
rect 1302 842 1305 848
rect 1342 842 1345 848
rect 1346 838 1353 841
rect 1330 828 1334 831
rect 1094 792 1097 818
rect 1142 792 1145 798
rect 1166 792 1169 828
rect 1254 822 1257 828
rect 1122 768 1126 771
rect 1170 768 1174 771
rect 1010 748 1014 751
rect 1050 748 1054 751
rect 1030 732 1033 738
rect 1086 732 1089 738
rect 982 662 985 718
rect 990 672 993 728
rect 1022 702 1025 728
rect 1094 692 1097 748
rect 1118 732 1121 758
rect 1150 752 1153 768
rect 1186 758 1190 761
rect 1230 752 1233 808
rect 1310 802 1313 818
rect 1342 762 1345 768
rect 1314 758 1321 761
rect 1186 748 1193 751
rect 1262 751 1265 758
rect 1142 742 1145 748
rect 1174 742 1177 748
rect 1182 732 1185 738
rect 1006 662 1009 678
rect 1022 672 1025 678
rect 1030 672 1033 688
rect 1078 672 1081 688
rect 1134 682 1137 698
rect 1166 692 1169 698
rect 1190 692 1193 748
rect 1310 742 1313 748
rect 1298 738 1302 741
rect 1318 732 1321 758
rect 1350 752 1353 838
rect 1430 822 1433 858
rect 1368 803 1370 807
rect 1374 803 1377 807
rect 1381 803 1384 807
rect 1358 742 1361 798
rect 1430 792 1433 798
rect 1410 758 1414 761
rect 1438 752 1441 828
rect 1446 802 1449 848
rect 1454 772 1457 858
rect 1542 852 1545 868
rect 1558 852 1561 928
rect 1590 892 1593 978
rect 1606 932 1609 958
rect 1614 942 1617 1058
rect 1622 932 1625 948
rect 1610 928 1614 931
rect 1622 921 1625 928
rect 1614 918 1625 921
rect 1614 892 1617 918
rect 1606 862 1609 868
rect 1630 862 1633 948
rect 1654 922 1657 1058
rect 1726 1052 1729 1059
rect 1742 1042 1745 1068
rect 1830 1062 1833 1068
rect 1838 1052 1841 1068
rect 1878 1062 1881 1078
rect 1942 1072 1945 1078
rect 1926 1062 1929 1068
rect 2014 1062 2017 1108
rect 2038 1062 2041 1128
rect 2110 1092 2113 1118
rect 1846 1052 1849 1058
rect 1942 1052 1945 1058
rect 1966 1052 1969 1058
rect 1906 1048 1910 1051
rect 2038 1042 2041 1058
rect 1714 988 1718 991
rect 1702 962 1705 978
rect 1718 962 1721 968
rect 1750 962 1753 978
rect 1758 972 1761 978
rect 1690 958 1694 961
rect 1690 948 1694 951
rect 1706 948 1710 951
rect 1734 942 1737 948
rect 1782 942 1785 948
rect 1838 942 1841 958
rect 1846 952 1849 958
rect 2022 951 2025 958
rect 2054 952 2057 1088
rect 2070 1062 2073 1088
rect 2126 1072 2129 1098
rect 2142 1092 2145 1138
rect 1670 932 1673 938
rect 1758 932 1761 938
rect 1638 872 1641 918
rect 1662 912 1665 928
rect 1726 892 1729 898
rect 1690 888 1697 891
rect 1694 872 1697 888
rect 1734 878 1737 908
rect 1774 902 1777 938
rect 1790 932 1793 938
rect 1818 918 1822 921
rect 1846 902 1849 948
rect 1886 942 1889 948
rect 1934 942 1937 948
rect 1866 938 1870 941
rect 2054 932 2057 938
rect 2078 932 2081 1068
rect 2134 1062 2137 1078
rect 2142 1072 2145 1078
rect 2102 992 2105 1008
rect 2122 958 2126 961
rect 2142 952 2145 958
rect 2098 948 2102 951
rect 2118 942 2121 948
rect 2134 942 2137 948
rect 2098 938 2102 941
rect 2150 932 2153 1158
rect 2158 1132 2161 1268
rect 2166 1182 2169 1218
rect 2174 1152 2177 1238
rect 2190 1172 2193 1268
rect 2198 1162 2201 1268
rect 2302 1262 2305 1268
rect 2310 1262 2313 1268
rect 2274 1258 2278 1261
rect 2214 1242 2217 1248
rect 2254 1242 2257 1258
rect 2206 1152 2209 1158
rect 2230 1152 2233 1158
rect 2254 1151 2257 1238
rect 2286 1192 2289 1198
rect 2310 1192 2313 1258
rect 2266 1158 2270 1161
rect 2254 1148 2265 1151
rect 2174 1142 2177 1148
rect 2182 1142 2185 1148
rect 2158 1102 2161 1128
rect 2190 1112 2193 1128
rect 2246 1122 2249 1138
rect 2166 1092 2169 1108
rect 2174 1072 2177 1078
rect 2190 1072 2193 1078
rect 2198 1072 2201 1118
rect 2214 1082 2217 1118
rect 2214 1061 2217 1078
rect 2254 1062 2257 1118
rect 2262 1112 2265 1148
rect 2270 1142 2273 1148
rect 2302 1082 2305 1098
rect 2294 1072 2297 1078
rect 2310 1062 2313 1068
rect 2210 1058 2217 1061
rect 2234 1058 2238 1061
rect 2170 1048 2174 1051
rect 2278 1042 2281 1048
rect 2266 1038 2270 1041
rect 1918 912 1921 918
rect 1872 903 1874 907
rect 1878 903 1881 907
rect 1885 903 1888 907
rect 1882 888 1886 891
rect 1954 888 1958 891
rect 1902 872 1905 878
rect 1974 872 1977 878
rect 1986 868 1990 871
rect 1630 852 1633 858
rect 1554 848 1558 851
rect 1466 768 1470 771
rect 1506 768 1510 771
rect 1546 768 1550 771
rect 1518 762 1521 768
rect 1526 762 1529 768
rect 1574 762 1577 768
rect 1482 758 1486 761
rect 1450 748 1454 751
rect 1474 748 1478 751
rect 1374 742 1377 748
rect 1330 738 1334 741
rect 1486 741 1489 748
rect 1482 738 1489 741
rect 1366 732 1369 738
rect 1438 732 1441 738
rect 1510 732 1513 758
rect 1542 752 1545 758
rect 1594 748 1598 751
rect 1558 742 1561 748
rect 1546 738 1550 741
rect 1582 732 1585 738
rect 1590 732 1593 738
rect 1598 732 1601 738
rect 1322 728 1326 731
rect 1378 728 1382 731
rect 1410 728 1414 731
rect 1450 728 1454 731
rect 1490 728 1494 731
rect 1206 692 1209 728
rect 1146 688 1150 691
rect 1250 688 1254 691
rect 1042 668 1046 671
rect 914 658 918 661
rect 1050 658 1054 661
rect 902 642 905 648
rect 942 632 945 648
rect 838 618 849 621
rect 818 568 822 571
rect 742 562 745 568
rect 710 552 713 558
rect 718 542 721 548
rect 750 542 753 558
rect 766 542 769 558
rect 774 552 777 568
rect 830 552 833 618
rect 782 542 785 548
rect 714 538 718 541
rect 702 528 710 531
rect 722 528 726 531
rect 754 528 758 531
rect 662 492 665 508
rect 702 492 705 528
rect 766 502 769 538
rect 838 532 841 558
rect 802 528 806 531
rect 790 492 793 498
rect 846 492 849 618
rect 886 602 889 618
rect 902 592 905 618
rect 966 572 969 648
rect 982 642 985 648
rect 990 592 993 658
rect 1022 652 1025 658
rect 1022 602 1025 648
rect 1038 592 1041 598
rect 862 552 865 568
rect 910 552 913 558
rect 870 542 873 548
rect 910 532 913 538
rect 882 528 886 531
rect 898 528 902 531
rect 934 522 937 558
rect 990 552 993 588
rect 958 522 961 528
rect 856 503 858 507
rect 862 503 865 507
rect 869 503 872 507
rect 822 482 825 488
rect 654 392 657 418
rect 670 362 673 478
rect 678 452 681 468
rect 686 452 689 458
rect 710 442 713 468
rect 734 462 737 468
rect 686 392 689 438
rect 718 432 721 458
rect 742 432 745 458
rect 758 442 761 478
rect 798 472 801 478
rect 770 468 774 471
rect 770 458 774 461
rect 790 452 793 468
rect 838 462 841 478
rect 862 462 865 468
rect 802 458 806 461
rect 822 452 825 458
rect 870 452 873 478
rect 830 422 833 448
rect 846 422 849 438
rect 666 358 670 361
rect 710 352 713 358
rect 658 348 662 351
rect 690 348 694 351
rect 702 342 705 348
rect 662 332 665 338
rect 694 332 697 338
rect 718 332 721 368
rect 750 352 753 368
rect 778 358 782 361
rect 726 332 729 348
rect 738 340 742 343
rect 750 342 753 348
rect 798 342 801 358
rect 830 352 833 358
rect 854 352 857 358
rect 886 352 889 498
rect 966 492 969 538
rect 982 532 985 538
rect 1014 532 1017 538
rect 906 458 910 461
rect 926 442 929 468
rect 942 462 945 468
rect 954 458 958 461
rect 954 448 958 451
rect 942 441 945 448
rect 942 438 953 441
rect 910 422 913 438
rect 950 432 953 438
rect 898 418 902 421
rect 950 392 953 428
rect 966 422 969 438
rect 978 418 982 421
rect 926 352 929 368
rect 882 348 886 351
rect 838 342 841 348
rect 982 342 985 378
rect 990 342 993 438
rect 998 432 1001 468
rect 1006 442 1009 478
rect 1014 442 1017 448
rect 1022 392 1025 548
rect 1030 542 1033 558
rect 1030 532 1033 538
rect 1046 462 1049 608
rect 1070 572 1073 648
rect 1094 572 1097 658
rect 1102 622 1105 648
rect 1110 621 1113 678
rect 1118 652 1121 658
rect 1126 642 1129 658
rect 1134 642 1137 678
rect 1150 652 1153 658
rect 1106 618 1113 621
rect 1102 592 1105 608
rect 1126 592 1129 628
rect 1158 562 1161 678
rect 1310 672 1313 678
rect 1318 672 1321 718
rect 1470 692 1473 718
rect 1574 712 1577 718
rect 1606 692 1609 838
rect 1630 792 1633 848
rect 1646 842 1649 868
rect 1766 862 1769 868
rect 1794 858 1798 861
rect 1742 792 1745 828
rect 1830 802 1833 838
rect 1846 792 1849 848
rect 1870 792 1873 838
rect 1690 748 1694 751
rect 1662 742 1665 748
rect 1710 742 1713 788
rect 1718 752 1721 778
rect 1862 772 1865 788
rect 1790 762 1793 768
rect 1814 742 1817 748
rect 1862 742 1865 768
rect 1654 702 1657 738
rect 1686 692 1689 718
rect 1750 692 1753 728
rect 1758 692 1761 738
rect 1806 732 1809 738
rect 1886 722 1889 728
rect 1714 688 1721 691
rect 1366 672 1369 688
rect 1502 672 1505 678
rect 1258 668 1262 671
rect 1170 658 1174 661
rect 1078 542 1081 558
rect 1182 552 1185 648
rect 1198 642 1201 668
rect 1222 652 1225 658
rect 1230 642 1233 668
rect 1238 612 1241 668
rect 1390 662 1393 668
rect 1278 652 1281 658
rect 1422 652 1425 658
rect 1254 572 1257 648
rect 1438 642 1441 668
rect 1230 551 1233 558
rect 1334 552 1337 638
rect 1070 512 1073 528
rect 1086 512 1089 548
rect 1110 502 1113 538
rect 1158 502 1161 538
rect 1166 482 1169 518
rect 1198 511 1201 548
rect 1342 542 1345 598
rect 1350 592 1353 618
rect 1446 612 1449 668
rect 1494 632 1497 668
rect 1566 662 1569 668
rect 1368 603 1370 607
rect 1374 603 1377 607
rect 1381 603 1384 607
rect 1446 592 1449 598
rect 1478 592 1481 628
rect 1406 542 1409 568
rect 1494 562 1497 628
rect 1574 572 1577 618
rect 1606 592 1609 688
rect 1718 672 1721 688
rect 1726 672 1729 678
rect 1774 672 1777 698
rect 1854 692 1857 718
rect 1872 703 1874 707
rect 1878 703 1881 707
rect 1885 703 1888 707
rect 1830 672 1833 678
rect 1894 672 1897 838
rect 1906 758 1910 761
rect 1906 728 1910 731
rect 1918 721 1921 868
rect 1990 858 1998 861
rect 1978 848 1982 851
rect 1926 732 1929 758
rect 1934 742 1937 778
rect 1958 772 1961 778
rect 1950 762 1953 768
rect 1918 718 1929 721
rect 1926 692 1929 718
rect 1966 692 1969 828
rect 1618 668 1622 671
rect 1906 668 1910 671
rect 1634 659 1638 662
rect 1670 641 1673 668
rect 1662 638 1673 641
rect 1802 658 1806 661
rect 1662 592 1665 638
rect 1726 592 1729 598
rect 1662 562 1665 588
rect 1414 542 1417 548
rect 1190 508 1201 511
rect 1470 541 1473 558
rect 1550 552 1553 558
rect 1466 538 1473 541
rect 1486 542 1489 548
rect 1626 538 1630 541
rect 1690 538 1694 541
rect 1190 492 1193 508
rect 1190 472 1193 488
rect 1206 472 1209 478
rect 1078 462 1081 468
rect 1142 462 1145 468
rect 1174 463 1177 468
rect 1070 422 1073 458
rect 1078 352 1081 458
rect 1098 348 1102 351
rect 930 338 934 341
rect 1042 338 1046 341
rect 758 332 761 338
rect 526 262 529 268
rect 574 182 577 218
rect 582 212 585 268
rect 622 192 625 238
rect 430 168 441 171
rect 438 162 441 168
rect 374 142 377 158
rect 398 152 401 158
rect 410 148 414 151
rect 338 138 342 141
rect 174 122 177 128
rect 78 72 81 88
rect 174 82 177 98
rect 110 72 113 79
rect 126 72 129 78
rect 174 72 177 78
rect 230 72 233 128
rect 238 72 241 118
rect 246 102 249 138
rect 102 68 110 71
rect 102 62 105 68
rect 138 66 142 69
rect 162 58 166 61
rect 178 58 182 61
rect 254 61 257 138
rect 382 132 385 148
rect 446 142 449 148
rect 434 128 438 131
rect 262 82 265 88
rect 266 68 270 71
rect 250 58 262 61
rect 94 52 97 58
rect 294 52 297 88
rect 302 82 305 98
rect 422 92 425 118
rect 438 82 441 128
rect 454 92 457 168
rect 470 132 473 168
rect 490 148 494 151
rect 490 138 494 141
rect 502 132 505 158
rect 518 142 521 158
rect 530 148 534 151
rect 542 142 545 168
rect 558 162 561 178
rect 570 168 574 171
rect 590 162 593 168
rect 630 162 633 268
rect 682 258 686 261
rect 654 242 657 258
rect 694 252 697 298
rect 726 282 729 298
rect 714 268 721 271
rect 706 258 710 261
rect 666 248 670 251
rect 718 242 721 268
rect 750 262 753 308
rect 758 282 761 328
rect 766 312 769 318
rect 766 282 769 298
rect 782 242 785 318
rect 806 272 809 338
rect 862 332 865 338
rect 798 242 801 248
rect 642 238 646 241
rect 682 238 686 241
rect 746 238 750 241
rect 726 222 729 228
rect 654 182 657 218
rect 726 192 729 208
rect 750 202 753 218
rect 638 172 641 178
rect 790 172 793 178
rect 702 162 705 168
rect 570 158 574 161
rect 558 152 561 158
rect 582 152 585 158
rect 598 152 601 158
rect 646 152 649 158
rect 706 148 710 151
rect 530 138 534 141
rect 550 141 553 148
rect 550 138 561 141
rect 478 122 481 128
rect 454 82 457 88
rect 462 82 465 118
rect 510 92 513 118
rect 318 72 321 78
rect 366 72 369 78
rect 470 72 473 88
rect 518 82 521 98
rect 542 92 545 138
rect 558 132 561 138
rect 582 132 585 148
rect 602 138 606 141
rect 630 132 633 148
rect 650 138 654 141
rect 558 92 561 128
rect 598 92 601 128
rect 606 88 614 91
rect 550 82 553 88
rect 494 72 497 78
rect 510 72 513 78
rect 550 72 553 78
rect 566 72 569 88
rect 606 72 609 88
rect 654 72 657 88
rect 662 82 665 148
rect 702 138 710 141
rect 790 142 793 168
rect 798 152 801 158
rect 806 152 809 198
rect 814 182 817 328
rect 822 262 825 318
rect 838 302 841 318
rect 856 303 858 307
rect 862 303 865 307
rect 869 303 872 307
rect 1046 302 1049 318
rect 838 252 841 298
rect 862 288 870 291
rect 882 288 886 291
rect 862 272 865 288
rect 982 282 985 288
rect 1078 282 1081 298
rect 1102 292 1105 338
rect 1110 322 1113 418
rect 1174 392 1177 438
rect 1214 392 1217 538
rect 1262 532 1265 538
rect 1310 522 1313 538
rect 1290 518 1294 521
rect 1222 492 1225 518
rect 1342 512 1345 538
rect 1362 518 1366 521
rect 1318 492 1321 508
rect 1406 492 1409 528
rect 1462 522 1465 538
rect 1494 532 1497 538
rect 1258 468 1262 471
rect 1222 462 1225 468
rect 1226 448 1230 451
rect 1246 442 1249 448
rect 1270 442 1273 478
rect 1438 472 1441 488
rect 1350 462 1353 468
rect 1294 452 1297 458
rect 1374 432 1377 468
rect 1422 452 1425 468
rect 1454 463 1457 468
rect 1368 403 1370 407
rect 1374 403 1377 407
rect 1381 403 1384 407
rect 1198 342 1201 388
rect 1390 382 1393 408
rect 1406 392 1409 448
rect 1462 392 1465 498
rect 1526 482 1529 518
rect 1542 492 1545 538
rect 1574 532 1577 538
rect 1590 492 1593 518
rect 1562 478 1566 481
rect 1526 452 1529 478
rect 1614 475 1617 508
rect 1622 492 1625 528
rect 1554 468 1558 471
rect 1590 468 1598 471
rect 1542 462 1545 468
rect 1538 448 1542 451
rect 1502 382 1505 388
rect 1270 352 1273 358
rect 1298 348 1302 351
rect 1358 342 1361 368
rect 1370 348 1374 351
rect 1422 348 1430 351
rect 1422 342 1425 348
rect 1322 338 1326 341
rect 1338 338 1342 341
rect 1142 332 1145 338
rect 1190 322 1193 338
rect 1174 292 1177 318
rect 1198 312 1201 338
rect 1202 288 1206 291
rect 1014 272 1017 278
rect 1038 272 1041 278
rect 822 171 825 218
rect 910 172 913 268
rect 930 258 934 261
rect 954 258 958 261
rect 970 258 974 261
rect 918 242 921 248
rect 938 238 942 241
rect 818 168 825 171
rect 830 162 833 168
rect 894 158 902 161
rect 894 142 897 158
rect 906 148 910 151
rect 926 151 929 218
rect 950 212 953 248
rect 998 232 1001 258
rect 922 148 929 151
rect 958 152 961 218
rect 1014 192 1017 268
rect 1022 262 1025 268
rect 1042 258 1046 261
rect 1030 232 1033 258
rect 918 142 921 148
rect 1022 142 1025 218
rect 1038 172 1041 218
rect 1046 152 1049 198
rect 1054 162 1057 258
rect 1078 212 1081 278
rect 1086 272 1089 278
rect 1134 272 1137 278
rect 1206 272 1209 278
rect 1238 272 1241 298
rect 1254 292 1257 338
rect 1382 332 1385 338
rect 1274 328 1278 331
rect 1430 331 1433 338
rect 1422 328 1433 331
rect 1078 162 1081 198
rect 1086 162 1089 258
rect 1142 241 1145 268
rect 1142 238 1153 241
rect 1094 192 1097 238
rect 1030 142 1033 148
rect 670 132 673 138
rect 678 82 681 98
rect 702 92 705 138
rect 782 132 785 140
rect 842 138 846 141
rect 890 138 894 141
rect 930 138 934 141
rect 822 122 825 138
rect 846 132 849 138
rect 854 122 857 138
rect 942 132 945 138
rect 958 132 961 138
rect 1070 132 1073 138
rect 874 128 881 131
rect 922 128 926 131
rect 1026 128 1030 131
rect 702 82 705 88
rect 306 68 310 71
rect 418 68 422 71
rect 442 68 446 71
rect 486 62 489 68
rect 518 62 521 68
rect 526 62 529 68
rect 386 58 390 61
rect 418 58 422 61
rect 586 58 590 61
rect 626 58 630 61
rect 658 58 662 61
rect 478 52 481 58
rect 566 52 569 58
rect 686 52 689 68
rect 718 62 721 118
rect 734 52 737 58
rect 742 52 745 98
rect 758 72 761 108
rect 766 102 769 118
rect 766 72 769 78
rect 798 72 801 78
rect 786 68 790 71
rect 750 62 753 68
rect 806 62 809 78
rect 790 52 793 58
rect 822 52 825 118
rect 830 92 833 118
rect 856 103 858 107
rect 862 103 865 107
rect 869 103 872 107
rect 846 92 849 98
rect 878 92 881 128
rect 830 82 833 88
rect 902 82 905 118
rect 902 72 905 78
rect 926 62 929 128
rect 942 52 945 88
rect 950 72 953 78
rect 966 62 969 118
rect 990 92 993 128
rect 998 92 1001 118
rect 1038 92 1041 108
rect 1010 78 1014 81
rect 1026 78 1030 81
rect 1054 72 1057 88
rect 1066 78 1070 81
rect 1078 72 1081 158
rect 1102 152 1105 168
rect 1118 162 1121 208
rect 1126 192 1129 198
rect 1150 192 1153 238
rect 1134 152 1137 168
rect 1174 162 1177 228
rect 1190 212 1193 268
rect 1262 262 1265 328
rect 1334 322 1337 328
rect 1242 258 1246 261
rect 1262 252 1265 258
rect 1270 252 1273 318
rect 1302 292 1305 298
rect 1310 272 1313 278
rect 1318 272 1321 308
rect 1282 268 1286 271
rect 1330 268 1334 271
rect 1230 242 1233 248
rect 1250 238 1254 241
rect 1190 152 1193 158
rect 1142 148 1150 151
rect 1094 142 1097 148
rect 1126 142 1129 148
rect 1142 112 1145 148
rect 1214 142 1217 228
rect 1270 192 1273 248
rect 1286 222 1289 258
rect 1306 248 1313 251
rect 1290 147 1294 150
rect 1170 138 1174 141
rect 1290 138 1294 141
rect 1190 132 1193 138
rect 1226 128 1230 131
rect 1166 122 1169 128
rect 1234 118 1238 121
rect 1090 88 1094 91
rect 1130 78 1134 81
rect 1010 68 1014 71
rect 974 52 977 68
rect 990 62 993 68
rect 1042 58 1046 61
rect 982 52 985 58
rect 1094 52 1097 78
rect 1114 68 1118 71
rect 1138 68 1142 71
rect 1150 62 1153 108
rect 1166 62 1169 78
rect 1182 72 1185 118
rect 1222 82 1225 108
rect 1246 72 1249 118
rect 1310 82 1313 248
rect 1326 222 1329 248
rect 1342 242 1345 328
rect 1350 272 1353 328
rect 1414 292 1417 328
rect 1422 292 1425 328
rect 1430 322 1433 328
rect 1438 292 1441 338
rect 1486 332 1489 338
rect 1494 312 1497 338
rect 1510 322 1513 358
rect 1518 352 1521 358
rect 1542 352 1545 378
rect 1550 372 1553 378
rect 1582 362 1585 368
rect 1530 348 1534 351
rect 1566 342 1569 348
rect 1574 342 1577 358
rect 1542 332 1545 338
rect 1582 332 1585 338
rect 1590 322 1593 468
rect 1646 462 1649 532
rect 1654 412 1657 458
rect 1678 432 1681 538
rect 1702 532 1705 558
rect 1694 482 1697 518
rect 1702 472 1705 528
rect 1710 462 1713 538
rect 1734 492 1737 532
rect 1774 512 1777 658
rect 1838 622 1841 668
rect 1894 581 1897 668
rect 1950 602 1953 628
rect 1958 612 1961 668
rect 1894 578 1905 581
rect 1890 568 1894 571
rect 1798 552 1801 568
rect 1814 532 1817 558
rect 1830 542 1833 568
rect 1858 558 1862 561
rect 1842 548 1846 551
rect 1858 548 1862 551
rect 1882 548 1886 551
rect 1774 492 1777 508
rect 1734 482 1737 488
rect 1722 468 1726 471
rect 1698 458 1702 461
rect 1726 452 1729 458
rect 1706 448 1710 451
rect 1742 442 1745 468
rect 1678 382 1681 418
rect 1622 342 1625 378
rect 1682 348 1686 351
rect 1654 342 1657 348
rect 1602 338 1606 341
rect 1666 338 1670 341
rect 1682 338 1686 341
rect 1694 332 1697 398
rect 1702 392 1705 438
rect 1750 382 1753 428
rect 1790 392 1793 518
rect 1798 402 1801 448
rect 1742 372 1745 378
rect 1706 348 1710 351
rect 1702 342 1705 348
rect 1726 342 1729 358
rect 1750 352 1753 378
rect 1790 361 1793 388
rect 1782 358 1793 361
rect 1782 352 1785 358
rect 1762 348 1766 351
rect 1602 328 1606 331
rect 1470 292 1473 308
rect 1518 292 1521 318
rect 1386 278 1390 281
rect 1426 278 1430 281
rect 1534 272 1537 308
rect 1614 302 1617 318
rect 1622 292 1625 318
rect 1630 282 1633 328
rect 1638 322 1641 328
rect 1718 322 1721 328
rect 1734 292 1737 348
rect 1754 338 1758 341
rect 1602 278 1606 281
rect 1546 268 1550 271
rect 1358 222 1361 268
rect 1398 252 1401 268
rect 1326 152 1329 208
rect 1368 203 1370 207
rect 1374 203 1377 207
rect 1381 203 1384 207
rect 1398 192 1401 238
rect 1406 222 1409 258
rect 1446 242 1449 268
rect 1478 262 1481 268
rect 1458 258 1462 261
rect 1462 242 1465 248
rect 1478 192 1481 198
rect 1350 152 1353 178
rect 1390 162 1393 188
rect 1450 158 1457 161
rect 1330 148 1334 151
rect 1390 142 1393 158
rect 1442 138 1446 141
rect 1406 122 1409 138
rect 1414 132 1417 138
rect 1442 128 1446 131
rect 1454 131 1457 158
rect 1462 142 1465 188
rect 1486 162 1489 268
rect 1558 262 1561 268
rect 1566 252 1569 278
rect 1678 272 1681 278
rect 1710 272 1713 288
rect 1742 282 1745 318
rect 1758 312 1761 328
rect 1790 322 1793 348
rect 1806 332 1809 348
rect 1814 342 1817 398
rect 1822 392 1825 468
rect 1838 442 1841 478
rect 1846 472 1849 538
rect 1862 512 1865 528
rect 1872 503 1874 507
rect 1878 503 1881 507
rect 1885 503 1888 507
rect 1874 488 1878 491
rect 1858 468 1862 471
rect 1846 462 1849 468
rect 1882 458 1886 461
rect 1854 422 1857 448
rect 1886 422 1889 448
rect 1830 382 1833 418
rect 1846 372 1849 378
rect 1830 362 1833 368
rect 1862 362 1865 418
rect 1894 392 1897 448
rect 1850 348 1854 351
rect 1890 348 1894 351
rect 1826 338 1830 341
rect 1838 322 1841 338
rect 1886 322 1889 338
rect 1872 303 1874 307
rect 1878 303 1881 307
rect 1885 303 1888 307
rect 1718 278 1737 281
rect 1594 268 1598 271
rect 1574 262 1577 268
rect 1554 238 1558 241
rect 1494 162 1497 218
rect 1526 192 1529 238
rect 1574 231 1577 248
rect 1582 242 1585 268
rect 1606 262 1609 268
rect 1574 228 1585 231
rect 1582 192 1585 228
rect 1470 131 1473 148
rect 1450 128 1457 131
rect 1462 128 1473 131
rect 1450 118 1454 121
rect 1462 92 1465 128
rect 1486 102 1489 158
rect 1494 132 1497 158
rect 1518 142 1521 148
rect 1534 142 1537 168
rect 1542 152 1545 168
rect 1558 162 1561 188
rect 1598 172 1601 218
rect 1614 162 1617 268
rect 1686 262 1689 268
rect 1702 262 1705 268
rect 1718 262 1721 278
rect 1734 271 1737 278
rect 1734 268 1742 271
rect 1658 258 1662 261
rect 1726 252 1729 268
rect 1750 252 1753 278
rect 1774 272 1777 288
rect 1782 282 1785 298
rect 1822 272 1825 288
rect 1902 281 1905 578
rect 1926 562 1929 568
rect 1918 482 1921 548
rect 1926 532 1929 538
rect 1942 532 1945 578
rect 1950 552 1953 598
rect 1958 562 1961 608
rect 1974 572 1977 678
rect 1982 582 1985 618
rect 1990 592 1993 858
rect 2006 852 2009 878
rect 2014 862 2017 868
rect 2022 802 2025 928
rect 2070 922 2073 928
rect 2054 892 2057 898
rect 2094 892 2097 908
rect 2134 892 2137 898
rect 2166 892 2169 978
rect 2190 952 2193 1018
rect 2214 952 2217 1038
rect 2274 1018 2278 1021
rect 2230 972 2233 1018
rect 2274 948 2278 951
rect 2190 892 2193 948
rect 2214 942 2217 948
rect 2262 932 2265 938
rect 2110 872 2113 888
rect 2206 882 2209 898
rect 2214 882 2217 928
rect 2178 878 2182 881
rect 2222 872 2225 878
rect 2230 872 2233 888
rect 2238 872 2241 908
rect 2262 892 2265 918
rect 2294 882 2297 898
rect 2302 892 2305 1048
rect 2318 1002 2321 1328
rect 2382 1312 2385 1328
rect 2478 1321 2481 1338
rect 2546 1328 2550 1331
rect 2478 1318 2486 1321
rect 2570 1318 2574 1321
rect 2462 1308 2470 1311
rect 2326 1272 2329 1278
rect 2334 1252 2337 1298
rect 2342 1262 2345 1308
rect 2342 1222 2345 1258
rect 2366 1192 2369 1288
rect 2390 1262 2393 1268
rect 2406 1252 2409 1259
rect 2454 1242 2457 1248
rect 2392 1203 2394 1207
rect 2398 1203 2401 1207
rect 2405 1203 2408 1207
rect 2462 1192 2465 1308
rect 2474 1288 2478 1291
rect 2418 1178 2422 1181
rect 2326 1142 2329 1168
rect 2342 1152 2345 1158
rect 2446 1152 2449 1168
rect 2470 1162 2473 1178
rect 2478 1172 2481 1218
rect 2494 1192 2497 1268
rect 2438 1142 2441 1148
rect 2398 1122 2401 1138
rect 2454 1132 2457 1138
rect 2478 1122 2481 1148
rect 2486 1142 2489 1168
rect 2502 1162 2505 1318
rect 2590 1262 2593 1308
rect 2598 1302 2601 1338
rect 2654 1322 2657 1338
rect 2662 1332 2665 1338
rect 2626 1318 2630 1321
rect 2630 1292 2633 1298
rect 2690 1288 2694 1291
rect 2674 1268 2678 1271
rect 2614 1262 2617 1268
rect 2526 1242 2529 1258
rect 2558 1252 2561 1259
rect 2518 1192 2521 1218
rect 2638 1192 2641 1248
rect 2662 1212 2665 1268
rect 2670 1252 2673 1258
rect 2610 1158 2614 1161
rect 2502 1132 2505 1138
rect 2326 1092 2329 1118
rect 2326 1022 2329 1048
rect 2334 1041 2337 1118
rect 2350 1072 2353 1078
rect 2366 1072 2369 1098
rect 2382 1092 2385 1108
rect 2454 1092 2457 1118
rect 2558 1082 2561 1158
rect 2566 1092 2569 1158
rect 2622 1152 2625 1158
rect 2574 1102 2577 1148
rect 2634 1138 2638 1141
rect 2650 1138 2654 1141
rect 2590 1092 2593 1138
rect 2606 1082 2609 1128
rect 2614 1092 2617 1138
rect 2634 1128 2638 1131
rect 2622 1082 2625 1128
rect 2670 1122 2673 1138
rect 2638 1092 2641 1118
rect 2362 1068 2366 1071
rect 2490 1068 2494 1071
rect 2438 1062 2441 1068
rect 2526 1062 2529 1068
rect 2542 1062 2545 1078
rect 2346 1058 2350 1061
rect 2506 1058 2510 1061
rect 2334 1038 2342 1041
rect 2318 872 2321 988
rect 2326 962 2329 1018
rect 2350 972 2353 1038
rect 2358 1022 2361 1048
rect 2382 1041 2385 1058
rect 2374 1038 2385 1041
rect 2462 1042 2465 1048
rect 2358 992 2361 1008
rect 2374 992 2377 1038
rect 2392 1003 2394 1007
rect 2398 1003 2401 1007
rect 2405 1003 2408 1007
rect 2478 982 2481 1058
rect 2494 1022 2497 1048
rect 2514 1018 2518 1021
rect 2346 968 2350 971
rect 2378 968 2382 971
rect 2366 962 2369 968
rect 2526 962 2529 1058
rect 2550 1042 2553 1058
rect 2574 1052 2577 1078
rect 2598 1072 2601 1078
rect 2606 1052 2609 1078
rect 2614 1058 2622 1061
rect 2658 1058 2662 1061
rect 2582 1022 2585 1048
rect 2358 942 2361 948
rect 2338 938 2342 941
rect 2358 872 2361 908
rect 2366 902 2369 958
rect 2390 952 2393 958
rect 2414 942 2417 958
rect 2430 942 2433 948
rect 2438 932 2441 958
rect 2462 942 2465 958
rect 2494 952 2497 958
rect 2558 952 2561 958
rect 2538 948 2542 951
rect 2602 948 2606 951
rect 2490 938 2494 941
rect 2522 938 2526 941
rect 2034 868 2038 871
rect 2162 868 2166 871
rect 2178 868 2182 871
rect 2290 868 2294 871
rect 2038 852 2041 858
rect 2054 852 2057 868
rect 2130 858 2134 861
rect 2146 858 2150 861
rect 2050 848 2054 851
rect 2006 752 2009 798
rect 2038 772 2041 828
rect 2094 792 2097 858
rect 2146 848 2150 851
rect 2158 842 2161 868
rect 2214 862 2217 868
rect 2250 858 2254 861
rect 2214 852 2217 858
rect 2138 838 2142 841
rect 2166 792 2169 848
rect 2270 842 2273 868
rect 2290 848 2297 851
rect 2138 768 2142 771
rect 2038 751 2041 768
rect 2082 758 2086 761
rect 2086 742 2089 748
rect 2110 742 2113 758
rect 2182 752 2185 758
rect 2070 732 2073 738
rect 2158 732 2161 738
rect 2206 732 2209 748
rect 2186 728 2190 731
rect 2030 662 2033 688
rect 2038 672 2041 728
rect 2102 692 2105 728
rect 2110 692 2113 728
rect 2150 692 2153 718
rect 2174 702 2177 728
rect 2214 722 2217 738
rect 2078 672 2081 678
rect 2182 672 2185 708
rect 2062 642 2065 668
rect 2006 592 2009 598
rect 2062 552 2065 638
rect 2126 612 2129 668
rect 2134 662 2137 668
rect 1974 542 1977 548
rect 1982 532 1985 538
rect 1942 522 1945 528
rect 1954 527 1958 530
rect 1926 482 1929 498
rect 1934 472 1937 478
rect 1918 432 1921 468
rect 1974 462 1977 468
rect 1982 462 1985 518
rect 1998 502 2001 528
rect 1990 452 1993 478
rect 2006 472 2009 488
rect 2014 482 2017 528
rect 2022 522 2025 528
rect 2058 488 2065 491
rect 2062 472 2065 488
rect 2070 482 2073 558
rect 2086 551 2089 558
rect 2102 492 2105 608
rect 2118 592 2121 598
rect 2174 552 2177 568
rect 2070 472 2073 478
rect 2166 472 2169 538
rect 2182 502 2185 668
rect 2198 642 2201 668
rect 2222 662 2225 808
rect 2270 792 2273 818
rect 2286 792 2289 838
rect 2294 822 2297 848
rect 2310 842 2313 868
rect 2366 862 2369 868
rect 2386 858 2390 861
rect 2406 852 2409 898
rect 2414 862 2417 878
rect 2422 862 2425 918
rect 2430 902 2433 928
rect 2462 922 2465 938
rect 2474 928 2478 931
rect 2486 892 2489 928
rect 2494 882 2497 928
rect 2502 882 2505 898
rect 2446 862 2449 878
rect 2542 872 2545 938
rect 2550 912 2553 928
rect 2574 922 2577 938
rect 2606 922 2609 938
rect 2614 932 2617 1058
rect 2670 1052 2673 1108
rect 2678 1092 2681 1208
rect 2686 1162 2689 1168
rect 2694 1162 2697 1228
rect 2702 1212 2705 1248
rect 2710 1192 2713 1328
rect 2726 1281 2729 1338
rect 2722 1278 2729 1281
rect 2718 1272 2721 1278
rect 2726 1261 2729 1268
rect 2722 1258 2729 1261
rect 2686 1142 2689 1148
rect 2694 1070 2697 1158
rect 2702 1148 2710 1151
rect 2702 1132 2705 1148
rect 2718 1142 2721 1258
rect 2734 1252 2737 1348
rect 2750 1332 2753 1378
rect 2806 1372 2809 1378
rect 2862 1362 2865 1408
rect 2830 1358 2838 1361
rect 2846 1358 2854 1361
rect 2830 1351 2833 1358
rect 2794 1348 2833 1351
rect 2826 1338 2830 1341
rect 2766 1322 2769 1328
rect 2774 1302 2777 1328
rect 2782 1292 2785 1338
rect 2826 1328 2830 1331
rect 2798 1292 2801 1298
rect 2806 1282 2809 1328
rect 2818 1278 2822 1281
rect 2786 1268 2790 1271
rect 2758 1262 2761 1268
rect 2750 1252 2753 1258
rect 2750 1192 2753 1238
rect 2758 1212 2761 1248
rect 2774 1222 2777 1268
rect 2814 1262 2817 1268
rect 2786 1258 2790 1261
rect 2838 1232 2841 1348
rect 2846 1282 2849 1358
rect 2870 1352 2873 1418
rect 2942 1362 2945 1368
rect 2982 1362 2985 1398
rect 2930 1358 2934 1361
rect 2886 1302 2889 1338
rect 2902 1332 2905 1358
rect 2982 1342 2985 1358
rect 2970 1338 2977 1341
rect 2942 1332 2945 1338
rect 2914 1328 2918 1331
rect 2974 1312 2977 1338
rect 2986 1328 2990 1331
rect 2998 1312 3001 1338
rect 3014 1332 3017 1438
rect 3062 1362 3065 1378
rect 3102 1352 3105 1378
rect 3142 1352 3145 1378
rect 3174 1352 3177 1458
rect 3182 1452 3185 1458
rect 3190 1432 3193 1468
rect 3286 1462 3289 1478
rect 3214 1432 3217 1458
rect 3230 1442 3233 1448
rect 3294 1442 3297 1558
rect 3306 1548 3310 1551
rect 3314 1538 3318 1541
rect 3326 1541 3329 1558
rect 3322 1538 3329 1541
rect 3310 1462 3313 1498
rect 3334 1482 3337 1678
rect 3366 1672 3369 1678
rect 3422 1662 3425 1698
rect 3478 1692 3481 1728
rect 3502 1722 3505 1738
rect 3510 1731 3513 1738
rect 3510 1728 3518 1731
rect 3434 1668 3438 1671
rect 3362 1658 3369 1661
rect 3366 1652 3369 1658
rect 3446 1652 3449 1678
rect 3458 1658 3462 1661
rect 3474 1658 3478 1661
rect 3502 1661 3505 1718
rect 3498 1658 3505 1661
rect 3510 1692 3513 1728
rect 3526 1702 3529 1718
rect 3510 1662 3513 1688
rect 3526 1682 3529 1688
rect 3518 1652 3521 1668
rect 3506 1648 3510 1651
rect 3534 1651 3537 1738
rect 3546 1728 3550 1731
rect 3598 1691 3601 1718
rect 3606 1702 3609 1758
rect 3614 1752 3617 1768
rect 3598 1688 3609 1691
rect 3658 1688 3662 1691
rect 3606 1682 3609 1688
rect 3594 1678 3598 1681
rect 3546 1658 3550 1661
rect 3530 1648 3537 1651
rect 3486 1642 3489 1648
rect 3382 1592 3385 1638
rect 3494 1632 3497 1638
rect 3342 1562 3345 1568
rect 3342 1542 3345 1548
rect 3366 1542 3369 1558
rect 3354 1538 3358 1541
rect 3390 1532 3393 1538
rect 3350 1512 3353 1528
rect 3358 1492 3361 1528
rect 3346 1478 3350 1481
rect 3186 1388 3190 1391
rect 3314 1388 3318 1391
rect 3026 1348 3030 1351
rect 3182 1348 3190 1351
rect 3246 1351 3249 1358
rect 3150 1342 3153 1348
rect 3174 1342 3177 1348
rect 3050 1338 3054 1341
rect 3006 1322 3009 1328
rect 3014 1322 3017 1328
rect 2904 1303 2906 1307
rect 2910 1303 2913 1307
rect 2917 1303 2920 1307
rect 2862 1282 2865 1288
rect 2846 1252 2849 1278
rect 2854 1232 2857 1278
rect 2910 1272 2913 1278
rect 2874 1268 2878 1271
rect 2902 1262 2905 1268
rect 2882 1258 2886 1261
rect 2886 1242 2889 1248
rect 2738 1168 2742 1171
rect 2714 1138 2718 1141
rect 2718 1092 2721 1128
rect 2726 1122 2729 1158
rect 2734 1142 2737 1148
rect 2774 1142 2777 1208
rect 2782 1152 2785 1218
rect 2902 1192 2905 1258
rect 2942 1242 2945 1258
rect 2950 1252 2953 1258
rect 2958 1252 2961 1278
rect 2966 1262 2969 1268
rect 2974 1252 2977 1308
rect 2982 1272 2985 1278
rect 3054 1272 3057 1318
rect 3038 1262 3041 1268
rect 3002 1258 3006 1261
rect 3022 1252 3025 1258
rect 3046 1252 3049 1258
rect 3062 1252 3065 1338
rect 3094 1332 3097 1338
rect 3118 1332 3121 1338
rect 3102 1282 3105 1288
rect 3070 1262 3073 1268
rect 3094 1262 3097 1278
rect 3110 1261 3113 1318
rect 3126 1272 3129 1318
rect 3154 1268 3158 1271
rect 3110 1258 3118 1261
rect 3158 1252 3161 1258
rect 2970 1248 2974 1251
rect 2918 1212 2921 1218
rect 2822 1152 2825 1158
rect 2762 1138 2766 1141
rect 2902 1141 2905 1168
rect 2954 1158 2958 1161
rect 2898 1138 2905 1141
rect 2754 1128 2758 1131
rect 2822 1102 2825 1135
rect 2838 1112 2841 1138
rect 2846 1102 2849 1138
rect 2862 1092 2865 1118
rect 2870 1112 2873 1118
rect 2894 1082 2897 1138
rect 2934 1132 2937 1138
rect 2914 1128 2918 1131
rect 2904 1103 2906 1107
rect 2910 1103 2913 1107
rect 2917 1103 2920 1107
rect 2742 1072 2745 1078
rect 2690 1066 2694 1069
rect 2730 1068 2734 1071
rect 2702 1052 2705 1068
rect 2742 1052 2745 1058
rect 2706 1048 2710 1051
rect 2650 1038 2654 1041
rect 2662 1032 2665 1048
rect 2734 992 2737 1048
rect 2750 1042 2753 1058
rect 2766 1042 2769 1048
rect 2774 1042 2777 1078
rect 2782 1062 2785 1068
rect 2790 1022 2793 1048
rect 2798 1042 2801 1048
rect 2806 1042 2809 1078
rect 2854 1072 2857 1078
rect 2886 1072 2889 1078
rect 2814 1062 2817 1068
rect 2926 1062 2929 1078
rect 2834 1058 2838 1061
rect 2850 1058 2854 1061
rect 2882 1058 2886 1061
rect 2914 1058 2918 1061
rect 2834 1048 2838 1051
rect 2810 1038 2814 1041
rect 2742 992 2745 998
rect 2854 992 2857 1048
rect 2862 1022 2865 1048
rect 2862 992 2865 1018
rect 2874 968 2878 971
rect 2650 948 2654 951
rect 2678 951 2681 958
rect 2798 952 2801 968
rect 2710 942 2713 948
rect 2822 942 2825 948
rect 2758 932 2761 938
rect 2622 922 2625 928
rect 2550 882 2553 908
rect 2558 882 2561 918
rect 2582 912 2585 918
rect 2614 902 2617 918
rect 2582 882 2585 898
rect 2646 882 2649 888
rect 2570 878 2574 881
rect 2498 868 2502 871
rect 2518 862 2521 868
rect 2558 862 2561 878
rect 2638 872 2641 878
rect 2726 872 2729 888
rect 2742 872 2745 908
rect 2774 892 2777 938
rect 2870 922 2873 928
rect 2858 918 2862 921
rect 2830 882 2833 888
rect 2586 868 2590 871
rect 2794 868 2801 871
rect 2826 868 2830 871
rect 2566 862 2569 868
rect 2710 863 2713 868
rect 2466 858 2470 861
rect 2438 852 2441 858
rect 2526 852 2529 858
rect 2790 852 2793 858
rect 2330 848 2334 851
rect 2422 842 2425 848
rect 2454 842 2457 848
rect 2414 832 2417 838
rect 2618 818 2622 821
rect 2358 792 2361 818
rect 2392 803 2394 807
rect 2398 803 2401 807
rect 2405 803 2408 807
rect 2498 778 2502 781
rect 2294 772 2297 778
rect 2766 771 2769 828
rect 2774 782 2777 818
rect 2798 792 2801 868
rect 2814 842 2817 858
rect 2886 792 2889 1048
rect 2934 1042 2937 1128
rect 2942 1072 2945 1148
rect 2950 1070 2953 1158
rect 2966 1142 2969 1168
rect 2966 1101 2969 1138
rect 2974 1132 2977 1138
rect 2982 1122 2985 1248
rect 3030 1242 3033 1248
rect 3062 1242 3065 1248
rect 3006 1232 3009 1238
rect 2998 1222 3001 1228
rect 3054 1222 3057 1228
rect 3006 1192 3009 1208
rect 3102 1192 3105 1238
rect 3182 1202 3185 1348
rect 3194 1328 3198 1331
rect 3230 1282 3233 1328
rect 3230 1263 3233 1278
rect 3246 1272 3249 1328
rect 3262 1282 3265 1288
rect 3246 1262 3249 1268
rect 3294 1262 3297 1268
rect 2990 1162 2993 1178
rect 2990 1142 2993 1158
rect 2998 1132 3001 1168
rect 3198 1162 3201 1188
rect 3198 1152 3201 1158
rect 3294 1152 3297 1258
rect 2958 1098 2969 1101
rect 2958 1072 2961 1098
rect 2966 1082 2969 1088
rect 2950 1062 2953 1066
rect 2958 951 2961 978
rect 2990 962 2993 968
rect 2974 942 2977 948
rect 2904 903 2906 907
rect 2910 903 2913 907
rect 2917 903 2920 907
rect 2966 892 2969 908
rect 2998 892 3001 1118
rect 3046 1072 3049 1138
rect 3062 1122 3065 1148
rect 3134 1142 3137 1148
rect 3062 1079 3070 1081
rect 3062 1078 3073 1079
rect 2894 863 2897 888
rect 3006 882 3009 928
rect 3022 912 3025 1058
rect 3046 942 3049 1068
rect 3062 1062 3065 1078
rect 3086 1072 3089 1138
rect 3102 952 3105 1038
rect 3142 992 3145 1148
rect 3150 1072 3153 1078
rect 3158 1062 3161 1068
rect 3166 1042 3169 1058
rect 3182 1052 3185 1088
rect 3214 1072 3217 1118
rect 3294 1072 3297 1148
rect 3310 1092 3313 1118
rect 3310 1082 3313 1088
rect 3318 1071 3321 1258
rect 3310 1068 3321 1071
rect 3326 1152 3329 1448
rect 3346 1438 3350 1441
rect 3366 1422 3369 1458
rect 3382 1442 3385 1478
rect 3390 1462 3393 1488
rect 3398 1452 3401 1608
rect 3406 1572 3409 1608
rect 3416 1603 3418 1607
rect 3422 1603 3425 1607
rect 3429 1603 3432 1607
rect 3422 1552 3425 1558
rect 3414 1542 3417 1548
rect 3462 1542 3465 1558
rect 3418 1518 3425 1521
rect 3414 1492 3417 1508
rect 3422 1482 3425 1518
rect 3406 1462 3409 1468
rect 3342 1272 3345 1328
rect 3358 1272 3361 1348
rect 3366 1272 3369 1318
rect 3390 1282 3393 1418
rect 3406 1332 3409 1458
rect 3450 1438 3454 1441
rect 3462 1432 3465 1518
rect 3478 1462 3481 1468
rect 3494 1462 3497 1488
rect 3502 1472 3505 1508
rect 3470 1432 3473 1438
rect 3486 1431 3489 1448
rect 3494 1432 3497 1458
rect 3486 1428 3494 1431
rect 3416 1403 3418 1407
rect 3422 1403 3425 1407
rect 3429 1403 3432 1407
rect 3478 1361 3481 1418
rect 3510 1402 3513 1648
rect 3558 1642 3561 1668
rect 3578 1658 3582 1661
rect 3566 1652 3569 1658
rect 3590 1652 3593 1658
rect 3614 1652 3617 1678
rect 3662 1672 3665 1678
rect 3634 1668 3638 1671
rect 3630 1658 3638 1661
rect 3630 1652 3633 1658
rect 3582 1642 3585 1648
rect 3566 1592 3569 1628
rect 3522 1548 3526 1551
rect 3550 1502 3553 1538
rect 3598 1501 3601 1618
rect 3670 1602 3673 1859
rect 3686 1791 3689 1868
rect 3718 1862 3721 1868
rect 3774 1863 3777 1888
rect 3934 1882 3937 1888
rect 3806 1862 3809 1868
rect 3854 1862 3857 1868
rect 3718 1842 3721 1848
rect 3686 1788 3697 1791
rect 3678 1722 3681 1747
rect 3694 1742 3697 1788
rect 3726 1752 3729 1858
rect 3742 1762 3745 1858
rect 3870 1822 3873 1859
rect 3714 1748 3718 1751
rect 3694 1692 3697 1708
rect 3710 1692 3713 1698
rect 3718 1692 3721 1738
rect 3730 1718 3734 1721
rect 3742 1672 3745 1758
rect 3758 1752 3761 1758
rect 3754 1748 3758 1751
rect 3762 1738 3766 1741
rect 3774 1741 3777 1758
rect 3770 1738 3777 1741
rect 3782 1742 3785 1748
rect 3790 1742 3793 1758
rect 3894 1751 3897 1758
rect 3862 1742 3865 1748
rect 3902 1742 3905 1858
rect 3810 1738 3814 1741
rect 3966 1741 3969 2068
rect 3982 2042 3985 2118
rect 4006 2102 4009 2118
rect 4018 2088 4022 2091
rect 4054 2082 4057 2118
rect 3994 2078 4001 2081
rect 4058 2078 4062 2081
rect 3998 2072 4001 2078
rect 4070 2072 4073 2098
rect 4058 2068 4062 2071
rect 4102 2071 4105 2078
rect 4110 2071 4113 2118
rect 4102 2068 4113 2071
rect 3990 2062 3993 2068
rect 4006 1962 4009 1968
rect 3974 1952 3977 1958
rect 4022 1942 4025 1968
rect 4042 1958 4046 1961
rect 4030 1942 4033 1948
rect 4046 1942 4049 1948
rect 3974 1932 3977 1938
rect 4054 1932 4057 1958
rect 4062 1942 4065 1948
rect 3982 1882 3985 1898
rect 4070 1892 4073 1988
rect 4078 1962 4081 1968
rect 4086 1962 4089 2058
rect 4094 2052 4097 2058
rect 4102 2052 4105 2068
rect 4142 2062 4145 2078
rect 4114 2058 4118 2061
rect 4138 2048 4142 2051
rect 4106 2038 4110 2041
rect 4110 1952 4113 2018
rect 4118 1992 4121 2018
rect 4150 1982 4153 2148
rect 4158 2112 4161 2268
rect 4214 2242 4217 2268
rect 4222 2262 4225 2268
rect 4270 2252 4273 2268
rect 4186 2218 4190 2221
rect 4222 2182 4225 2248
rect 4278 2232 4281 2338
rect 4310 2331 4313 2348
rect 4334 2342 4337 2368
rect 4306 2328 4313 2331
rect 4350 2332 4353 2358
rect 4286 2312 4289 2328
rect 4310 2292 4313 2318
rect 4326 2272 4329 2278
rect 4334 2272 4337 2288
rect 4342 2272 4345 2278
rect 4310 2262 4313 2268
rect 4298 2258 4302 2261
rect 4334 2252 4337 2268
rect 4290 2238 4294 2241
rect 4282 2228 4289 2231
rect 4254 2202 4257 2218
rect 4270 2192 4273 2208
rect 4226 2178 4230 2181
rect 4238 2172 4241 2178
rect 4250 2168 4254 2171
rect 4214 2162 4217 2168
rect 4262 2162 4265 2178
rect 4278 2172 4281 2178
rect 4226 2158 4230 2161
rect 4242 2148 4246 2151
rect 4274 2148 4278 2151
rect 4206 2092 4209 2128
rect 4286 2092 4289 2228
rect 4294 2222 4297 2228
rect 4302 2222 4305 2248
rect 4310 2242 4313 2248
rect 4294 2162 4297 2188
rect 4342 2172 4345 2258
rect 4350 2242 4353 2288
rect 4358 2241 4361 2448
rect 4542 2442 4545 2488
rect 4586 2478 4590 2481
rect 4602 2478 4606 2481
rect 4630 2472 4633 2498
rect 4638 2482 4641 2488
rect 4586 2468 4590 2471
rect 4610 2468 4614 2471
rect 4570 2458 4574 2461
rect 4594 2458 4598 2461
rect 4630 2452 4633 2458
rect 4638 2452 4641 2458
rect 4558 2442 4561 2448
rect 4530 2438 4534 2441
rect 4394 2418 4398 2421
rect 4440 2403 4442 2407
rect 4446 2403 4449 2407
rect 4453 2403 4456 2407
rect 4542 2372 4545 2378
rect 4530 2368 4534 2371
rect 4366 2352 4369 2358
rect 4398 2352 4401 2358
rect 4422 2342 4425 2348
rect 4470 2342 4473 2358
rect 4494 2342 4497 2368
rect 4446 2322 4449 2338
rect 4474 2328 4478 2331
rect 4502 2322 4505 2348
rect 4510 2332 4513 2358
rect 4518 2322 4521 2348
rect 4550 2332 4553 2418
rect 4574 2362 4577 2418
rect 4586 2358 4590 2361
rect 4590 2342 4593 2348
rect 4654 2342 4657 2588
rect 4662 2572 4665 2578
rect 4670 2572 4673 2578
rect 4678 2562 4681 2628
rect 4670 2552 4673 2558
rect 4686 2542 4689 2548
rect 4682 2538 4686 2541
rect 4702 2532 4705 2558
rect 4710 2552 4713 2558
rect 4718 2542 4721 2618
rect 4734 2542 4737 2638
rect 4758 2592 4761 2618
rect 4798 2552 4801 2598
rect 4790 2542 4793 2548
rect 4702 2502 4705 2518
rect 4726 2482 4729 2518
rect 4734 2512 4737 2528
rect 4662 2472 4665 2478
rect 4670 2472 4673 2478
rect 4678 2461 4681 2468
rect 4674 2458 4681 2461
rect 4694 2462 4697 2478
rect 4734 2462 4737 2508
rect 4742 2472 4745 2528
rect 4770 2518 4774 2521
rect 4766 2482 4769 2488
rect 4790 2482 4793 2498
rect 4782 2472 4785 2478
rect 4798 2472 4801 2548
rect 4814 2542 4817 2618
rect 4846 2572 4849 2598
rect 4830 2552 4833 2558
rect 4862 2552 4865 2558
rect 4870 2552 4873 2618
rect 4886 2612 4889 2708
rect 4934 2692 4937 2858
rect 4982 2852 4985 2868
rect 4990 2862 4993 2878
rect 5014 2862 5017 2878
rect 5038 2872 5041 2878
rect 5022 2852 5025 2868
rect 5062 2862 5065 2868
rect 5110 2862 5113 2928
rect 5126 2922 5129 2948
rect 5118 2862 5121 2918
rect 4942 2832 4945 2848
rect 4950 2842 4953 2848
rect 4998 2842 5001 2848
rect 5046 2842 5049 2848
rect 4990 2772 4993 2818
rect 5010 2748 5014 2751
rect 5026 2748 5030 2751
rect 4966 2742 4969 2748
rect 4942 2732 4945 2738
rect 4974 2722 4977 2738
rect 5022 2732 5025 2738
rect 5002 2728 5006 2731
rect 4952 2703 4954 2707
rect 4958 2703 4961 2707
rect 4965 2703 4968 2707
rect 4914 2668 4918 2671
rect 4894 2652 4897 2658
rect 4898 2638 4902 2641
rect 4898 2618 4902 2621
rect 4910 2592 4913 2648
rect 4982 2602 4985 2718
rect 4990 2672 4993 2728
rect 5006 2702 5009 2718
rect 4998 2652 5001 2658
rect 4990 2632 4993 2648
rect 5006 2642 5009 2688
rect 5022 2642 5025 2648
rect 5030 2642 5033 2718
rect 5038 2692 5041 2818
rect 5046 2692 5049 2718
rect 5038 2662 5041 2678
rect 5054 2672 5057 2718
rect 5070 2682 5073 2738
rect 5046 2652 5049 2668
rect 5070 2662 5073 2678
rect 5086 2652 5089 2758
rect 5098 2748 5102 2751
rect 5110 2742 5113 2858
rect 5142 2801 5145 2948
rect 5206 2942 5209 3058
rect 5182 2932 5185 2938
rect 5174 2872 5177 2888
rect 5206 2862 5209 2938
rect 5246 2911 5249 3078
rect 5254 3062 5257 3088
rect 5262 3082 5265 3128
rect 5270 3072 5273 3078
rect 5278 3062 5281 3148
rect 5274 3048 5278 3051
rect 5286 3032 5289 3058
rect 5294 3022 5297 3038
rect 5262 2932 5265 3018
rect 5286 2952 5289 3018
rect 5294 2942 5297 2948
rect 5266 2928 5270 2931
rect 5258 2918 5262 2921
rect 5246 2908 5257 2911
rect 5222 2862 5225 2868
rect 5142 2798 5153 2801
rect 5150 2792 5153 2798
rect 5206 2742 5209 2858
rect 5222 2832 5225 2858
rect 5214 2751 5217 2758
rect 5134 2662 5137 2698
rect 5142 2672 5145 2688
rect 5182 2672 5185 2678
rect 5074 2648 5078 2651
rect 5094 2642 5097 2658
rect 5182 2652 5185 2668
rect 5194 2658 5198 2661
rect 5122 2648 5126 2651
rect 5190 2642 5193 2648
rect 5058 2638 5062 2641
rect 5106 2638 5110 2641
rect 5134 2632 5137 2638
rect 5158 2632 5161 2638
rect 5230 2632 5233 2908
rect 5254 2742 5257 2908
rect 5270 2862 5273 2918
rect 5278 2772 5281 2918
rect 5286 2912 5289 2938
rect 5302 2902 5305 3118
rect 5310 3052 5313 3068
rect 5310 2952 5313 2968
rect 5302 2861 5305 2879
rect 5302 2858 5310 2861
rect 5286 2842 5289 2848
rect 5274 2758 5278 2761
rect 5302 2752 5305 2858
rect 5262 2711 5265 2748
rect 5278 2712 5281 2728
rect 5262 2708 5278 2711
rect 4998 2572 5001 2618
rect 4886 2552 4889 2568
rect 4842 2548 4846 2551
rect 4806 2502 4809 2538
rect 4822 2532 4825 2538
rect 4814 2492 4817 2518
rect 4814 2472 4817 2478
rect 4766 2462 4769 2468
rect 4838 2462 4841 2538
rect 4870 2532 4873 2548
rect 4894 2542 4897 2558
rect 4934 2552 4937 2558
rect 4934 2542 4937 2548
rect 4942 2542 4945 2568
rect 4982 2562 4985 2568
rect 5094 2562 5097 2618
rect 5238 2612 5241 2658
rect 5018 2558 5022 2561
rect 4966 2542 4969 2558
rect 4990 2542 4993 2548
rect 5014 2542 5017 2548
rect 4914 2528 4929 2531
rect 4926 2522 4929 2528
rect 4978 2518 4982 2521
rect 4854 2482 4857 2488
rect 4870 2472 4873 2518
rect 4878 2492 4881 2508
rect 4754 2458 4758 2461
rect 4826 2458 4830 2461
rect 4886 2452 4889 2468
rect 4894 2452 4897 2478
rect 4910 2472 4913 2488
rect 4918 2472 4921 2518
rect 4952 2503 4954 2507
rect 4958 2503 4961 2507
rect 4965 2503 4968 2507
rect 4942 2482 4945 2498
rect 4990 2478 4993 2538
rect 5022 2532 5025 2538
rect 4934 2472 4937 2478
rect 5022 2472 5025 2508
rect 5038 2482 5041 2518
rect 5070 2502 5073 2538
rect 5078 2482 5081 2518
rect 5094 2502 5097 2538
rect 5102 2532 5105 2578
rect 5138 2568 5142 2571
rect 5182 2542 5185 2548
rect 5198 2542 5201 2568
rect 5254 2542 5257 2548
rect 5102 2522 5105 2528
rect 5102 2512 5105 2518
rect 5094 2472 5097 2498
rect 5110 2492 5113 2538
rect 5158 2532 5161 2538
rect 5246 2532 5249 2538
rect 5262 2532 5265 2688
rect 5270 2662 5273 2708
rect 5270 2642 5273 2648
rect 5270 2532 5273 2608
rect 4962 2468 4966 2471
rect 5026 2458 5030 2461
rect 5038 2452 5041 2468
rect 5126 2462 5129 2468
rect 5058 2458 5062 2461
rect 5090 2458 5094 2461
rect 5102 2452 5105 2458
rect 5142 2452 5145 2478
rect 5158 2472 5161 2478
rect 5154 2458 5158 2461
rect 4722 2448 4726 2451
rect 5074 2448 5078 2451
rect 5154 2448 5158 2451
rect 4750 2442 4753 2448
rect 4686 2392 4689 2418
rect 4754 2378 4758 2381
rect 4670 2342 4673 2378
rect 4730 2368 4734 2371
rect 4754 2368 4758 2371
rect 4766 2362 4769 2378
rect 4826 2358 4830 2361
rect 4734 2352 4737 2358
rect 4714 2348 4721 2351
rect 4562 2338 4566 2341
rect 4574 2332 4577 2338
rect 4466 2318 4470 2321
rect 4530 2318 4534 2321
rect 4366 2252 4369 2288
rect 4398 2282 4401 2318
rect 4470 2272 4473 2278
rect 4486 2272 4489 2318
rect 4526 2292 4529 2318
rect 4566 2312 4569 2328
rect 4598 2321 4601 2338
rect 4678 2332 4681 2348
rect 4718 2342 4721 2348
rect 4742 2332 4745 2358
rect 4766 2352 4769 2358
rect 4790 2332 4793 2358
rect 4862 2352 4865 2358
rect 4894 2352 4897 2448
rect 5058 2438 5062 2441
rect 5082 2438 5086 2441
rect 5114 2438 5118 2441
rect 4910 2382 4913 2438
rect 5094 2432 5097 2438
rect 4910 2352 4913 2378
rect 4918 2372 4921 2418
rect 4954 2368 4958 2371
rect 4818 2348 4822 2351
rect 4882 2348 4886 2351
rect 4798 2342 4801 2348
rect 4846 2342 4849 2348
rect 4918 2342 4921 2368
rect 4982 2342 4985 2348
rect 4826 2338 4830 2341
rect 4906 2338 4910 2341
rect 4598 2318 4606 2321
rect 4542 2292 4545 2308
rect 4590 2302 4593 2318
rect 4570 2288 4574 2291
rect 4534 2272 4537 2278
rect 4434 2268 4438 2271
rect 4514 2268 4521 2271
rect 4374 2262 4377 2268
rect 4422 2262 4425 2268
rect 4486 2262 4489 2268
rect 4402 2258 4406 2261
rect 4506 2258 4510 2261
rect 4414 2252 4417 2258
rect 4518 2251 4521 2268
rect 4514 2248 4521 2251
rect 4446 2242 4449 2248
rect 4358 2238 4369 2241
rect 4386 2238 4390 2241
rect 4366 2192 4369 2238
rect 4398 2232 4401 2238
rect 4310 2162 4313 2168
rect 4298 2158 4302 2161
rect 4294 2142 4297 2148
rect 4334 2142 4337 2158
rect 4410 2148 4414 2151
rect 4310 2112 4313 2138
rect 4334 2102 4337 2138
rect 4342 2112 4345 2128
rect 4350 2122 4353 2138
rect 4414 2122 4417 2138
rect 4422 2082 4425 2198
rect 4430 2192 4433 2218
rect 4440 2203 4442 2207
rect 4446 2203 4449 2207
rect 4453 2203 4456 2207
rect 4502 2172 4505 2248
rect 4526 2232 4529 2268
rect 4550 2262 4553 2278
rect 4558 2232 4561 2278
rect 4614 2272 4617 2308
rect 4638 2282 4641 2288
rect 4654 2282 4657 2328
rect 4686 2322 4689 2328
rect 4662 2272 4665 2318
rect 4694 2292 4697 2318
rect 4814 2292 4817 2338
rect 4894 2322 4897 2338
rect 4938 2328 4942 2331
rect 4834 2318 4838 2321
rect 4910 2312 4913 2328
rect 4942 2318 4950 2321
rect 4694 2281 4697 2288
rect 4694 2278 4702 2281
rect 4738 2278 4742 2281
rect 4686 2272 4689 2278
rect 4758 2272 4761 2278
rect 4566 2268 4574 2271
rect 4674 2268 4678 2271
rect 4738 2268 4742 2271
rect 4566 2262 4569 2268
rect 4638 2262 4641 2268
rect 4718 2262 4721 2268
rect 4574 2252 4577 2258
rect 4590 2252 4593 2258
rect 4574 2192 4577 2248
rect 4598 2232 4601 2248
rect 4606 2242 4609 2258
rect 4622 2232 4625 2258
rect 4766 2252 4769 2268
rect 4774 2262 4777 2288
rect 4854 2272 4857 2278
rect 4910 2272 4913 2278
rect 4942 2272 4945 2318
rect 4952 2303 4954 2307
rect 4958 2303 4961 2307
rect 4965 2303 4968 2307
rect 4990 2302 4993 2418
rect 5026 2368 5030 2371
rect 5014 2362 5017 2368
rect 5046 2362 5049 2398
rect 5054 2362 5057 2418
rect 5062 2382 5065 2418
rect 5102 2372 5105 2378
rect 5074 2368 5078 2371
rect 5002 2358 5006 2361
rect 5058 2358 5062 2361
rect 4998 2342 5001 2358
rect 5086 2352 5089 2358
rect 5042 2348 5046 2351
rect 5098 2348 5102 2351
rect 5018 2338 5022 2341
rect 5006 2281 5009 2318
rect 5062 2312 5065 2348
rect 5070 2342 5073 2348
rect 5094 2332 5097 2338
rect 5022 2282 5025 2288
rect 5006 2278 5014 2281
rect 4982 2272 4985 2278
rect 4962 2268 4966 2271
rect 4798 2262 4801 2268
rect 4846 2262 4849 2268
rect 4902 2262 4905 2268
rect 4922 2258 4926 2261
rect 4930 2258 4934 2261
rect 4886 2252 4889 2258
rect 4942 2252 4945 2268
rect 5006 2262 5009 2278
rect 5046 2272 5049 2288
rect 5086 2272 5089 2298
rect 5110 2292 5113 2418
rect 5134 2402 5137 2448
rect 5118 2342 5121 2348
rect 5126 2302 5129 2368
rect 5134 2312 5137 2348
rect 5150 2332 5153 2358
rect 5166 2322 5169 2518
rect 5190 2512 5193 2528
rect 5270 2522 5273 2528
rect 5174 2462 5177 2508
rect 5182 2472 5185 2478
rect 5206 2462 5209 2508
rect 5214 2502 5217 2518
rect 5262 2512 5265 2518
rect 5214 2472 5217 2478
rect 5238 2462 5241 2508
rect 5270 2492 5273 2508
rect 5246 2479 5254 2481
rect 5246 2478 5257 2479
rect 5246 2462 5249 2478
rect 5190 2452 5193 2458
rect 5206 2412 5209 2418
rect 5182 2392 5185 2398
rect 5214 2382 5217 2388
rect 5194 2358 5198 2361
rect 5182 2342 5185 2348
rect 5190 2332 5193 2338
rect 5166 2292 5169 2298
rect 5146 2278 5150 2281
rect 5174 2272 5177 2308
rect 5198 2282 5201 2358
rect 5214 2342 5217 2348
rect 5214 2292 5217 2338
rect 5222 2332 5225 2338
rect 5230 2331 5233 2348
rect 5254 2331 5257 2348
rect 5278 2342 5281 2698
rect 5294 2672 5297 2678
rect 5286 2662 5289 2668
rect 5302 2662 5305 2738
rect 5290 2658 5297 2661
rect 5286 2562 5289 2618
rect 5286 2542 5289 2548
rect 5294 2522 5297 2658
rect 5294 2482 5297 2498
rect 5302 2482 5305 2518
rect 5286 2462 5289 2468
rect 5290 2348 5294 2351
rect 5310 2342 5313 2538
rect 5230 2328 5238 2331
rect 5254 2328 5262 2331
rect 5278 2291 5281 2318
rect 5270 2288 5281 2291
rect 5206 2282 5209 2288
rect 5246 2272 5249 2278
rect 5058 2268 5062 2271
rect 5226 2268 5230 2271
rect 4994 2258 4998 2261
rect 4754 2248 4758 2251
rect 5002 2248 5006 2251
rect 4734 2202 4737 2218
rect 4594 2168 4598 2171
rect 4626 2168 4630 2171
rect 4550 2162 4553 2168
rect 4442 2148 4446 2151
rect 4526 2142 4529 2148
rect 4434 2128 4438 2131
rect 4462 2091 4465 2138
rect 4470 2132 4473 2138
rect 4542 2122 4545 2158
rect 4550 2142 4553 2148
rect 4566 2142 4569 2158
rect 4582 2152 4585 2168
rect 4590 2152 4593 2158
rect 4594 2148 4598 2151
rect 4606 2142 4609 2148
rect 4614 2142 4617 2148
rect 4638 2142 4641 2188
rect 4654 2162 4657 2178
rect 4662 2162 4665 2168
rect 4678 2142 4681 2178
rect 4714 2148 4718 2151
rect 4650 2138 4654 2141
rect 4682 2138 4686 2141
rect 4606 2132 4609 2138
rect 4554 2128 4558 2131
rect 4486 2112 4489 2118
rect 4522 2108 4529 2111
rect 4526 2092 4529 2108
rect 4622 2092 4625 2118
rect 4686 2112 4689 2128
rect 4694 2122 4697 2128
rect 4702 2122 4705 2128
rect 4726 2122 4729 2188
rect 4734 2142 4737 2158
rect 4766 2152 4769 2158
rect 4758 2142 4761 2148
rect 4774 2142 4777 2238
rect 4790 2182 4793 2218
rect 4830 2162 4833 2168
rect 4862 2152 4865 2188
rect 4794 2148 4798 2151
rect 4822 2142 4825 2148
rect 4846 2142 4849 2148
rect 4870 2142 4873 2178
rect 4898 2158 4902 2161
rect 4918 2151 4921 2218
rect 4934 2192 4937 2248
rect 5030 2242 5033 2268
rect 5134 2262 5137 2268
rect 5062 2242 5065 2248
rect 4990 2212 4993 2218
rect 4950 2172 4953 2178
rect 5078 2172 5081 2218
rect 4986 2168 4990 2171
rect 5030 2162 5033 2168
rect 4930 2158 4934 2161
rect 5018 2158 5022 2161
rect 4918 2148 4926 2151
rect 4962 2148 4966 2151
rect 4954 2138 4958 2141
rect 4746 2128 4750 2131
rect 4462 2088 4470 2091
rect 4166 2042 4169 2058
rect 4198 2041 4201 2078
rect 4226 2068 4230 2071
rect 4206 2052 4209 2068
rect 4246 2062 4249 2068
rect 4222 2052 4225 2058
rect 4210 2048 4214 2051
rect 4254 2042 4257 2078
rect 4550 2072 4553 2078
rect 4598 2072 4601 2078
rect 4638 2075 4641 2108
rect 4750 2092 4753 2118
rect 4806 2112 4809 2128
rect 4862 2122 4865 2138
rect 4790 2092 4793 2098
rect 4662 2088 4670 2091
rect 4682 2088 4686 2091
rect 4850 2088 4854 2091
rect 4654 2072 4657 2088
rect 4662 2072 4665 2088
rect 4886 2082 4889 2138
rect 4898 2128 4902 2131
rect 4902 2072 4905 2088
rect 4274 2068 4278 2071
rect 4490 2068 4494 2071
rect 4338 2058 4342 2061
rect 4542 2062 4545 2068
rect 4278 2042 4281 2048
rect 4198 2038 4209 2041
rect 4166 1992 4169 2028
rect 4206 1992 4209 2038
rect 4122 1958 4126 1961
rect 4126 1942 4129 1958
rect 4270 1951 4273 1998
rect 4318 1972 4321 2058
rect 4406 2052 4409 2059
rect 4570 2038 4574 2041
rect 4440 2003 4442 2007
rect 4446 2003 4449 2007
rect 4453 2003 4456 2007
rect 4510 1952 4513 1958
rect 4182 1942 4185 1948
rect 4418 1948 4422 1951
rect 4382 1942 4385 1948
rect 4106 1938 4110 1941
rect 4410 1938 4414 1941
rect 4442 1938 4446 1941
rect 4190 1922 4193 1938
rect 4090 1918 4094 1921
rect 4142 1892 4145 1918
rect 4238 1912 4241 1938
rect 4254 1902 4257 1938
rect 4350 1932 4353 1938
rect 4394 1928 4398 1931
rect 4342 1902 4345 1928
rect 4110 1872 4113 1878
rect 4158 1872 4161 1878
rect 4166 1872 4169 1888
rect 4182 1872 4185 1878
rect 4190 1872 4193 1888
rect 4246 1882 4249 1898
rect 4306 1888 4310 1891
rect 4358 1891 4361 1918
rect 4358 1888 4366 1891
rect 3982 1792 3985 1859
rect 4046 1842 4049 1848
rect 4054 1842 4057 1868
rect 3982 1752 3985 1788
rect 3966 1738 3974 1741
rect 3798 1712 3801 1728
rect 3806 1692 3809 1718
rect 3830 1702 3833 1728
rect 3706 1668 3710 1671
rect 3678 1652 3681 1668
rect 3678 1612 3681 1648
rect 3702 1642 3705 1668
rect 3666 1558 3670 1561
rect 3686 1552 3689 1558
rect 3714 1548 3718 1551
rect 3630 1542 3633 1547
rect 3590 1498 3601 1501
rect 3546 1488 3550 1491
rect 3546 1478 3550 1481
rect 3518 1472 3521 1478
rect 3574 1472 3577 1478
rect 3582 1461 3585 1468
rect 3554 1458 3585 1461
rect 3558 1392 3561 1418
rect 3530 1388 3534 1391
rect 3478 1358 3489 1361
rect 3434 1348 3438 1351
rect 3454 1272 3457 1338
rect 3466 1278 3470 1281
rect 3478 1272 3481 1348
rect 3486 1282 3489 1358
rect 3494 1271 3497 1338
rect 3486 1268 3497 1271
rect 3342 1262 3345 1268
rect 3358 1261 3361 1268
rect 3390 1262 3393 1268
rect 3358 1258 3369 1261
rect 3334 1192 3337 1208
rect 3206 1062 3209 1068
rect 3198 1052 3201 1058
rect 3122 978 3126 981
rect 3182 972 3185 1048
rect 3150 952 3153 958
rect 3130 948 3134 951
rect 3054 942 3057 947
rect 3086 942 3089 948
rect 3158 942 3161 968
rect 3182 952 3185 958
rect 3198 952 3201 1038
rect 3206 942 3209 1058
rect 3222 1032 3225 1038
rect 3230 1022 3233 1068
rect 3262 1052 3265 1059
rect 3230 952 3233 1018
rect 3310 992 3313 1068
rect 3326 1032 3329 1148
rect 3358 1092 3361 1108
rect 3366 1092 3369 1258
rect 3410 1258 3414 1261
rect 3334 1072 3337 1078
rect 3322 1018 3326 1021
rect 3218 948 3222 951
rect 3242 948 3246 951
rect 3294 942 3297 948
rect 3202 938 3206 941
rect 3090 928 3094 931
rect 3114 928 3118 931
rect 3138 928 3142 931
rect 3026 888 3030 891
rect 3054 882 3057 888
rect 3078 882 3081 888
rect 2974 872 2977 878
rect 3030 872 3033 878
rect 2910 792 2913 868
rect 2942 802 2945 868
rect 3038 862 3041 878
rect 3118 872 3121 878
rect 3126 872 3129 878
rect 3134 872 3137 918
rect 3150 892 3153 938
rect 2954 858 2958 861
rect 2990 852 2993 858
rect 3054 852 3057 858
rect 3078 852 3081 868
rect 3042 848 3046 851
rect 2766 768 2777 771
rect 2250 758 2254 761
rect 2274 758 2278 761
rect 2238 752 2241 758
rect 2278 742 2281 758
rect 2286 752 2289 768
rect 2314 748 2318 751
rect 2222 492 2225 658
rect 2230 561 2233 738
rect 2238 732 2241 738
rect 2254 732 2257 738
rect 2310 732 2313 738
rect 2326 732 2329 768
rect 2478 762 2481 768
rect 2434 758 2438 761
rect 2474 758 2478 761
rect 2610 758 2614 761
rect 2354 748 2358 751
rect 2426 748 2430 751
rect 2466 748 2470 751
rect 2370 738 2374 741
rect 2446 732 2449 738
rect 2454 732 2457 738
rect 2462 732 2465 738
rect 2502 732 2505 738
rect 2434 728 2438 731
rect 2230 558 2241 561
rect 2230 502 2233 548
rect 2238 542 2241 558
rect 2262 552 2265 728
rect 2374 722 2377 728
rect 2278 672 2281 688
rect 2286 682 2289 688
rect 2286 632 2289 678
rect 2294 652 2297 668
rect 2290 548 2294 551
rect 2286 521 2289 538
rect 2282 518 2289 521
rect 2270 502 2273 518
rect 2270 488 2278 491
rect 2014 462 2017 468
rect 2182 462 2185 488
rect 2222 472 2225 478
rect 2270 472 2273 488
rect 2206 462 2209 468
rect 2278 462 2281 468
rect 2002 458 2006 461
rect 1994 448 1998 451
rect 2034 448 2038 451
rect 1950 442 1953 448
rect 1962 438 1966 441
rect 1918 392 1921 398
rect 1910 362 1913 388
rect 1926 372 1929 388
rect 1934 352 1937 368
rect 1950 362 1953 368
rect 1958 352 1961 418
rect 1974 392 1977 428
rect 2086 372 2089 378
rect 1966 332 1969 368
rect 2034 348 2038 351
rect 2062 342 2065 348
rect 1870 272 1873 279
rect 1894 278 1905 281
rect 1778 268 1782 271
rect 1766 262 1769 268
rect 1830 262 1833 268
rect 1854 262 1857 268
rect 1818 258 1822 261
rect 1846 252 1849 258
rect 1810 248 1814 251
rect 1642 238 1646 241
rect 1654 232 1657 248
rect 1654 192 1657 198
rect 1622 162 1625 178
rect 1662 172 1665 198
rect 1710 192 1713 198
rect 1846 192 1849 248
rect 1682 188 1686 191
rect 1778 188 1782 191
rect 1834 188 1838 191
rect 1878 172 1881 258
rect 1758 168 1870 171
rect 1550 142 1553 158
rect 1578 138 1582 141
rect 1510 132 1513 138
rect 1338 88 1342 91
rect 1402 88 1406 91
rect 1302 72 1305 78
rect 1358 72 1361 88
rect 1502 82 1505 88
rect 1474 78 1478 81
rect 1518 72 1521 138
rect 1558 132 1561 138
rect 1598 132 1601 148
rect 1526 82 1529 128
rect 1582 92 1585 128
rect 1606 122 1609 158
rect 1614 148 1622 151
rect 1614 92 1617 148
rect 1630 112 1633 168
rect 1686 162 1689 168
rect 1718 162 1721 168
rect 1758 162 1761 168
rect 1646 122 1649 158
rect 1654 152 1657 158
rect 1694 142 1697 148
rect 1702 132 1705 158
rect 1726 142 1729 148
rect 1726 122 1729 138
rect 1742 132 1745 138
rect 1702 92 1705 118
rect 1734 92 1737 108
rect 1766 92 1769 158
rect 1774 112 1777 148
rect 1790 142 1793 158
rect 1802 138 1806 141
rect 1782 102 1785 138
rect 1814 112 1817 138
rect 1822 132 1825 138
rect 1534 72 1537 78
rect 1630 72 1633 88
rect 1678 82 1681 88
rect 1766 82 1769 88
rect 1218 68 1222 71
rect 1434 68 1438 71
rect 1274 58 1278 61
rect 1102 52 1105 58
rect 1206 52 1209 58
rect 1310 52 1313 68
rect 1382 62 1385 68
rect 1442 58 1446 61
rect 1482 58 1486 61
rect 266 48 270 51
rect 714 48 718 51
rect 1074 48 1078 51
rect 1154 48 1158 51
rect 1242 48 1246 51
rect 1282 48 1286 51
rect 278 42 281 48
rect 702 42 705 48
rect 958 42 961 48
rect 1550 42 1553 68
rect 1562 58 1574 61
rect 1578 58 1582 61
rect 1590 52 1593 68
rect 1618 58 1622 61
rect 1630 52 1633 58
rect 1646 52 1649 78
rect 1670 72 1673 78
rect 1686 72 1689 78
rect 1726 72 1729 78
rect 1758 72 1761 78
rect 1762 68 1766 71
rect 1670 52 1673 68
rect 1678 62 1681 68
rect 1686 62 1689 68
rect 1718 62 1721 68
rect 1750 62 1753 68
rect 1782 62 1785 88
rect 1806 70 1809 88
rect 1814 72 1817 78
rect 1822 72 1825 128
rect 1838 122 1841 148
rect 1830 92 1833 118
rect 1790 62 1793 68
rect 1734 52 1737 58
rect 1782 52 1785 58
rect 1838 52 1841 118
rect 1846 112 1849 118
rect 1854 92 1857 128
rect 1862 122 1865 148
rect 1874 138 1878 141
rect 1872 103 1874 107
rect 1878 103 1881 107
rect 1885 103 1888 107
rect 1618 48 1622 51
rect 1654 42 1657 48
rect 1138 38 1142 41
rect 1578 38 1582 41
rect 1610 38 1614 41
rect 344 3 346 7
rect 350 3 353 7
rect 357 3 360 7
rect 486 -18 489 8
rect 526 -18 529 8
rect 558 -18 561 8
rect 798 -18 801 8
rect 1078 -18 1081 8
rect 1110 -18 1113 8
rect 1174 -18 1177 8
rect 1230 -18 1233 18
rect 1254 -18 1257 8
rect 1278 -18 1281 8
rect 1294 -18 1297 8
rect 1358 -18 1361 8
rect 1368 3 1370 7
rect 1374 3 1377 7
rect 1381 3 1384 7
rect 1390 -18 1393 8
rect 1462 -18 1465 8
rect 1478 -18 1481 8
rect 1638 -18 1641 8
rect 1678 -18 1681 8
rect 1734 -18 1737 8
rect 1798 -18 1801 8
rect 1894 -18 1897 278
rect 1950 272 1953 308
rect 1958 282 1961 298
rect 1982 282 1985 318
rect 1990 272 1993 308
rect 2014 292 2017 298
rect 2054 292 2057 308
rect 2078 302 2081 338
rect 2086 312 2089 348
rect 2034 288 2038 291
rect 2022 272 2025 288
rect 2062 282 2065 298
rect 2094 278 2097 378
rect 2102 362 2105 368
rect 2110 302 2113 348
rect 2118 312 2121 338
rect 2126 332 2129 368
rect 2142 342 2145 438
rect 2254 372 2257 418
rect 2178 368 2182 371
rect 2242 368 2246 371
rect 2182 352 2185 358
rect 2190 332 2193 338
rect 2130 318 2134 321
rect 2206 282 2209 338
rect 2214 302 2217 348
rect 2222 342 2225 358
rect 2234 348 2238 351
rect 2230 332 2233 338
rect 2254 322 2257 338
rect 2218 288 2222 291
rect 2230 272 2233 278
rect 1978 268 1982 271
rect 1902 152 1905 268
rect 1958 262 1961 268
rect 1954 258 1958 261
rect 1994 258 1998 261
rect 2042 258 2046 261
rect 2038 252 2041 258
rect 1918 142 1921 218
rect 1926 192 1929 238
rect 2086 212 2089 218
rect 1978 188 1982 191
rect 2082 188 2086 191
rect 1942 142 1945 188
rect 2030 168 2049 171
rect 2014 141 2017 148
rect 2010 138 2017 141
rect 1910 122 1913 138
rect 1918 132 1921 138
rect 1950 112 1953 128
rect 1958 102 1961 138
rect 2006 121 2009 138
rect 2002 118 2009 121
rect 2030 112 2033 168
rect 2038 142 2041 158
rect 2046 141 2049 168
rect 2110 142 2113 188
rect 2118 162 2121 268
rect 2150 263 2153 268
rect 2182 262 2185 268
rect 2270 262 2273 368
rect 2302 352 2305 698
rect 2318 692 2321 718
rect 2422 712 2425 728
rect 2510 722 2513 758
rect 2534 752 2537 758
rect 2510 702 2513 718
rect 2462 692 2465 698
rect 2318 682 2321 688
rect 2350 672 2353 688
rect 2430 672 2433 678
rect 2438 672 2441 688
rect 2486 682 2489 688
rect 2370 668 2377 671
rect 2330 658 2334 661
rect 2342 652 2345 668
rect 2350 652 2353 658
rect 2366 652 2369 658
rect 2374 652 2377 668
rect 2486 662 2489 668
rect 2502 662 2505 698
rect 2510 662 2513 668
rect 2518 662 2521 668
rect 2442 658 2446 661
rect 2466 658 2470 661
rect 2390 652 2393 658
rect 2494 652 2497 658
rect 2362 648 2366 651
rect 2434 648 2438 651
rect 2322 638 2326 641
rect 2378 638 2382 641
rect 2514 638 2518 641
rect 2310 632 2313 638
rect 2390 632 2393 638
rect 2310 552 2313 588
rect 2318 542 2321 618
rect 2392 603 2394 607
rect 2398 603 2401 607
rect 2405 603 2408 607
rect 2462 592 2465 608
rect 2534 592 2537 748
rect 2550 712 2553 738
rect 2586 718 2590 721
rect 2590 692 2593 698
rect 2606 682 2609 758
rect 2630 722 2633 748
rect 2638 702 2641 738
rect 2646 732 2649 738
rect 2662 732 2665 738
rect 2670 732 2673 768
rect 2694 752 2697 758
rect 2714 748 2718 751
rect 2774 742 2777 768
rect 2838 742 2841 748
rect 2886 742 2889 788
rect 2898 748 2902 751
rect 2934 751 2937 798
rect 3034 758 3038 761
rect 3054 752 3057 818
rect 3062 762 3065 838
rect 3094 822 3097 858
rect 3102 832 3105 868
rect 3110 852 3113 868
rect 3134 842 3137 868
rect 3158 862 3161 878
rect 3150 842 3153 848
rect 3158 842 3161 858
rect 3118 762 3121 798
rect 3134 752 3137 838
rect 2718 702 2721 738
rect 2726 732 2729 738
rect 2782 732 2785 738
rect 2758 712 2761 718
rect 2614 682 2617 698
rect 2630 672 2633 698
rect 2718 692 2721 698
rect 2726 692 2729 698
rect 2766 692 2769 718
rect 2782 692 2785 728
rect 2830 722 2833 738
rect 2814 692 2817 718
rect 2674 688 2678 691
rect 2650 678 2654 681
rect 2546 658 2550 661
rect 2558 658 2566 661
rect 2546 648 2550 651
rect 2558 642 2561 658
rect 2566 632 2569 638
rect 2574 632 2577 648
rect 2582 612 2585 648
rect 2606 642 2609 668
rect 2654 662 2657 668
rect 2334 542 2337 588
rect 2358 562 2361 568
rect 2374 562 2377 588
rect 2430 572 2433 578
rect 2606 572 2609 638
rect 2650 628 2654 631
rect 2538 568 2542 571
rect 2518 562 2521 568
rect 2614 562 2617 568
rect 2630 562 2633 608
rect 2654 592 2657 598
rect 2426 548 2430 551
rect 2414 542 2417 548
rect 2446 542 2449 558
rect 2458 548 2462 551
rect 2530 548 2534 551
rect 2546 548 2550 551
rect 2354 538 2358 541
rect 2398 532 2401 538
rect 2414 532 2417 538
rect 2454 532 2457 538
rect 2486 532 2489 538
rect 2510 522 2513 548
rect 2370 518 2374 521
rect 2526 492 2529 538
rect 2558 512 2561 558
rect 2566 522 2569 548
rect 2574 542 2577 558
rect 2598 541 2601 558
rect 2622 552 2625 558
rect 2594 538 2601 541
rect 2634 548 2638 551
rect 2590 532 2593 538
rect 2606 522 2609 548
rect 2646 522 2649 568
rect 2662 542 2665 688
rect 2782 672 2785 678
rect 2714 668 2718 671
rect 2762 668 2766 671
rect 2798 670 2801 678
rect 2822 672 2825 698
rect 2854 692 2857 708
rect 2904 703 2906 707
rect 2910 703 2913 707
rect 2917 703 2920 707
rect 2934 692 2937 728
rect 2966 702 2969 748
rect 3110 742 3113 748
rect 3150 742 3153 838
rect 3174 761 3177 918
rect 3206 862 3209 888
rect 3222 872 3225 928
rect 3254 922 3257 938
rect 3270 932 3273 938
rect 3290 928 3294 931
rect 3230 902 3233 918
rect 3214 792 3217 868
rect 3222 862 3225 868
rect 3262 862 3265 898
rect 3286 872 3289 898
rect 3326 881 3329 928
rect 3334 922 3337 938
rect 3342 902 3345 1058
rect 3350 962 3353 1018
rect 3370 968 3374 971
rect 3382 952 3385 1218
rect 3390 1142 3393 1258
rect 3416 1203 3418 1207
rect 3422 1203 3425 1207
rect 3429 1203 3432 1207
rect 3398 1151 3401 1158
rect 3434 1148 3438 1151
rect 3466 1148 3470 1151
rect 3478 1142 3481 1218
rect 3386 948 3390 951
rect 3354 888 3358 891
rect 3326 878 3337 881
rect 3334 872 3337 878
rect 3342 872 3345 878
rect 3306 868 3313 871
rect 3254 852 3257 858
rect 3274 838 3278 841
rect 3278 822 3281 828
rect 3174 758 3185 761
rect 3182 752 3185 758
rect 3170 748 3174 751
rect 3162 738 3166 741
rect 3054 692 3057 738
rect 3126 732 3129 738
rect 3146 728 3150 731
rect 3090 718 3094 721
rect 3126 692 3129 708
rect 3158 702 3161 718
rect 2834 688 2838 691
rect 2862 672 2865 678
rect 3086 672 3089 678
rect 2670 652 2673 668
rect 2686 662 2689 668
rect 2726 662 2729 668
rect 2734 662 2737 668
rect 2790 662 2793 668
rect 2886 662 2889 668
rect 2910 662 2913 668
rect 2970 658 2974 661
rect 2678 652 2681 658
rect 2710 652 2713 658
rect 2726 652 2729 658
rect 2734 652 2737 658
rect 2766 652 2769 658
rect 2822 652 2825 658
rect 2834 648 2838 651
rect 2690 638 2694 641
rect 2742 592 2745 608
rect 2758 592 2761 638
rect 2766 602 2769 648
rect 2870 642 2873 658
rect 2878 652 2881 658
rect 2998 652 3001 668
rect 3030 662 3033 668
rect 3018 658 3022 661
rect 3026 648 3030 651
rect 2814 592 2817 598
rect 2850 558 2854 561
rect 2694 552 2697 558
rect 2722 548 2726 551
rect 2778 548 2782 551
rect 2818 548 2825 551
rect 2734 542 2737 548
rect 2722 538 2726 541
rect 2710 521 2713 538
rect 2710 518 2718 521
rect 2354 468 2358 471
rect 2446 462 2449 468
rect 2462 463 2465 468
rect 2418 458 2422 461
rect 2542 462 2545 468
rect 2258 258 2262 261
rect 2174 162 2177 238
rect 2118 142 2121 158
rect 2174 142 2177 158
rect 2190 142 2193 148
rect 2046 138 2054 141
rect 2162 138 2166 141
rect 2042 128 2046 131
rect 2062 131 2065 138
rect 2054 128 2065 131
rect 2134 132 2137 138
rect 2142 132 2145 138
rect 2178 128 2182 131
rect 2054 92 2057 128
rect 2118 112 2121 118
rect 2086 92 2089 108
rect 1942 72 1945 78
rect 2070 72 2073 78
rect 1918 62 1921 68
rect 1910 58 1918 61
rect 2006 59 2014 61
rect 2018 59 2022 62
rect 2038 62 2041 68
rect 2006 58 2017 59
rect 1910 -18 1913 58
rect 1958 42 1961 58
rect 2006 -18 2009 58
rect 2078 52 2081 78
rect 2102 72 2105 78
rect 2158 62 2161 68
rect 2190 63 2193 68
rect 2246 63 2249 208
rect 2270 152 2273 198
rect 2090 48 2094 51
rect 2046 -18 2049 8
rect 2062 -18 2065 18
rect 2078 -18 2081 28
rect 2094 -18 2097 38
rect 2126 -18 2129 8
rect 2150 -18 2153 8
rect 2182 -18 2185 8
rect 2198 -18 2201 8
rect 2214 -18 2217 28
rect 2246 22 2249 59
rect 2246 -18 2249 8
rect 2262 -18 2265 68
rect 2270 12 2273 148
rect 2278 -18 2281 258
rect 2294 142 2297 238
rect 2302 202 2305 348
rect 2334 342 2337 458
rect 2558 452 2561 459
rect 2392 403 2394 407
rect 2398 403 2401 407
rect 2405 403 2408 407
rect 2370 348 2374 351
rect 2402 348 2406 351
rect 2402 338 2406 341
rect 2310 292 2313 308
rect 2334 301 2337 338
rect 2334 298 2345 301
rect 2342 282 2345 298
rect 2350 292 2353 338
rect 2350 262 2353 278
rect 2414 232 2417 398
rect 2442 378 2446 381
rect 2486 352 2489 368
rect 2510 342 2513 348
rect 2422 292 2425 338
rect 2470 332 2473 338
rect 2478 322 2481 338
rect 2466 318 2470 321
rect 2510 312 2513 328
rect 2518 322 2521 328
rect 2430 272 2433 308
rect 2458 288 2462 291
rect 2478 282 2481 298
rect 2526 292 2529 438
rect 2542 392 2545 428
rect 2574 392 2577 508
rect 2622 492 2625 498
rect 2602 388 2606 391
rect 2534 352 2537 368
rect 2534 322 2537 338
rect 2542 332 2545 348
rect 2558 342 2561 358
rect 2566 342 2569 348
rect 2566 322 2569 338
rect 2574 332 2577 348
rect 2606 342 2609 368
rect 2614 342 2617 488
rect 2630 482 2633 498
rect 2670 492 2673 518
rect 2714 488 2718 491
rect 2666 478 2673 481
rect 2630 382 2633 468
rect 2630 362 2633 378
rect 2638 362 2641 388
rect 2654 382 2657 418
rect 2662 392 2665 468
rect 2654 372 2657 378
rect 2670 372 2673 478
rect 2698 468 2702 471
rect 2678 382 2681 468
rect 2698 458 2702 461
rect 2678 372 2681 378
rect 2670 362 2673 368
rect 2686 352 2689 458
rect 2718 442 2721 478
rect 2726 462 2729 508
rect 2734 492 2737 538
rect 2750 492 2753 528
rect 2790 492 2793 538
rect 2798 522 2801 528
rect 2750 472 2753 488
rect 2782 482 2785 488
rect 2766 478 2774 481
rect 2758 472 2761 478
rect 2766 472 2769 478
rect 2806 471 2809 538
rect 2822 472 2825 548
rect 2830 532 2833 558
rect 2838 522 2841 538
rect 2806 468 2814 471
rect 2734 432 2737 468
rect 2758 442 2761 458
rect 2694 392 2697 428
rect 2766 392 2769 468
rect 2774 462 2777 468
rect 2798 462 2801 468
rect 2806 452 2809 458
rect 2814 442 2817 468
rect 2822 462 2825 468
rect 2838 462 2841 488
rect 2830 452 2833 458
rect 2838 452 2841 458
rect 2806 392 2809 428
rect 2838 412 2841 448
rect 2846 441 2849 468
rect 2854 462 2857 518
rect 2862 492 2865 588
rect 2878 552 2881 648
rect 2942 642 2945 648
rect 2950 642 2953 648
rect 2898 638 2902 641
rect 2886 632 2889 638
rect 2982 632 2985 648
rect 2998 582 3001 648
rect 3038 612 3041 668
rect 3094 662 3097 668
rect 3030 592 3033 598
rect 3038 572 3041 608
rect 3094 592 3097 658
rect 2894 552 2897 568
rect 2990 562 2993 568
rect 2958 552 2961 558
rect 2974 552 2977 558
rect 2946 548 2950 551
rect 3002 548 3006 551
rect 2870 492 2873 518
rect 2878 492 2881 528
rect 2904 503 2906 507
rect 2910 503 2913 507
rect 2917 503 2920 507
rect 2926 492 2929 528
rect 2942 512 2945 528
rect 2958 522 2961 538
rect 2958 482 2961 498
rect 2914 478 2918 481
rect 2870 462 2873 478
rect 2974 472 2977 548
rect 3014 542 3017 548
rect 3022 532 3025 558
rect 3046 552 3049 588
rect 3106 568 3110 571
rect 3058 558 3062 561
rect 3058 538 3062 541
rect 3078 532 3081 538
rect 3086 492 3089 558
rect 3094 542 3097 548
rect 2954 468 2958 471
rect 2878 462 2881 468
rect 3094 462 3097 518
rect 3102 472 3105 548
rect 3118 542 3121 618
rect 3142 592 3145 668
rect 3150 662 3153 698
rect 3174 692 3177 748
rect 3190 742 3193 748
rect 3198 732 3201 758
rect 3214 742 3217 788
rect 3230 742 3233 747
rect 3262 722 3265 748
rect 3278 742 3281 818
rect 3294 792 3297 858
rect 3302 852 3305 858
rect 3310 852 3313 868
rect 3322 858 3326 861
rect 3326 822 3329 828
rect 3310 762 3313 768
rect 3326 752 3329 818
rect 3334 752 3337 868
rect 3342 842 3345 868
rect 3366 792 3369 848
rect 3374 832 3377 948
rect 3406 941 3409 1078
rect 3446 1072 3449 1098
rect 3470 1082 3473 1138
rect 3430 1063 3433 1068
rect 3478 1062 3481 1118
rect 3486 1092 3489 1268
rect 3534 1261 3537 1348
rect 3546 1338 3550 1341
rect 3566 1332 3569 1388
rect 3590 1362 3593 1498
rect 3606 1482 3609 1488
rect 3606 1462 3609 1468
rect 3622 1462 3625 1518
rect 3630 1502 3633 1528
rect 3646 1482 3649 1548
rect 3678 1532 3681 1538
rect 3666 1518 3670 1521
rect 3686 1512 3689 1548
rect 3702 1532 3705 1538
rect 3634 1478 3641 1481
rect 3590 1352 3593 1358
rect 3622 1352 3625 1418
rect 3594 1338 3598 1341
rect 3554 1328 3558 1331
rect 3602 1328 3606 1331
rect 3542 1302 3545 1318
rect 3566 1292 3569 1328
rect 3542 1272 3545 1278
rect 3530 1258 3537 1261
rect 3550 1262 3553 1288
rect 3562 1278 3566 1281
rect 3574 1271 3577 1318
rect 3622 1292 3625 1348
rect 3638 1292 3641 1478
rect 3678 1462 3681 1468
rect 3646 1422 3649 1458
rect 3654 1452 3657 1458
rect 3686 1452 3689 1458
rect 3654 1392 3657 1438
rect 3702 1432 3705 1528
rect 3650 1358 3654 1361
rect 3710 1332 3713 1468
rect 3718 1452 3721 1518
rect 3726 1492 3729 1548
rect 3730 1468 3734 1471
rect 3742 1471 3745 1668
rect 3774 1663 3777 1688
rect 3850 1668 3854 1671
rect 3758 1551 3761 1558
rect 3790 1552 3793 1668
rect 3786 1548 3790 1551
rect 3822 1522 3825 1538
rect 3750 1492 3753 1508
rect 3738 1468 3745 1471
rect 3774 1462 3777 1488
rect 3786 1478 3790 1481
rect 3830 1472 3833 1668
rect 3838 1632 3841 1658
rect 3838 1502 3841 1518
rect 3862 1512 3865 1728
rect 3886 1492 3889 1688
rect 3898 1628 3902 1631
rect 3910 1552 3913 1738
rect 3928 1703 3930 1707
rect 3934 1703 3937 1707
rect 3941 1703 3944 1707
rect 3962 1668 3966 1671
rect 3950 1652 3953 1658
rect 3914 1548 3918 1551
rect 3898 1538 3902 1541
rect 3894 1462 3897 1468
rect 3918 1462 3921 1508
rect 3928 1503 3930 1507
rect 3934 1503 3937 1507
rect 3941 1503 3944 1507
rect 3966 1492 3969 1598
rect 3974 1542 3977 1738
rect 4006 1692 4009 1718
rect 4014 1692 4017 1828
rect 4062 1792 4065 1808
rect 4070 1742 4073 1818
rect 4086 1752 4089 1818
rect 4102 1792 4105 1868
rect 4190 1862 4193 1868
rect 4198 1862 4201 1878
rect 4238 1872 4241 1878
rect 4254 1872 4257 1878
rect 4270 1872 4273 1888
rect 4278 1870 4281 1878
rect 4238 1862 4241 1868
rect 4298 1868 4302 1871
rect 4310 1862 4313 1868
rect 4342 1862 4345 1878
rect 4354 1868 4358 1871
rect 4386 1868 4390 1871
rect 4258 1858 4262 1861
rect 4350 1858 4358 1861
rect 4182 1852 4185 1858
rect 4326 1852 4329 1858
rect 4210 1838 4214 1841
rect 4226 1838 4230 1841
rect 4182 1752 4185 1838
rect 4214 1802 4217 1818
rect 4190 1762 4193 1768
rect 4198 1762 4201 1788
rect 4202 1748 4206 1751
rect 4182 1742 4185 1748
rect 4214 1742 4217 1788
rect 4238 1762 4241 1798
rect 4266 1768 4270 1771
rect 4278 1762 4281 1798
rect 4282 1748 4286 1751
rect 4254 1742 4257 1748
rect 4294 1742 4297 1758
rect 4310 1752 4313 1818
rect 4334 1752 4337 1798
rect 4350 1772 4353 1778
rect 4350 1762 4353 1768
rect 4358 1762 4361 1778
rect 4366 1772 4369 1868
rect 4398 1862 4401 1878
rect 4382 1762 4385 1798
rect 4342 1752 4345 1758
rect 4362 1748 4366 1751
rect 4406 1742 4409 1918
rect 4470 1912 4473 1928
rect 4486 1922 4489 1948
rect 4510 1922 4513 1938
rect 4534 1922 4537 1940
rect 4414 1882 4417 1898
rect 4422 1882 4425 1898
rect 4450 1858 4454 1861
rect 4462 1842 4465 1868
rect 4470 1852 4473 1898
rect 4494 1862 4497 1918
rect 4518 1872 4521 1918
rect 4550 1902 4553 1938
rect 4570 1918 4574 1921
rect 4598 1902 4601 1938
rect 4526 1882 4529 1898
rect 4482 1858 4486 1861
rect 4534 1852 4537 1878
rect 4558 1862 4561 1868
rect 4590 1862 4593 1868
rect 4582 1852 4585 1858
rect 4578 1848 4582 1851
rect 4606 1851 4609 1918
rect 4614 1882 4617 1898
rect 4602 1848 4609 1851
rect 4490 1838 4494 1841
rect 4570 1838 4574 1841
rect 4602 1838 4606 1841
rect 4502 1832 4505 1838
rect 4414 1762 4417 1768
rect 4422 1751 4425 1818
rect 4440 1803 4442 1807
rect 4446 1803 4449 1807
rect 4453 1803 4456 1807
rect 4478 1782 4481 1818
rect 4542 1772 4545 1818
rect 4434 1758 4438 1761
rect 4486 1752 4489 1768
rect 4542 1752 4545 1758
rect 4418 1748 4430 1751
rect 4046 1672 4049 1738
rect 4054 1722 4057 1728
rect 4118 1722 4121 1738
rect 4126 1732 4129 1738
rect 4230 1732 4233 1738
rect 4382 1732 4385 1738
rect 4430 1732 4433 1748
rect 4510 1742 4513 1748
rect 4442 1738 4446 1741
rect 4558 1741 4561 1818
rect 4582 1762 4585 1768
rect 4590 1742 4593 1818
rect 4598 1752 4601 1758
rect 4614 1752 4617 1858
rect 4622 1851 4625 1948
rect 4686 1942 4689 2048
rect 4710 1982 4713 2068
rect 4718 2062 4721 2068
rect 4766 2062 4769 2068
rect 4774 2052 4777 2068
rect 4822 2042 4825 2068
rect 4830 2032 4833 2068
rect 4910 2062 4913 2138
rect 4926 2092 4929 2138
rect 4952 2103 4954 2107
rect 4958 2103 4961 2107
rect 4965 2103 4968 2107
rect 4958 2072 4961 2088
rect 4990 2072 4993 2118
rect 4998 2112 5001 2148
rect 5014 2132 5017 2138
rect 5022 2081 5025 2158
rect 5058 2138 5062 2141
rect 5030 2122 5033 2138
rect 5070 2131 5073 2158
rect 5086 2152 5089 2248
rect 5142 2202 5145 2268
rect 5150 2262 5153 2268
rect 5174 2262 5177 2268
rect 5218 2258 5222 2261
rect 5146 2188 5150 2191
rect 5190 2182 5193 2258
rect 5250 2248 5254 2251
rect 5206 2192 5209 2238
rect 5262 2222 5265 2228
rect 5094 2142 5097 2168
rect 5102 2162 5105 2168
rect 5118 2162 5121 2178
rect 5122 2158 5129 2161
rect 5082 2138 5086 2141
rect 5066 2128 5073 2131
rect 5062 2102 5065 2128
rect 5074 2118 5078 2121
rect 5086 2092 5089 2098
rect 5094 2082 5097 2138
rect 5102 2132 5105 2148
rect 5126 2132 5129 2158
rect 5190 2152 5193 2178
rect 5214 2172 5217 2178
rect 5198 2162 5201 2168
rect 5202 2148 5206 2151
rect 5214 2142 5217 2168
rect 5182 2132 5185 2138
rect 5162 2128 5166 2131
rect 5110 2082 5113 2108
rect 5022 2078 5030 2081
rect 5046 2072 5049 2078
rect 5002 2068 5006 2071
rect 4982 2062 4985 2068
rect 5022 2032 5025 2048
rect 5054 2022 5057 2028
rect 5014 2012 5017 2018
rect 5070 2012 5073 2058
rect 5078 2052 5081 2068
rect 5094 2062 5097 2068
rect 5110 2062 5113 2078
rect 5174 2072 5177 2078
rect 5222 2072 5225 2208
rect 5230 2152 5233 2158
rect 5254 2152 5257 2168
rect 5250 2148 5254 2151
rect 5250 2138 5254 2141
rect 5234 2128 5238 2131
rect 5250 2128 5254 2131
rect 5094 2022 5097 2048
rect 5118 2022 5121 2068
rect 4798 1942 4801 2008
rect 5006 1992 5009 1998
rect 5038 1992 5041 2008
rect 5078 1992 5081 2018
rect 4946 1988 4950 1991
rect 4838 1962 4841 1968
rect 4886 1951 4889 1988
rect 5042 1958 5046 1961
rect 4806 1942 4809 1948
rect 4914 1948 4918 1951
rect 5026 1938 5030 1941
rect 4630 1902 4633 1938
rect 4638 1902 4641 1938
rect 4654 1882 4657 1918
rect 4686 1912 4689 1938
rect 4694 1921 4697 1938
rect 4742 1932 4745 1938
rect 4694 1918 4702 1921
rect 4770 1918 4774 1921
rect 4638 1862 4641 1878
rect 4686 1872 4689 1888
rect 4710 1872 4713 1918
rect 4718 1882 4721 1898
rect 4758 1875 4761 1908
rect 4854 1892 4857 1938
rect 4952 1903 4954 1907
rect 4958 1903 4961 1907
rect 4965 1903 4968 1907
rect 4974 1892 4977 1938
rect 5054 1932 5057 1958
rect 5142 1952 5145 2028
rect 5166 2002 5169 2068
rect 5250 2058 5254 2061
rect 5230 2052 5233 2058
rect 5194 2038 5198 2041
rect 5170 1988 5174 1991
rect 5198 1952 5201 2018
rect 5210 1958 5214 1961
rect 5094 1942 5097 1948
rect 5062 1932 5065 1938
rect 4998 1892 5001 1932
rect 5110 1922 5113 1947
rect 4782 1888 4790 1891
rect 4802 1888 4806 1891
rect 4922 1888 4926 1891
rect 5050 1888 5054 1891
rect 4774 1872 4777 1888
rect 4782 1872 4785 1888
rect 4894 1872 4897 1878
rect 5014 1872 5017 1878
rect 5022 1872 5025 1878
rect 5078 1872 5081 1878
rect 4674 1868 4678 1871
rect 4834 1868 4838 1871
rect 4662 1862 4665 1868
rect 4694 1862 4697 1868
rect 4630 1852 4633 1858
rect 4622 1848 4630 1851
rect 4674 1848 4678 1851
rect 4694 1842 4697 1858
rect 4710 1852 4713 1868
rect 4886 1862 4889 1868
rect 4942 1862 4945 1868
rect 4638 1802 4641 1818
rect 4622 1762 4625 1768
rect 4634 1758 4638 1761
rect 4662 1752 4665 1778
rect 4682 1758 4686 1761
rect 4554 1738 4561 1741
rect 4570 1738 4574 1741
rect 4610 1738 4614 1741
rect 4510 1732 4513 1738
rect 4490 1728 4494 1731
rect 4546 1728 4550 1731
rect 4086 1702 4089 1718
rect 4142 1712 4145 1718
rect 4110 1672 4113 1678
rect 4166 1672 4169 1678
rect 3994 1538 3998 1541
rect 4006 1492 4009 1668
rect 4046 1662 4049 1668
rect 4078 1621 4081 1659
rect 4158 1642 4161 1668
rect 4214 1662 4217 1668
rect 4222 1652 4225 1718
rect 4254 1682 4257 1688
rect 4230 1662 4233 1668
rect 4270 1662 4273 1718
rect 4286 1672 4289 1678
rect 4294 1672 4297 1718
rect 4286 1652 4289 1668
rect 4302 1652 4305 1728
rect 4462 1722 4465 1728
rect 4558 1722 4561 1728
rect 4314 1658 4318 1661
rect 4334 1652 4337 1698
rect 4382 1682 4385 1718
rect 4462 1692 4465 1708
rect 4470 1702 4473 1718
rect 4526 1682 4529 1718
rect 4346 1678 4350 1681
rect 4346 1668 4350 1671
rect 4358 1662 4361 1678
rect 4422 1672 4425 1678
rect 4394 1668 4398 1671
rect 4410 1668 4414 1671
rect 4342 1652 4345 1658
rect 4258 1648 4262 1651
rect 4446 1642 4449 1668
rect 4242 1638 4246 1641
rect 4362 1638 4366 1641
rect 4078 1618 4089 1621
rect 4018 1548 4022 1551
rect 4018 1538 4022 1541
rect 4006 1482 4009 1488
rect 4070 1482 4073 1488
rect 3766 1452 3769 1458
rect 3822 1452 3825 1459
rect 3782 1442 3785 1448
rect 3754 1358 3758 1361
rect 3718 1351 3721 1358
rect 3766 1352 3769 1428
rect 3790 1352 3793 1398
rect 3806 1362 3809 1428
rect 3846 1392 3849 1398
rect 3786 1338 3790 1341
rect 3646 1312 3649 1318
rect 3590 1272 3593 1288
rect 3654 1272 3657 1288
rect 3570 1268 3582 1271
rect 3642 1268 3646 1271
rect 3558 1262 3561 1268
rect 3502 1252 3505 1258
rect 3526 1232 3529 1258
rect 3582 1252 3585 1268
rect 3590 1262 3593 1268
rect 3614 1262 3617 1268
rect 3654 1262 3657 1268
rect 3610 1248 3614 1251
rect 3502 1162 3505 1218
rect 3498 1128 3502 1131
rect 3494 1082 3497 1118
rect 3526 1112 3529 1158
rect 3534 1142 3537 1248
rect 3622 1222 3625 1258
rect 3594 1158 3598 1161
rect 3546 1148 3550 1151
rect 3542 1142 3545 1148
rect 3558 1142 3561 1158
rect 3582 1142 3585 1148
rect 3606 1142 3609 1158
rect 3630 1151 3633 1168
rect 3626 1148 3633 1151
rect 3622 1132 3625 1148
rect 3610 1128 3614 1131
rect 3502 1092 3505 1108
rect 3416 1003 3418 1007
rect 3422 1003 3425 1007
rect 3429 1003 3432 1007
rect 3478 992 3481 1058
rect 3494 1042 3497 1078
rect 3558 1062 3561 1078
rect 3566 1072 3569 1118
rect 3574 1112 3577 1128
rect 3582 1072 3585 1098
rect 3638 1092 3641 1218
rect 3614 1082 3617 1088
rect 3638 1082 3641 1088
rect 3662 1082 3665 1308
rect 3670 1271 3673 1298
rect 3682 1278 3686 1281
rect 3670 1268 3678 1271
rect 3694 1262 3697 1308
rect 3702 1272 3705 1278
rect 3682 1258 3686 1261
rect 3710 1252 3713 1328
rect 3734 1292 3737 1338
rect 3774 1332 3777 1338
rect 3806 1332 3809 1358
rect 3822 1352 3825 1358
rect 3886 1352 3889 1358
rect 3826 1338 3830 1341
rect 3798 1282 3801 1288
rect 3718 1272 3721 1278
rect 3786 1258 3790 1261
rect 3746 1158 3750 1161
rect 3774 1152 3777 1158
rect 3690 1147 3694 1150
rect 3726 1142 3729 1148
rect 3710 1102 3713 1138
rect 3726 1122 3729 1128
rect 3742 1082 3745 1088
rect 3626 1078 3630 1081
rect 3682 1078 3686 1081
rect 3662 1072 3665 1078
rect 3602 1068 3606 1071
rect 3574 992 3577 1018
rect 3482 968 3486 971
rect 3426 958 3430 961
rect 3534 958 3542 961
rect 3470 942 3473 948
rect 3494 942 3497 948
rect 3406 938 3414 941
rect 3382 862 3385 878
rect 3390 872 3393 918
rect 3422 902 3425 928
rect 3462 922 3465 928
rect 3402 878 3406 881
rect 3422 872 3425 898
rect 3494 892 3497 938
rect 3502 932 3505 958
rect 3534 952 3537 958
rect 3510 922 3513 928
rect 3518 912 3521 918
rect 3518 892 3521 898
rect 3474 888 3478 891
rect 3510 882 3513 888
rect 3434 878 3438 881
rect 3458 878 3462 881
rect 3482 878 3486 881
rect 3434 868 3438 871
rect 3478 862 3481 868
rect 3458 858 3462 861
rect 3416 803 3418 807
rect 3422 803 3425 807
rect 3429 803 3432 807
rect 3350 762 3353 788
rect 3454 762 3457 788
rect 3458 758 3462 761
rect 3314 738 3318 741
rect 3214 672 3217 678
rect 3230 662 3233 668
rect 3254 662 3257 698
rect 3326 692 3329 748
rect 3306 688 3310 691
rect 3334 672 3337 748
rect 3374 742 3377 748
rect 3382 742 3385 748
rect 3390 742 3393 758
rect 3418 748 3422 751
rect 3430 742 3433 758
rect 3458 748 3462 751
rect 3402 738 3406 741
rect 3402 728 3406 731
rect 3350 672 3353 718
rect 3154 658 3158 661
rect 3150 552 3153 658
rect 3318 652 3321 658
rect 3350 602 3353 668
rect 3366 663 3369 718
rect 3430 692 3433 728
rect 3446 692 3449 748
rect 3470 742 3473 768
rect 3502 762 3505 768
rect 3526 752 3529 948
rect 3534 932 3537 938
rect 3542 902 3545 948
rect 3566 862 3569 908
rect 3582 882 3585 1068
rect 3622 1062 3625 1068
rect 3590 952 3593 1028
rect 3646 992 3649 1048
rect 3694 1042 3697 1068
rect 3766 1062 3769 1108
rect 3730 1058 3734 1061
rect 3702 1052 3705 1058
rect 3758 1052 3761 1058
rect 3642 968 3646 971
rect 3614 962 3617 968
rect 3614 942 3617 948
rect 3622 942 3625 958
rect 3630 952 3633 968
rect 3594 938 3598 941
rect 3654 932 3657 1038
rect 3670 972 3673 1018
rect 3694 982 3697 988
rect 3670 962 3673 968
rect 3670 948 3678 951
rect 3618 878 3622 881
rect 3630 852 3633 868
rect 3638 862 3641 898
rect 3670 892 3673 948
rect 3710 932 3713 1038
rect 3774 1022 3777 1138
rect 3782 1122 3785 1128
rect 3798 1112 3801 1128
rect 3726 992 3729 1018
rect 3758 952 3761 958
rect 3722 948 3726 951
rect 3718 902 3721 938
rect 3726 892 3729 928
rect 3774 892 3777 968
rect 3814 962 3817 1338
rect 3830 1292 3833 1318
rect 3894 1282 3897 1338
rect 3950 1321 3953 1478
rect 3974 1462 3977 1468
rect 4014 1402 4017 1458
rect 4078 1431 4081 1518
rect 4086 1512 4089 1618
rect 4194 1618 4198 1621
rect 4126 1592 4129 1618
rect 4150 1592 4153 1608
rect 4094 1542 4097 1578
rect 4142 1542 4145 1588
rect 4246 1562 4249 1618
rect 4210 1547 4214 1550
rect 4246 1542 4249 1548
rect 4302 1542 4305 1618
rect 4382 1552 4385 1618
rect 4440 1603 4442 1607
rect 4446 1603 4449 1607
rect 4453 1603 4456 1607
rect 4494 1572 4497 1668
rect 4502 1662 4505 1668
rect 4518 1662 4521 1668
rect 4526 1652 4529 1668
rect 4534 1662 4537 1668
rect 4558 1652 4561 1688
rect 4594 1678 4598 1681
rect 4574 1662 4577 1678
rect 4594 1668 4598 1671
rect 4582 1662 4585 1668
rect 4586 1658 4593 1661
rect 4514 1648 4518 1651
rect 4502 1642 4505 1648
rect 4534 1571 4537 1618
rect 4526 1568 4537 1571
rect 4410 1548 4414 1551
rect 4358 1542 4361 1548
rect 4422 1542 4425 1558
rect 4478 1552 4481 1558
rect 4506 1548 4510 1551
rect 4486 1542 4489 1548
rect 4526 1542 4529 1568
rect 4562 1558 4566 1561
rect 4534 1552 4537 1558
rect 4574 1552 4577 1618
rect 4410 1538 4414 1541
rect 4102 1492 4105 1508
rect 4110 1481 4113 1518
rect 4102 1478 4113 1481
rect 4086 1472 4089 1478
rect 4086 1452 4089 1458
rect 4078 1428 4089 1431
rect 4046 1392 4049 1418
rect 4078 1362 4081 1418
rect 4086 1352 4089 1428
rect 3950 1318 3961 1321
rect 3928 1303 3930 1307
rect 3934 1303 3937 1307
rect 3941 1303 3944 1307
rect 3958 1292 3961 1318
rect 3966 1292 3969 1348
rect 3982 1342 3985 1347
rect 4014 1342 4017 1348
rect 3894 1263 3897 1268
rect 3934 1192 3937 1288
rect 3958 1282 3961 1288
rect 4030 1282 4033 1348
rect 4086 1342 4089 1348
rect 4094 1342 4097 1478
rect 4102 1382 4105 1478
rect 4134 1462 4137 1478
rect 4174 1472 4177 1488
rect 4214 1472 4217 1528
rect 4266 1518 4270 1521
rect 4286 1492 4289 1508
rect 4294 1492 4297 1538
rect 4318 1502 4321 1518
rect 4258 1488 4262 1491
rect 4342 1472 4345 1518
rect 4350 1512 4353 1538
rect 4518 1532 4521 1538
rect 4442 1528 4446 1531
rect 4490 1528 4494 1531
rect 4486 1522 4489 1528
rect 4374 1512 4377 1518
rect 4374 1482 4377 1488
rect 4150 1462 4153 1468
rect 4114 1458 4118 1461
rect 4158 1452 4161 1468
rect 4202 1458 4206 1461
rect 4146 1448 4150 1451
rect 4126 1392 4129 1438
rect 4094 1292 4097 1338
rect 4102 1292 4105 1348
rect 4094 1282 4097 1288
rect 4134 1272 4137 1418
rect 4142 1392 4145 1438
rect 4150 1412 4153 1418
rect 4150 1392 4153 1398
rect 4158 1302 4161 1448
rect 4262 1432 4265 1468
rect 4178 1358 4182 1361
rect 4198 1352 4201 1408
rect 4270 1392 4273 1458
rect 4294 1452 4297 1458
rect 4222 1362 4225 1368
rect 4294 1362 4297 1428
rect 4310 1422 4313 1468
rect 4318 1462 4321 1468
rect 4358 1451 4361 1478
rect 4406 1472 4409 1498
rect 4414 1492 4417 1508
rect 4414 1482 4417 1488
rect 4430 1472 4433 1518
rect 4454 1462 4457 1468
rect 4470 1462 4473 1488
rect 4478 1462 4481 1468
rect 4494 1462 4497 1478
rect 4502 1472 4505 1518
rect 4510 1512 4513 1528
rect 4510 1472 4513 1478
rect 4358 1448 4366 1451
rect 4434 1448 4438 1451
rect 4318 1382 4321 1448
rect 4354 1388 4358 1391
rect 4214 1352 4217 1358
rect 4262 1352 4265 1358
rect 4294 1351 4297 1358
rect 4290 1348 4297 1351
rect 4302 1352 4305 1358
rect 4166 1312 4169 1348
rect 4214 1332 4217 1338
rect 4230 1332 4233 1348
rect 4258 1338 4262 1341
rect 4238 1332 4241 1338
rect 4270 1331 4273 1338
rect 4266 1328 4273 1331
rect 4238 1301 4241 1328
rect 4246 1312 4249 1318
rect 4230 1298 4241 1301
rect 4230 1282 4233 1298
rect 4242 1288 4246 1291
rect 3954 1258 3958 1261
rect 3942 1151 3945 1258
rect 3830 1142 3833 1148
rect 3942 1148 3950 1151
rect 3954 1148 3958 1151
rect 3986 1148 3990 1151
rect 3862 1142 3865 1147
rect 3998 1142 4001 1158
rect 4006 1142 4009 1158
rect 3830 1092 3833 1128
rect 3846 1102 3849 1138
rect 3822 1062 3825 1078
rect 3846 1062 3849 1098
rect 3854 992 3857 1008
rect 3806 952 3809 958
rect 3782 902 3785 948
rect 3790 942 3793 948
rect 3814 942 3817 958
rect 3822 942 3825 968
rect 3846 962 3849 968
rect 3834 958 3838 961
rect 3854 952 3857 968
rect 3862 952 3865 968
rect 3838 882 3841 918
rect 3870 892 3873 1138
rect 3958 1132 3961 1138
rect 3974 1132 3977 1138
rect 3882 1088 3886 1091
rect 3910 1072 3913 1128
rect 3928 1103 3930 1107
rect 3934 1103 3937 1107
rect 3941 1103 3944 1107
rect 3966 1082 3969 1118
rect 3990 1092 3993 1138
rect 3998 1132 4001 1138
rect 4014 1092 4017 1258
rect 4062 1222 4065 1258
rect 4042 1158 4046 1161
rect 4030 1142 4033 1158
rect 4054 1152 4057 1188
rect 3886 992 3889 1058
rect 3902 1042 3905 1048
rect 3910 1012 3913 1068
rect 3934 1052 3937 1068
rect 3962 1058 3966 1061
rect 3934 1022 3937 1048
rect 3934 962 3937 1018
rect 3974 962 3977 1088
rect 4022 1082 4025 1088
rect 4030 1072 4033 1138
rect 4046 1132 4049 1138
rect 4070 1082 4073 1118
rect 4094 1082 4097 1178
rect 4102 1152 4105 1158
rect 4110 1152 4113 1218
rect 4118 1152 4121 1218
rect 4134 1152 4137 1268
rect 4150 1172 4153 1248
rect 4190 1192 4193 1258
rect 4198 1182 4201 1268
rect 4254 1262 4257 1278
rect 4262 1262 4265 1328
rect 4278 1272 4281 1348
rect 4298 1328 4302 1331
rect 4310 1272 4313 1338
rect 4326 1331 4329 1348
rect 4334 1342 4337 1388
rect 4366 1362 4369 1448
rect 4390 1442 4393 1448
rect 4440 1403 4442 1407
rect 4446 1403 4449 1407
rect 4453 1403 4456 1407
rect 4462 1372 4465 1458
rect 4470 1452 4473 1458
rect 4510 1452 4513 1468
rect 4482 1448 4486 1451
rect 4470 1392 4473 1418
rect 4502 1382 4505 1388
rect 4474 1368 4478 1371
rect 4342 1352 4345 1358
rect 4486 1352 4489 1368
rect 4510 1362 4513 1368
rect 4498 1358 4502 1361
rect 4410 1348 4414 1351
rect 4350 1332 4353 1348
rect 4486 1332 4489 1348
rect 4526 1341 4529 1498
rect 4534 1492 4537 1548
rect 4542 1542 4545 1548
rect 4582 1542 4585 1548
rect 4590 1542 4593 1658
rect 4606 1642 4609 1668
rect 4618 1658 4622 1661
rect 4638 1652 4641 1658
rect 4622 1642 4625 1648
rect 4598 1562 4601 1568
rect 4630 1541 4633 1618
rect 4646 1572 4649 1718
rect 4662 1692 4665 1748
rect 4678 1742 4681 1758
rect 4694 1742 4697 1778
rect 4710 1772 4713 1798
rect 4702 1762 4705 1768
rect 4718 1752 4721 1798
rect 4742 1792 4745 1818
rect 4742 1772 4745 1778
rect 4750 1762 4753 1768
rect 4766 1762 4769 1768
rect 4810 1758 4814 1761
rect 4826 1758 4830 1761
rect 4726 1742 4729 1758
rect 4734 1752 4737 1758
rect 4746 1748 4750 1751
rect 4810 1748 4814 1751
rect 4826 1748 4830 1751
rect 4766 1742 4769 1748
rect 4662 1662 4665 1668
rect 4670 1652 4673 1738
rect 4678 1682 4681 1718
rect 4682 1658 4686 1661
rect 4682 1648 4686 1651
rect 4654 1622 4657 1638
rect 4678 1632 4681 1648
rect 4694 1592 4697 1638
rect 4658 1588 4662 1591
rect 4702 1572 4705 1718
rect 4798 1692 4801 1738
rect 4838 1731 4841 1858
rect 4950 1822 4953 1868
rect 5070 1862 5073 1868
rect 5126 1862 5129 1868
rect 5134 1852 5137 1858
rect 4910 1792 4913 1798
rect 4878 1772 4881 1778
rect 4858 1768 4862 1771
rect 4890 1768 4894 1771
rect 4922 1768 4926 1771
rect 4898 1758 4902 1761
rect 4846 1742 4849 1748
rect 4834 1728 4841 1731
rect 4854 1732 4857 1758
rect 4942 1752 4945 1768
rect 5014 1762 5017 1768
rect 4906 1748 4910 1751
rect 4930 1748 4934 1751
rect 4818 1688 4822 1691
rect 4838 1682 4841 1728
rect 4878 1692 4881 1748
rect 4942 1742 4945 1748
rect 4762 1678 4766 1681
rect 4714 1668 4718 1671
rect 4722 1658 4726 1661
rect 4750 1652 4753 1678
rect 4806 1672 4809 1678
rect 4830 1670 4833 1678
rect 4838 1672 4841 1678
rect 4870 1672 4873 1678
rect 4886 1672 4889 1738
rect 4958 1732 4961 1758
rect 5046 1752 5049 1808
rect 5070 1752 5073 1758
rect 4970 1748 4974 1751
rect 5010 1738 5014 1741
rect 4950 1722 4953 1728
rect 5006 1712 5009 1728
rect 4952 1703 4954 1707
rect 4958 1703 4961 1707
rect 4965 1703 4968 1707
rect 4950 1672 4953 1688
rect 4990 1672 4993 1688
rect 5006 1682 5009 1708
rect 5038 1692 5041 1708
rect 5046 1692 5049 1748
rect 5094 1742 5097 1818
rect 5142 1812 5145 1948
rect 5158 1832 5161 1878
rect 5166 1872 5169 1888
rect 5198 1882 5201 1948
rect 5218 1938 5222 1941
rect 5206 1862 5209 1918
rect 5230 1892 5233 2038
rect 5254 1992 5257 2048
rect 5262 1992 5265 2208
rect 5270 2171 5273 2288
rect 5278 2272 5281 2278
rect 5282 2258 5286 2261
rect 5278 2212 5281 2248
rect 5278 2182 5281 2188
rect 5270 2168 5281 2171
rect 5270 2051 5273 2158
rect 5278 2092 5281 2168
rect 5286 2152 5289 2158
rect 5294 2132 5297 2338
rect 5302 2292 5305 2328
rect 5302 2192 5305 2278
rect 5302 2152 5305 2158
rect 5306 2138 5310 2141
rect 5286 2101 5289 2118
rect 5286 2098 5297 2101
rect 5278 2079 5286 2081
rect 5278 2078 5289 2079
rect 5278 2062 5281 2078
rect 5294 2051 5297 2098
rect 5270 2048 5281 2051
rect 5266 1968 5270 1971
rect 5238 1944 5241 1958
rect 5266 1948 5270 1951
rect 5238 1892 5241 1940
rect 5214 1872 5217 1878
rect 5262 1871 5265 1918
rect 5254 1868 5265 1871
rect 5194 1858 5198 1861
rect 5234 1858 5238 1861
rect 5246 1852 5249 1868
rect 5182 1842 5185 1848
rect 5226 1838 5230 1841
rect 5214 1772 5217 1818
rect 5218 1758 5222 1761
rect 5238 1752 5241 1758
rect 5110 1742 5113 1748
rect 5242 1738 5246 1741
rect 4758 1662 4761 1668
rect 4782 1662 4785 1668
rect 4774 1652 4777 1658
rect 4626 1538 4633 1541
rect 4686 1542 4689 1548
rect 4542 1492 4545 1528
rect 4546 1478 4553 1481
rect 4550 1472 4553 1478
rect 4566 1472 4569 1488
rect 4574 1482 4577 1508
rect 4586 1478 4590 1481
rect 4598 1472 4601 1508
rect 4542 1462 4545 1468
rect 4582 1462 4585 1468
rect 4606 1462 4609 1488
rect 4614 1472 4617 1528
rect 4630 1522 4633 1528
rect 4694 1472 4697 1518
rect 4702 1492 4705 1568
rect 4718 1562 4721 1618
rect 4742 1572 4745 1618
rect 4750 1562 4753 1648
rect 4790 1592 4793 1618
rect 4798 1592 4801 1658
rect 4806 1602 4809 1668
rect 4846 1652 4849 1658
rect 4886 1652 4889 1668
rect 4758 1562 4761 1578
rect 4802 1568 4806 1571
rect 4766 1562 4769 1568
rect 4782 1562 4785 1568
rect 4798 1562 4801 1568
rect 4814 1562 4817 1588
rect 4738 1558 4742 1561
rect 4710 1552 4713 1558
rect 4762 1548 4766 1551
rect 4794 1548 4798 1551
rect 4710 1502 4713 1548
rect 4814 1542 4817 1548
rect 4822 1542 4825 1598
rect 4886 1542 4889 1638
rect 4894 1562 4897 1568
rect 4826 1538 4830 1541
rect 4838 1531 4841 1538
rect 4830 1528 4841 1531
rect 4734 1512 4737 1518
rect 4830 1492 4833 1528
rect 4858 1518 4862 1521
rect 4662 1462 4665 1468
rect 4694 1462 4697 1468
rect 4750 1462 4753 1478
rect 4766 1462 4769 1488
rect 4850 1478 4854 1481
rect 4890 1478 4894 1481
rect 4806 1472 4809 1478
rect 4814 1472 4817 1478
rect 4830 1468 4838 1471
rect 4774 1462 4777 1468
rect 4782 1462 4785 1468
rect 4674 1458 4678 1461
rect 4790 1452 4793 1458
rect 4818 1448 4822 1451
rect 4642 1438 4646 1441
rect 4558 1392 4561 1438
rect 4798 1432 4801 1448
rect 4830 1432 4833 1468
rect 4846 1452 4849 1468
rect 4886 1452 4889 1468
rect 4894 1462 4897 1468
rect 4838 1448 4846 1451
rect 4902 1451 4905 1668
rect 4918 1663 4921 1668
rect 4942 1592 4945 1668
rect 4910 1542 4913 1588
rect 4918 1542 4921 1558
rect 4918 1532 4921 1538
rect 4926 1532 4929 1538
rect 4922 1478 4926 1481
rect 4914 1468 4918 1471
rect 4934 1461 4937 1578
rect 5014 1572 5017 1618
rect 5070 1571 5073 1668
rect 5078 1652 5081 1688
rect 5102 1672 5105 1718
rect 5110 1682 5113 1688
rect 5098 1658 5102 1661
rect 5066 1568 5073 1571
rect 4974 1562 4977 1568
rect 5030 1542 5033 1558
rect 5038 1552 5041 1568
rect 5062 1562 5065 1568
rect 5058 1548 5062 1551
rect 5010 1538 5014 1541
rect 5058 1538 5062 1541
rect 4990 1532 4994 1535
rect 4942 1492 4945 1518
rect 4952 1503 4954 1507
rect 4958 1503 4961 1507
rect 4965 1503 4968 1507
rect 4946 1468 4950 1471
rect 4930 1458 4937 1461
rect 4974 1462 4977 1468
rect 4902 1448 4913 1451
rect 4650 1368 4654 1371
rect 4726 1371 4729 1418
rect 4822 1392 4825 1428
rect 4726 1368 4737 1371
rect 4762 1368 4766 1371
rect 4594 1358 4598 1361
rect 4550 1352 4553 1358
rect 4526 1338 4534 1341
rect 4570 1338 4574 1341
rect 4598 1332 4601 1358
rect 4626 1348 4630 1351
rect 4678 1342 4681 1368
rect 4702 1362 4705 1368
rect 4686 1342 4689 1348
rect 4734 1342 4737 1368
rect 4838 1362 4841 1448
rect 4846 1392 4849 1428
rect 4854 1372 4857 1388
rect 4842 1358 4846 1361
rect 4606 1332 4609 1338
rect 4326 1328 4334 1331
rect 4514 1328 4518 1331
rect 4322 1288 4326 1291
rect 4270 1262 4273 1268
rect 4234 1168 4238 1171
rect 4166 1162 4169 1168
rect 4210 1148 4214 1151
rect 4222 1142 4225 1158
rect 4234 1148 4238 1151
rect 4186 1138 4190 1141
rect 4126 1092 4129 1118
rect 3982 992 3985 1068
rect 4006 1042 4009 1068
rect 4082 1058 4086 1061
rect 4026 1038 4030 1041
rect 3990 1012 3993 1018
rect 3990 972 3993 988
rect 3898 948 3902 951
rect 3962 948 3966 951
rect 3878 932 3881 948
rect 3890 938 3894 941
rect 3954 938 3958 941
rect 3738 878 3742 881
rect 3878 881 3881 928
rect 3870 878 3881 881
rect 3946 918 3950 921
rect 3886 881 3889 918
rect 3928 903 3930 907
rect 3934 903 3937 907
rect 3941 903 3944 907
rect 3886 878 3897 881
rect 3694 872 3697 878
rect 3718 872 3721 878
rect 3666 858 3670 861
rect 3558 762 3561 768
rect 3574 742 3577 818
rect 3614 792 3617 808
rect 3638 802 3641 858
rect 3694 852 3697 858
rect 3682 848 3686 851
rect 3694 772 3697 828
rect 3702 762 3705 818
rect 3726 792 3729 798
rect 3734 792 3737 878
rect 3870 872 3873 878
rect 3770 868 3774 871
rect 3850 868 3854 871
rect 3882 868 3886 871
rect 3786 858 3790 861
rect 3858 858 3862 861
rect 3894 861 3897 878
rect 3890 858 3897 861
rect 3914 858 3918 861
rect 3838 842 3841 858
rect 3958 852 3961 938
rect 3966 902 3969 948
rect 3974 942 3977 958
rect 3982 952 3985 968
rect 4022 962 4025 968
rect 4042 948 4046 951
rect 4062 942 4065 1008
rect 4002 938 4006 941
rect 4090 938 4094 941
rect 4030 932 4033 938
rect 4050 928 4054 931
rect 3966 862 3969 888
rect 4038 882 4041 888
rect 4050 878 4054 881
rect 3990 863 3993 878
rect 4034 868 4038 871
rect 4050 868 4054 871
rect 4022 862 4025 868
rect 4070 862 4073 868
rect 3854 842 3857 848
rect 3930 838 3934 841
rect 3718 762 3721 788
rect 3822 772 3825 818
rect 3966 792 3969 858
rect 4078 852 4081 898
rect 4110 892 4113 1058
rect 4118 952 4121 978
rect 4134 972 4137 1138
rect 4206 1132 4209 1138
rect 4230 1132 4233 1138
rect 4186 1128 4190 1131
rect 4214 1092 4217 1098
rect 4246 1092 4249 1258
rect 4254 1192 4257 1258
rect 4262 1181 4265 1258
rect 4254 1178 4265 1181
rect 4150 1052 4153 1059
rect 4182 992 4185 1048
rect 4142 942 4145 988
rect 4150 952 4153 958
rect 4170 948 4174 951
rect 4122 938 4126 941
rect 4178 938 4182 941
rect 4134 932 4137 938
rect 4206 932 4209 1088
rect 4238 1082 4241 1088
rect 4238 1062 4241 1068
rect 4222 1052 4225 1058
rect 4254 982 4257 1178
rect 4262 1152 4265 1158
rect 4262 1132 4265 1138
rect 4278 1132 4281 1268
rect 4334 1262 4337 1298
rect 4382 1292 4385 1298
rect 4350 1282 4353 1288
rect 4422 1272 4425 1328
rect 4694 1292 4697 1308
rect 4494 1272 4497 1278
rect 4638 1272 4641 1288
rect 4654 1282 4657 1288
rect 4646 1272 4649 1278
rect 4710 1272 4713 1318
rect 4742 1312 4745 1338
rect 4790 1332 4793 1338
rect 4798 1322 4801 1348
rect 4846 1342 4849 1348
rect 4830 1332 4833 1338
rect 4862 1332 4865 1448
rect 4870 1362 4873 1368
rect 4886 1342 4889 1448
rect 4910 1412 4913 1448
rect 4966 1432 4969 1438
rect 4902 1352 4905 1358
rect 4846 1292 4849 1328
rect 4870 1292 4873 1338
rect 4890 1328 4894 1331
rect 4774 1272 4777 1278
rect 4790 1272 4793 1278
rect 4362 1268 4366 1271
rect 4318 1252 4321 1258
rect 4294 1142 4297 1158
rect 4302 1152 4305 1218
rect 4310 1132 4313 1138
rect 4318 1101 4321 1178
rect 4342 1162 4345 1268
rect 4362 1258 4366 1261
rect 4430 1182 4433 1268
rect 4514 1258 4518 1261
rect 4438 1252 4441 1258
rect 4440 1203 4442 1207
rect 4446 1203 4449 1207
rect 4453 1203 4456 1207
rect 4502 1182 4505 1188
rect 4374 1152 4377 1158
rect 4338 1148 4342 1151
rect 4434 1148 4438 1151
rect 4446 1142 4449 1178
rect 4310 1098 4321 1101
rect 4310 1082 4313 1098
rect 4326 1092 4329 1128
rect 4382 1122 4385 1138
rect 4350 1082 4353 1118
rect 4438 1092 4441 1128
rect 4454 1079 4462 1081
rect 4478 1082 4481 1088
rect 4502 1082 4505 1088
rect 4542 1082 4545 1268
rect 4558 1142 4561 1228
rect 4574 1192 4577 1268
rect 4662 1262 4665 1268
rect 4718 1262 4721 1268
rect 4582 1252 4585 1258
rect 4614 1142 4617 1218
rect 4558 1122 4561 1138
rect 4566 1132 4569 1138
rect 4594 1118 4598 1121
rect 4622 1112 4625 1118
rect 4638 1092 4641 1248
rect 4750 1242 4753 1248
rect 4678 1172 4681 1188
rect 4678 1152 4681 1168
rect 4742 1151 4745 1158
rect 4690 1088 4694 1091
rect 4742 1082 4745 1128
rect 4766 1122 4769 1268
rect 4798 1252 4801 1278
rect 4830 1272 4833 1278
rect 4910 1272 4913 1408
rect 4974 1342 4977 1348
rect 4926 1332 4929 1338
rect 4946 1318 4950 1321
rect 4952 1303 4954 1307
rect 4958 1303 4961 1307
rect 4965 1303 4968 1307
rect 4982 1292 4985 1532
rect 5010 1528 5014 1531
rect 5070 1522 5073 1558
rect 5094 1552 5097 1618
rect 5126 1582 5129 1618
rect 5134 1592 5137 1718
rect 5146 1688 5150 1691
rect 5146 1678 5150 1681
rect 5126 1562 5129 1578
rect 5158 1552 5161 1728
rect 5166 1722 5169 1738
rect 5190 1692 5193 1698
rect 5174 1682 5177 1688
rect 5186 1678 5190 1681
rect 5170 1668 5174 1671
rect 5182 1662 5185 1678
rect 5198 1672 5201 1688
rect 5214 1682 5217 1688
rect 5230 1672 5233 1678
rect 5238 1672 5241 1708
rect 5254 1691 5257 1868
rect 5278 1862 5281 2048
rect 5286 2048 5297 2051
rect 5286 1962 5289 2048
rect 5294 1872 5297 1878
rect 5266 1858 5270 1861
rect 5262 1842 5265 1848
rect 5262 1742 5265 1778
rect 5270 1762 5273 1818
rect 5302 1762 5305 2088
rect 5270 1722 5273 1748
rect 5282 1728 5286 1731
rect 5246 1688 5257 1691
rect 5262 1692 5265 1708
rect 5278 1692 5281 1718
rect 5294 1702 5297 1758
rect 5290 1688 5297 1691
rect 5202 1658 5206 1661
rect 5214 1652 5217 1668
rect 5214 1602 5217 1618
rect 5222 1572 5225 1658
rect 5230 1592 5233 1668
rect 5246 1662 5249 1688
rect 5294 1672 5297 1688
rect 5174 1562 5177 1568
rect 5234 1558 5238 1561
rect 5014 1492 5017 1508
rect 5022 1481 5025 1518
rect 5078 1492 5081 1538
rect 5086 1482 5089 1548
rect 5094 1532 5097 1538
rect 5102 1522 5105 1528
rect 5110 1492 5113 1518
rect 5150 1512 5153 1538
rect 5174 1492 5177 1518
rect 5190 1502 5193 1535
rect 5206 1522 5209 1538
rect 5214 1511 5217 1558
rect 5270 1552 5273 1658
rect 5206 1508 5217 1511
rect 5206 1492 5209 1508
rect 5014 1478 5025 1481
rect 5058 1478 5062 1481
rect 5146 1478 5150 1481
rect 4990 1472 4993 1478
rect 4998 1462 5001 1468
rect 5006 1432 5009 1448
rect 4998 1392 5001 1418
rect 5014 1362 5017 1478
rect 5026 1468 5030 1471
rect 5042 1468 5046 1471
rect 5098 1468 5102 1471
rect 5030 1462 5033 1468
rect 5054 1392 5057 1468
rect 5062 1422 5065 1468
rect 5114 1458 5118 1461
rect 5102 1442 5105 1458
rect 5126 1442 5129 1458
rect 5110 1392 5113 1428
rect 5006 1342 5009 1358
rect 5034 1348 5038 1351
rect 5014 1342 5017 1348
rect 5062 1332 5065 1358
rect 5078 1348 5086 1351
rect 5050 1328 5054 1331
rect 5062 1302 5065 1328
rect 5070 1312 5073 1318
rect 5014 1272 5017 1278
rect 5010 1268 5014 1271
rect 4806 1262 4809 1268
rect 4830 1252 4833 1258
rect 4846 1252 4849 1268
rect 4786 1248 4790 1251
rect 4842 1248 4846 1251
rect 4846 1192 4849 1238
rect 4886 1192 4889 1248
rect 4902 1242 4905 1268
rect 4934 1192 4937 1268
rect 4974 1232 4977 1268
rect 5062 1262 5065 1278
rect 5078 1272 5081 1348
rect 5106 1338 5110 1341
rect 5094 1275 5097 1338
rect 5134 1332 5137 1478
rect 5142 1468 5150 1471
rect 5154 1468 5158 1471
rect 5178 1468 5182 1471
rect 5142 1462 5145 1468
rect 5154 1458 5158 1461
rect 5178 1458 5182 1461
rect 5174 1422 5177 1448
rect 5182 1362 5185 1438
rect 5182 1352 5185 1358
rect 5154 1348 5158 1351
rect 5126 1272 5129 1308
rect 5134 1272 5137 1298
rect 5142 1292 5145 1338
rect 5150 1332 5153 1338
rect 5158 1292 5161 1338
rect 5166 1292 5169 1338
rect 5182 1332 5185 1338
rect 5190 1332 5193 1478
rect 5206 1462 5209 1488
rect 5230 1472 5233 1548
rect 5242 1538 5246 1541
rect 5246 1482 5249 1528
rect 5266 1518 5270 1521
rect 5278 1492 5281 1518
rect 5294 1502 5297 1538
rect 5302 1502 5305 1758
rect 5230 1452 5233 1468
rect 5206 1362 5209 1448
rect 5218 1418 5225 1421
rect 5214 1372 5217 1378
rect 5222 1351 5225 1418
rect 5246 1392 5249 1468
rect 5238 1372 5241 1378
rect 5230 1362 5233 1368
rect 5238 1351 5241 1358
rect 5222 1348 5241 1351
rect 5198 1342 5201 1348
rect 5230 1332 5233 1348
rect 5246 1332 5249 1348
rect 5190 1292 5193 1328
rect 5222 1292 5225 1298
rect 5154 1278 5158 1281
rect 5074 1268 5078 1271
rect 5074 1258 5078 1261
rect 4994 1248 4998 1251
rect 5014 1192 5017 1218
rect 4810 1168 4814 1171
rect 4814 1132 4817 1138
rect 4838 1092 4841 1132
rect 4886 1092 4889 1148
rect 4894 1092 4897 1168
rect 4902 1152 4905 1168
rect 4986 1148 4990 1151
rect 4902 1132 4905 1148
rect 4942 1142 4945 1148
rect 5022 1141 5025 1258
rect 5066 1248 5070 1251
rect 5142 1242 5145 1278
rect 5202 1268 5206 1271
rect 5174 1262 5177 1268
rect 5186 1258 5190 1261
rect 5150 1252 5153 1258
rect 5178 1248 5182 1251
rect 5050 1238 5054 1241
rect 5062 1232 5065 1238
rect 5102 1192 5105 1208
rect 5142 1192 5145 1238
rect 5098 1168 5102 1171
rect 5114 1158 5118 1161
rect 5082 1148 5086 1151
rect 5102 1142 5105 1148
rect 5118 1142 5121 1148
rect 5126 1142 5129 1168
rect 5154 1158 5158 1161
rect 5186 1158 5190 1161
rect 5022 1138 5030 1141
rect 4910 1132 4913 1138
rect 4454 1078 4465 1079
rect 4482 1078 4494 1081
rect 4522 1078 4526 1081
rect 4358 1072 4361 1078
rect 4290 1058 4294 1061
rect 4286 992 4289 1048
rect 4318 992 4321 1018
rect 4334 992 4337 1038
rect 4342 981 4345 1068
rect 4354 1048 4358 1051
rect 4366 1051 4369 1078
rect 4406 1062 4409 1068
rect 4378 1058 4382 1061
rect 4394 1058 4398 1061
rect 4362 1048 4369 1051
rect 4382 1042 4385 1048
rect 4398 1042 4401 1048
rect 4414 1022 4417 1068
rect 4454 1062 4457 1078
rect 4422 992 4425 1048
rect 4430 1042 4433 1048
rect 4440 1003 4442 1007
rect 4446 1003 4449 1007
rect 4453 1003 4456 1007
rect 4334 978 4345 981
rect 4314 968 4318 971
rect 4214 942 4217 948
rect 4222 942 4225 948
rect 4178 928 4182 931
rect 4194 928 4198 931
rect 4126 922 4129 928
rect 4126 892 4129 898
rect 4122 878 4126 881
rect 4062 842 4065 848
rect 4086 842 4089 878
rect 4174 862 4177 918
rect 4206 882 4209 928
rect 4222 892 4225 928
rect 4250 918 4254 921
rect 4182 862 4185 868
rect 4254 862 4257 868
rect 4098 858 4102 861
rect 3738 768 3742 771
rect 3806 768 3814 771
rect 3682 758 3686 761
rect 3634 748 3638 751
rect 3522 738 3526 741
rect 3454 732 3457 738
rect 3482 728 3486 731
rect 3478 702 3481 718
rect 3574 712 3577 738
rect 3582 732 3585 738
rect 3510 662 3513 698
rect 3654 692 3657 738
rect 3662 732 3665 758
rect 3710 752 3713 758
rect 3726 752 3729 758
rect 3806 742 3809 768
rect 3834 748 3838 751
rect 3906 748 3910 751
rect 3870 741 3873 748
rect 4022 742 4025 748
rect 4030 742 4033 808
rect 4058 758 4062 761
rect 4078 742 4081 808
rect 4102 742 4105 758
rect 4150 742 4153 748
rect 4182 742 4185 858
rect 4262 832 4265 928
rect 4270 812 4273 938
rect 4302 932 4305 948
rect 4322 928 4326 931
rect 4278 862 4281 918
rect 4302 912 4305 928
rect 4334 921 4337 978
rect 4342 952 4345 958
rect 4374 942 4377 948
rect 4326 918 4337 921
rect 4366 932 4369 938
rect 4326 892 4329 918
rect 4366 892 4369 928
rect 4354 879 4361 881
rect 4350 878 4361 879
rect 4334 852 4337 868
rect 4358 862 4361 878
rect 4362 848 4366 851
rect 4318 832 4321 848
rect 4334 812 4337 848
rect 4374 842 4377 938
rect 4382 932 4385 938
rect 4398 932 4401 958
rect 4438 952 4441 958
rect 4478 952 4481 958
rect 4466 948 4470 951
rect 4438 932 4441 948
rect 4486 942 4489 1008
rect 4494 962 4497 1068
rect 4502 1062 4505 1078
rect 4550 1072 4553 1078
rect 4662 1072 4665 1078
rect 4870 1072 4873 1088
rect 4594 1068 4598 1071
rect 4518 1052 4521 1058
rect 4526 992 4529 1068
rect 4566 992 4569 1068
rect 4574 1052 4577 1058
rect 4582 992 4585 1008
rect 4598 972 4601 1058
rect 4606 1012 4609 1068
rect 4654 1042 4657 1068
rect 4538 968 4542 971
rect 4574 962 4577 968
rect 4614 962 4617 978
rect 4506 948 4510 951
rect 4494 942 4497 948
rect 4518 942 4521 948
rect 4542 922 4545 948
rect 4558 942 4561 958
rect 4614 942 4617 948
rect 4638 942 4641 988
rect 4562 938 4566 941
rect 4598 932 4601 938
rect 4646 932 4649 948
rect 4630 892 4633 928
rect 4654 882 4657 958
rect 4662 952 4665 1068
rect 4670 992 4673 1038
rect 4710 982 4713 1068
rect 4742 1063 4745 1068
rect 4862 1062 4865 1068
rect 4774 1042 4777 1058
rect 4830 992 4833 1058
rect 4890 1048 4894 1051
rect 4910 992 4913 1118
rect 4918 1082 4921 1098
rect 4942 1091 4945 1138
rect 4970 1128 4974 1131
rect 4952 1103 4954 1107
rect 4958 1103 4961 1107
rect 4965 1103 4968 1107
rect 4982 1092 4985 1138
rect 5030 1122 5033 1138
rect 5078 1121 5081 1138
rect 5074 1118 5081 1121
rect 5142 1132 5145 1158
rect 5162 1148 5166 1151
rect 4942 1088 4950 1091
rect 4990 1082 4993 1098
rect 5142 1092 5145 1128
rect 4922 1078 4929 1081
rect 4926 1072 4929 1078
rect 4990 1072 4993 1078
rect 4918 1062 4921 1068
rect 5046 1062 5049 1068
rect 5078 1063 5081 1068
rect 4938 1058 4942 1061
rect 4978 1058 4982 1061
rect 4994 1058 4998 1061
rect 5022 992 5025 1058
rect 5110 1042 5113 1058
rect 5150 1052 5153 1148
rect 5158 1092 5161 1138
rect 5166 1072 5169 1088
rect 5174 1082 5177 1158
rect 5182 1112 5185 1128
rect 5190 1072 5193 1148
rect 5198 1082 5201 1268
rect 5222 1262 5225 1278
rect 5246 1262 5249 1318
rect 5254 1302 5257 1458
rect 5262 1412 5265 1468
rect 5270 1462 5273 1468
rect 5278 1392 5281 1478
rect 5282 1368 5286 1371
rect 5266 1358 5270 1361
rect 5278 1332 5281 1348
rect 5278 1292 5281 1308
rect 5266 1268 5270 1271
rect 5206 1242 5209 1258
rect 5214 1212 5217 1248
rect 5222 1202 5225 1258
rect 5230 1222 5233 1238
rect 5246 1222 5249 1248
rect 5262 1242 5265 1248
rect 5270 1232 5273 1258
rect 5278 1242 5281 1248
rect 5206 1192 5209 1198
rect 5246 1172 5249 1178
rect 5206 1142 5209 1148
rect 5214 1111 5217 1138
rect 5238 1131 5241 1148
rect 5234 1128 5241 1131
rect 5214 1108 5225 1111
rect 5222 1092 5225 1108
rect 5262 1101 5265 1138
rect 5270 1112 5273 1128
rect 5254 1098 5265 1101
rect 5222 1072 5225 1088
rect 5198 1062 5201 1068
rect 5254 1062 5257 1098
rect 5262 1072 5265 1078
rect 5278 1072 5281 1079
rect 5282 1068 5289 1071
rect 5286 1062 5289 1068
rect 5254 1052 5257 1058
rect 5110 1021 5113 1038
rect 5110 1018 5121 1021
rect 4854 982 4857 988
rect 4670 931 4673 948
rect 4678 942 4681 948
rect 4686 942 4689 948
rect 4694 942 4697 948
rect 4710 941 4713 978
rect 5098 968 5102 971
rect 4750 962 4753 968
rect 4722 948 4726 951
rect 4710 938 4721 941
rect 4670 928 4681 931
rect 4670 892 4673 918
rect 4678 882 4681 928
rect 4702 922 4705 928
rect 4710 892 4713 928
rect 4718 902 4721 938
rect 4726 922 4729 928
rect 4734 912 4737 958
rect 4778 948 4782 951
rect 4734 892 4737 898
rect 4742 892 4745 938
rect 4766 912 4769 938
rect 4790 922 4793 958
rect 4862 942 4865 968
rect 4882 958 4886 961
rect 4946 958 4950 961
rect 4986 948 4990 951
rect 4870 942 4873 948
rect 4934 942 4937 948
rect 5046 942 5049 958
rect 5062 942 5065 948
rect 4978 938 4982 941
rect 4798 892 4801 938
rect 4846 932 4849 938
rect 4886 922 4889 938
rect 4822 892 4825 898
rect 4814 882 4817 888
rect 4482 878 4486 881
rect 4462 872 4465 878
rect 4410 868 4414 871
rect 4398 852 4401 858
rect 4390 812 4393 848
rect 4410 838 4414 841
rect 4422 822 4425 858
rect 4294 792 4297 808
rect 4366 792 4369 808
rect 4430 792 4433 828
rect 4440 803 4442 807
rect 4446 803 4449 807
rect 4453 803 4456 807
rect 4462 802 4465 868
rect 4478 862 4481 868
rect 4486 851 4489 868
rect 4514 858 4518 861
rect 4482 848 4489 851
rect 4526 852 4529 868
rect 4318 772 4321 778
rect 4290 768 4294 771
rect 4418 768 4422 771
rect 4274 758 4278 761
rect 4198 751 4201 758
rect 4282 748 4286 751
rect 3870 738 3881 741
rect 3750 721 3753 738
rect 3750 718 3758 721
rect 3774 712 3777 718
rect 3806 682 3809 688
rect 3674 679 3681 681
rect 3670 678 3681 679
rect 3394 658 3398 661
rect 3678 662 3681 678
rect 3742 672 3745 678
rect 3774 672 3777 678
rect 3782 672 3785 678
rect 3734 662 3737 668
rect 3766 662 3769 668
rect 3486 652 3489 658
rect 3574 642 3577 659
rect 3706 658 3710 661
rect 3722 658 3726 661
rect 3706 648 3710 651
rect 3690 638 3694 641
rect 3416 603 3418 607
rect 3422 603 3425 607
rect 3429 603 3432 607
rect 3574 592 3577 608
rect 3678 592 3681 638
rect 3370 588 3374 591
rect 3314 568 3318 571
rect 3238 562 3241 568
rect 3262 562 3265 568
rect 3178 558 3182 561
rect 3274 558 3278 561
rect 3170 548 3174 551
rect 3190 548 3198 551
rect 3166 521 3169 538
rect 3178 528 3182 531
rect 3162 518 3169 521
rect 3190 512 3193 548
rect 3206 542 3209 548
rect 3390 542 3393 558
rect 3510 552 3513 568
rect 3582 562 3585 588
rect 3670 572 3673 578
rect 3642 558 3646 561
rect 3198 522 3201 538
rect 3166 492 3169 508
rect 3222 502 3225 535
rect 3234 518 3238 521
rect 3262 512 3265 538
rect 3334 532 3337 538
rect 3342 512 3345 538
rect 3398 531 3401 548
rect 3486 542 3489 548
rect 3566 542 3569 548
rect 3582 542 3585 558
rect 3630 552 3633 558
rect 3638 542 3641 558
rect 3686 552 3689 618
rect 3694 592 3697 628
rect 3718 562 3721 648
rect 3750 632 3753 648
rect 3734 578 3750 581
rect 3726 572 3729 578
rect 3734 562 3737 578
rect 3766 572 3769 618
rect 3782 602 3785 658
rect 3798 652 3801 678
rect 3814 662 3817 708
rect 3862 701 3865 738
rect 3862 698 3870 701
rect 3818 658 3822 661
rect 3830 632 3833 658
rect 3838 652 3841 658
rect 3846 652 3849 658
rect 3854 642 3857 688
rect 3870 682 3873 698
rect 3878 672 3881 738
rect 3894 722 3897 738
rect 3886 682 3889 718
rect 3906 668 3910 671
rect 3918 662 3921 728
rect 3926 722 3929 728
rect 4086 722 4089 738
rect 4126 732 4129 738
rect 4134 732 4137 738
rect 3928 703 3930 707
rect 3934 703 3937 707
rect 3941 703 3944 707
rect 3966 672 3969 718
rect 4070 682 4073 688
rect 3974 672 3977 678
rect 3966 662 3969 668
rect 3938 658 3942 661
rect 3978 658 3982 661
rect 3742 562 3745 568
rect 3750 562 3753 568
rect 3654 542 3657 548
rect 3610 538 3614 541
rect 3438 532 3441 538
rect 3398 528 3406 531
rect 3390 492 3393 508
rect 3454 502 3457 518
rect 3470 482 3473 488
rect 3310 472 3313 478
rect 3414 472 3417 478
rect 3178 468 3182 471
rect 3466 468 3470 471
rect 3238 462 3241 468
rect 3246 462 3249 468
rect 3294 462 3297 468
rect 3486 462 3489 528
rect 3494 481 3497 538
rect 3494 478 3502 481
rect 3502 472 3505 478
rect 3018 458 3022 461
rect 3514 458 3518 461
rect 3530 458 3534 461
rect 2858 448 2862 451
rect 2934 442 2937 448
rect 2846 438 2857 441
rect 2890 438 2894 441
rect 2750 372 2753 378
rect 2798 372 2801 378
rect 2814 372 2817 408
rect 2854 392 2857 438
rect 2958 418 2966 421
rect 2730 368 2734 371
rect 2738 368 2742 371
rect 2826 368 2830 371
rect 2642 348 2646 351
rect 2674 348 2678 351
rect 2630 342 2633 348
rect 2606 332 2609 338
rect 2574 292 2577 318
rect 2702 312 2705 328
rect 2538 278 2542 281
rect 2550 272 2553 288
rect 2582 282 2585 288
rect 2590 282 2593 308
rect 2614 278 2617 308
rect 2654 288 2662 291
rect 2674 288 2678 291
rect 2646 272 2649 288
rect 2654 272 2657 288
rect 2702 272 2705 278
rect 2490 268 2494 271
rect 2522 268 2526 271
rect 2550 262 2553 268
rect 2434 258 2438 261
rect 2458 258 2462 261
rect 2514 258 2518 261
rect 2462 252 2465 258
rect 2710 252 2713 338
rect 2726 272 2729 328
rect 2750 302 2753 348
rect 2758 312 2761 358
rect 2782 342 2785 368
rect 2798 362 2801 368
rect 2790 342 2793 348
rect 2766 312 2769 328
rect 2806 322 2809 348
rect 2830 322 2833 358
rect 2878 352 2881 418
rect 2934 352 2937 418
rect 2842 348 2846 351
rect 2734 292 2737 298
rect 2742 272 2745 288
rect 2786 278 2790 281
rect 2766 262 2769 268
rect 2722 248 2726 251
rect 2758 242 2761 258
rect 2774 252 2777 278
rect 2814 272 2817 288
rect 2862 282 2865 298
rect 2870 282 2873 318
rect 2904 303 2906 307
rect 2910 303 2913 307
rect 2917 303 2920 307
rect 2798 262 2801 268
rect 2806 262 2809 268
rect 2830 262 2833 268
rect 2830 242 2833 248
rect 2854 242 2857 268
rect 2902 262 2905 268
rect 2910 252 2913 278
rect 2894 242 2897 248
rect 2392 203 2394 207
rect 2398 203 2401 207
rect 2405 203 2408 207
rect 2294 -18 2297 8
rect 2310 -18 2313 18
rect 486 -22 490 -18
rect 526 -22 530 -18
rect 558 -22 562 -18
rect 798 -22 802 -18
rect 1078 -22 1082 -18
rect 1110 -22 1114 -18
rect 1174 -22 1178 -18
rect 1230 -22 1234 -18
rect 1254 -22 1258 -18
rect 1278 -22 1282 -18
rect 1294 -22 1298 -18
rect 1358 -22 1362 -18
rect 1390 -22 1394 -18
rect 1462 -22 1466 -18
rect 1478 -22 1482 -18
rect 1638 -22 1642 -18
rect 1678 -22 1682 -18
rect 1734 -22 1738 -18
rect 1798 -22 1802 -18
rect 1894 -22 1898 -18
rect 1910 -22 1914 -18
rect 2006 -22 2010 -18
rect 2046 -22 2050 -18
rect 2062 -22 2066 -18
rect 2078 -22 2082 -18
rect 2094 -22 2098 -18
rect 2126 -22 2130 -18
rect 2150 -22 2154 -18
rect 2182 -22 2186 -18
rect 2198 -22 2202 -18
rect 2214 -22 2218 -18
rect 2246 -22 2250 -18
rect 2262 -22 2266 -18
rect 2278 -22 2282 -18
rect 2294 -22 2298 -18
rect 2310 -22 2314 -18
rect 2318 -19 2321 198
rect 2614 192 2617 218
rect 2630 192 2633 218
rect 2354 188 2358 191
rect 2326 152 2329 158
rect 2386 138 2390 141
rect 2334 92 2337 138
rect 2366 72 2369 98
rect 2390 72 2393 128
rect 2398 102 2401 148
rect 2430 142 2433 178
rect 2478 142 2481 148
rect 2486 142 2489 168
rect 2542 142 2545 188
rect 2558 162 2561 168
rect 2654 162 2657 188
rect 2590 142 2593 158
rect 2678 152 2681 158
rect 2686 142 2689 188
rect 2710 162 2713 218
rect 2750 192 2753 218
rect 2750 171 2753 188
rect 2746 168 2753 171
rect 2738 158 2742 161
rect 2766 152 2769 158
rect 2782 152 2785 218
rect 2878 212 2881 218
rect 2862 162 2865 168
rect 2870 162 2873 188
rect 2818 158 2822 161
rect 2714 138 2718 141
rect 2534 132 2537 138
rect 2438 72 2441 108
rect 2446 92 2449 118
rect 2462 92 2465 118
rect 2502 112 2505 118
rect 2526 82 2529 98
rect 2446 72 2449 78
rect 2494 72 2497 78
rect 2590 72 2593 88
rect 2598 72 2601 128
rect 2622 122 2625 132
rect 2702 122 2705 128
rect 2614 92 2617 118
rect 2662 112 2665 118
rect 2654 72 2657 88
rect 2694 82 2697 118
rect 2726 102 2729 148
rect 2782 142 2785 148
rect 2738 138 2742 141
rect 2754 128 2758 131
rect 2790 122 2793 138
rect 2702 92 2705 98
rect 2734 82 2737 98
rect 2670 72 2673 78
rect 2530 59 2534 62
rect 2406 42 2409 48
rect 2358 -18 2361 8
rect 2392 3 2394 7
rect 2398 3 2401 7
rect 2405 3 2408 7
rect 2446 -18 2449 8
rect 2510 -18 2513 58
rect 2646 52 2649 68
rect 2678 62 2681 68
rect 2686 62 2689 78
rect 2726 62 2729 68
rect 2670 52 2673 58
rect 2742 52 2745 98
rect 2750 92 2753 118
rect 2758 72 2761 78
rect 2758 52 2761 58
rect 2774 42 2777 108
rect 2798 101 2801 158
rect 2902 152 2905 218
rect 2814 142 2817 148
rect 2822 122 2825 138
rect 2830 132 2833 138
rect 2838 132 2841 138
rect 2846 122 2849 148
rect 2862 142 2865 148
rect 2870 132 2873 138
rect 2794 98 2801 101
rect 2782 62 2785 78
rect 2790 52 2793 98
rect 2838 88 2857 91
rect 2798 72 2801 78
rect 2806 72 2809 78
rect 2838 72 2841 88
rect 2846 72 2849 78
rect 2854 72 2857 88
rect 2862 82 2865 98
rect 2886 92 2889 148
rect 2894 132 2897 138
rect 2918 132 2921 188
rect 2934 151 2937 348
rect 2958 332 2961 418
rect 2982 342 2985 438
rect 2998 351 3001 388
rect 3094 351 3097 458
rect 3134 352 3137 438
rect 3262 402 3265 418
rect 3334 372 3337 458
rect 3446 452 3449 458
rect 3474 448 3478 451
rect 3542 451 3545 538
rect 3586 528 3590 531
rect 3602 528 3606 531
rect 3670 522 3673 538
rect 3678 532 3681 548
rect 3702 532 3705 558
rect 3750 552 3753 558
rect 3718 532 3721 548
rect 3758 542 3761 568
rect 3770 558 3774 561
rect 3778 548 3782 551
rect 3750 538 3758 541
rect 3558 472 3561 488
rect 3574 472 3577 478
rect 3590 472 3593 478
rect 3566 462 3569 468
rect 3590 452 3593 468
rect 3614 462 3617 518
rect 3638 492 3641 518
rect 3654 472 3657 498
rect 3662 462 3665 468
rect 3670 462 3673 518
rect 3702 512 3705 528
rect 3694 472 3697 478
rect 3650 458 3654 461
rect 3682 458 3686 461
rect 3694 452 3697 468
rect 3538 448 3545 451
rect 3510 442 3513 448
rect 3526 442 3529 448
rect 3416 403 3418 407
rect 3422 403 3425 407
rect 3429 403 3432 407
rect 3094 348 3102 351
rect 3182 351 3185 368
rect 3074 318 3078 321
rect 3006 292 3009 318
rect 3062 311 3065 318
rect 3062 308 3073 311
rect 2974 272 2977 278
rect 3006 272 3009 288
rect 2950 262 2953 268
rect 3002 258 3006 261
rect 3014 252 3017 278
rect 3038 272 3041 288
rect 3046 282 3049 298
rect 3062 262 3065 298
rect 3070 292 3073 308
rect 3086 302 3089 348
rect 3166 342 3169 348
rect 3094 292 3097 338
rect 3102 332 3105 338
rect 3150 322 3153 338
rect 3254 321 3257 338
rect 3254 318 3262 321
rect 3070 282 3073 288
rect 3086 262 3089 268
rect 3094 262 3097 268
rect 3034 258 3038 261
rect 3074 258 3078 261
rect 3102 252 3105 298
rect 3118 272 3121 288
rect 3118 252 3121 258
rect 2942 242 2945 248
rect 3126 222 3129 318
rect 3142 272 3145 298
rect 3150 282 3153 298
rect 3150 272 3153 278
rect 3206 272 3209 308
rect 3246 282 3249 318
rect 3270 302 3273 318
rect 3302 302 3305 338
rect 3310 301 3313 318
rect 3310 298 3321 301
rect 3246 262 3249 278
rect 3254 272 3257 278
rect 3234 258 3238 261
rect 3158 242 3161 258
rect 3262 252 3265 258
rect 3242 248 3246 251
rect 3218 238 3222 241
rect 2950 192 2953 218
rect 2998 202 3001 218
rect 2962 158 2966 161
rect 2998 152 3001 198
rect 2934 148 2945 151
rect 2926 112 2929 148
rect 2904 103 2906 107
rect 2910 103 2913 107
rect 2917 103 2920 107
rect 2934 102 2937 138
rect 2874 78 2878 81
rect 2818 68 2822 71
rect 2830 62 2833 68
rect 2894 62 2897 68
rect 2918 62 2921 68
rect 2850 58 2854 61
rect 2698 38 2702 41
rect 2710 32 2713 38
rect 2558 -18 2561 8
rect 2926 -18 2929 8
rect 2942 -18 2945 148
rect 2962 148 2966 151
rect 2950 142 2953 148
rect 3006 142 3009 188
rect 3022 162 3025 208
rect 3030 151 3033 218
rect 3026 148 3033 151
rect 3046 142 3049 158
rect 2978 138 2982 141
rect 3018 138 3022 141
rect 2982 132 2985 138
rect 3062 132 3065 208
rect 3142 162 3145 168
rect 3078 152 3081 158
rect 3158 152 3161 238
rect 3270 222 3273 288
rect 3290 278 3294 281
rect 3302 271 3305 278
rect 3298 268 3305 271
rect 3310 262 3313 288
rect 3318 282 3321 298
rect 3326 292 3329 348
rect 3342 342 3345 378
rect 3334 332 3337 338
rect 3342 312 3345 338
rect 3390 332 3393 338
rect 3398 331 3401 348
rect 3398 328 3406 331
rect 3362 318 3366 321
rect 3430 292 3433 358
rect 3486 352 3489 438
rect 3510 392 3513 428
rect 3550 352 3553 448
rect 3574 442 3577 448
rect 3618 438 3622 441
rect 3630 432 3633 448
rect 3710 442 3713 448
rect 3562 358 3566 361
rect 3466 348 3470 351
rect 3498 348 3502 351
rect 3454 342 3457 348
rect 3542 342 3545 348
rect 3318 272 3321 278
rect 3318 251 3321 258
rect 3342 252 3345 258
rect 3310 248 3321 251
rect 3310 242 3313 248
rect 3326 242 3329 248
rect 3194 168 3198 171
rect 3138 148 3142 151
rect 3074 138 3078 141
rect 3106 138 3110 141
rect 2990 122 2993 128
rect 3074 118 3078 121
rect 2974 82 2977 118
rect 2998 72 3001 118
rect 3118 112 3121 128
rect 3034 88 3038 91
rect 2990 62 2993 68
rect 2970 58 2974 61
rect 2982 42 2985 48
rect 3014 42 3017 68
rect 3070 52 3073 88
rect 3094 72 3097 78
rect 3086 52 3089 58
rect 3118 52 3121 58
rect 3126 52 3129 108
rect 3174 102 3177 148
rect 3222 142 3225 168
rect 3230 162 3233 218
rect 3234 148 3238 151
rect 3250 148 3254 151
rect 3230 132 3233 138
rect 3150 82 3153 98
rect 3198 92 3201 132
rect 3246 122 3249 128
rect 3254 102 3257 128
rect 3174 82 3177 88
rect 3214 82 3217 98
rect 3222 88 3230 91
rect 3202 78 3206 81
rect 3222 72 3225 88
rect 3270 72 3273 218
rect 3278 192 3281 218
rect 3350 202 3353 248
rect 3358 242 3361 258
rect 3382 252 3385 268
rect 3390 262 3393 268
rect 3366 242 3369 248
rect 3398 242 3401 278
rect 3438 272 3441 318
rect 3454 312 3457 338
rect 3462 332 3465 338
rect 3530 328 3534 331
rect 3478 322 3481 328
rect 3538 318 3542 321
rect 3438 262 3441 268
rect 3430 252 3433 258
rect 3390 232 3393 238
rect 3438 232 3441 248
rect 3446 242 3449 278
rect 3474 268 3478 271
rect 3462 262 3465 268
rect 3486 262 3489 278
rect 3494 272 3497 278
rect 3510 272 3513 288
rect 3518 282 3521 308
rect 3558 302 3561 358
rect 3566 332 3569 338
rect 3582 332 3585 358
rect 3606 352 3609 418
rect 3646 372 3649 418
rect 3718 372 3721 518
rect 3726 482 3729 488
rect 3750 472 3753 538
rect 3774 512 3777 548
rect 3790 542 3793 568
rect 3798 542 3801 548
rect 3806 542 3809 548
rect 3822 532 3825 618
rect 3830 562 3833 598
rect 3846 592 3849 618
rect 3886 592 3889 648
rect 3894 642 3897 648
rect 3906 638 3910 641
rect 3854 582 3857 588
rect 3830 552 3833 558
rect 3846 542 3849 578
rect 3894 572 3897 588
rect 3902 572 3905 638
rect 3918 572 3921 658
rect 3950 652 3953 658
rect 3990 652 3993 678
rect 3998 672 4001 678
rect 4006 662 4009 668
rect 4042 658 4046 661
rect 4062 652 4065 678
rect 4018 648 4022 651
rect 3870 542 3873 548
rect 3830 532 3833 538
rect 3878 532 3881 568
rect 3914 558 3918 561
rect 3906 548 3910 551
rect 3926 542 3929 568
rect 3934 552 3937 568
rect 3958 562 3961 648
rect 4034 638 4038 641
rect 4006 632 4009 638
rect 4054 632 4057 648
rect 4078 642 4081 668
rect 4102 662 4105 718
rect 4090 658 4094 661
rect 4098 648 4102 651
rect 4110 642 4113 718
rect 4134 712 4137 728
rect 4150 692 4153 738
rect 4166 702 4169 718
rect 4182 682 4185 738
rect 4310 702 4313 768
rect 4378 758 4382 761
rect 4402 758 4406 761
rect 4442 758 4446 761
rect 4138 658 4142 661
rect 4158 652 4161 678
rect 4166 672 4169 678
rect 4170 648 4174 651
rect 4130 638 4134 641
rect 4030 622 4033 628
rect 3950 542 3953 548
rect 3958 532 3961 558
rect 3986 548 3990 551
rect 4018 548 4022 551
rect 4034 548 4038 551
rect 3822 522 3825 528
rect 3758 482 3761 508
rect 3774 492 3777 498
rect 3766 472 3769 478
rect 3798 472 3801 508
rect 3814 492 3817 518
rect 3928 503 3930 507
rect 3934 503 3937 507
rect 3941 503 3944 507
rect 3966 492 3969 528
rect 3726 462 3729 468
rect 3782 451 3785 468
rect 3790 462 3793 468
rect 3782 448 3793 451
rect 3790 392 3793 448
rect 3798 372 3801 468
rect 3846 462 3849 468
rect 3854 452 3857 488
rect 3890 468 3894 471
rect 3930 468 3934 471
rect 3906 458 3910 461
rect 3870 442 3873 448
rect 3822 392 3825 418
rect 3614 342 3617 368
rect 3822 362 3825 368
rect 3846 362 3849 388
rect 3870 362 3873 398
rect 3634 358 3638 361
rect 3650 348 3654 351
rect 3610 328 3614 331
rect 3542 292 3545 298
rect 3582 282 3585 298
rect 3598 272 3601 318
rect 3646 272 3649 318
rect 3662 282 3665 348
rect 3718 342 3721 358
rect 3726 342 3729 348
rect 3670 302 3673 338
rect 3718 331 3721 338
rect 3774 332 3777 338
rect 3718 328 3729 331
rect 3686 312 3689 318
rect 3726 292 3729 328
rect 3782 322 3785 358
rect 3794 348 3798 351
rect 3866 348 3870 351
rect 3818 338 3822 341
rect 3830 332 3833 348
rect 3878 342 3881 458
rect 3918 451 3921 468
rect 3934 452 3937 458
rect 3914 448 3921 451
rect 3910 442 3913 448
rect 3862 332 3865 338
rect 3746 318 3750 321
rect 3766 292 3769 318
rect 3774 282 3777 298
rect 3666 278 3670 281
rect 3782 272 3785 308
rect 3838 272 3841 308
rect 3846 302 3849 318
rect 3886 272 3889 378
rect 3902 372 3905 428
rect 3910 352 3913 388
rect 3926 362 3929 448
rect 3958 432 3961 448
rect 3966 442 3969 488
rect 3974 462 3977 508
rect 3982 482 3985 548
rect 4070 542 4073 598
rect 4078 552 4081 628
rect 4102 602 4105 618
rect 4110 572 4113 598
rect 4110 552 4113 568
rect 4046 532 4049 538
rect 3994 528 3998 531
rect 4010 528 4014 531
rect 4086 531 4089 548
rect 4134 542 4137 548
rect 4142 541 4145 618
rect 4182 572 4185 678
rect 4198 672 4201 698
rect 4230 672 4233 698
rect 4194 658 4198 661
rect 4206 652 4209 668
rect 4238 662 4241 688
rect 4254 682 4257 698
rect 4318 692 4321 748
rect 4342 732 4345 758
rect 4430 752 4433 758
rect 4394 748 4398 751
rect 4374 732 4377 738
rect 4342 692 4345 698
rect 4382 692 4385 748
rect 4402 738 4406 741
rect 4398 692 4401 738
rect 4306 688 4313 691
rect 4310 672 4313 688
rect 4366 672 4369 678
rect 4422 672 4425 698
rect 4446 672 4449 728
rect 4258 668 4262 671
rect 4418 668 4422 671
rect 4454 670 4457 778
rect 4462 732 4465 798
rect 4478 782 4481 848
rect 4534 842 4537 858
rect 4542 842 4545 878
rect 4702 872 4705 878
rect 4658 868 4662 871
rect 4718 870 4721 878
rect 4766 872 4769 878
rect 4570 858 4574 861
rect 4610 858 4614 861
rect 4630 852 4633 868
rect 4646 862 4649 868
rect 4582 842 4585 848
rect 4606 842 4609 848
rect 4622 842 4625 848
rect 4478 752 4481 778
rect 4494 762 4497 768
rect 4510 762 4513 778
rect 4542 762 4545 838
rect 4646 832 4649 858
rect 4686 822 4689 848
rect 4558 782 4561 818
rect 4566 792 4569 808
rect 4574 771 4577 818
rect 4598 781 4601 818
rect 4606 792 4609 818
rect 4694 792 4697 868
rect 4702 812 4705 868
rect 4710 822 4713 868
rect 4754 868 4758 871
rect 4778 868 4782 871
rect 4762 858 4769 861
rect 4766 792 4769 858
rect 4790 852 4793 878
rect 4814 792 4817 878
rect 4862 872 4865 878
rect 4870 872 4873 918
rect 4878 892 4881 908
rect 4934 892 4937 938
rect 4962 928 4966 931
rect 4952 903 4954 907
rect 4958 903 4961 907
rect 4965 903 4968 907
rect 4974 892 4977 918
rect 5006 892 5009 928
rect 5030 882 5033 888
rect 4830 792 4833 848
rect 4838 832 4841 858
rect 4846 852 4849 858
rect 4590 778 4601 781
rect 4674 778 4678 781
rect 4566 768 4577 771
rect 4558 762 4561 768
rect 4534 752 4537 758
rect 4566 752 4569 768
rect 4582 762 4585 768
rect 4574 752 4577 758
rect 4590 752 4593 778
rect 4602 768 4606 771
rect 4666 768 4670 771
rect 4682 768 4686 771
rect 4614 762 4617 768
rect 4490 748 4494 751
rect 4522 748 4526 751
rect 4470 742 4473 748
rect 4630 742 4633 768
rect 4638 752 4641 758
rect 4646 742 4649 758
rect 4514 738 4518 741
rect 4478 731 4481 738
rect 4470 728 4481 731
rect 4470 692 4473 728
rect 4566 692 4569 738
rect 4614 732 4617 738
rect 4618 688 4625 691
rect 4486 672 4489 678
rect 4226 658 4230 661
rect 4250 658 4254 661
rect 4314 648 4318 651
rect 4290 638 4294 641
rect 4222 632 4225 638
rect 4190 552 4193 618
rect 4334 602 4337 668
rect 4358 652 4361 668
rect 4390 652 4393 658
rect 4414 652 4417 658
rect 4430 612 4433 668
rect 4502 663 4505 688
rect 4622 672 4625 688
rect 4570 668 4574 671
rect 4646 662 4649 708
rect 4654 692 4657 748
rect 4678 692 4681 768
rect 4694 752 4697 758
rect 4730 748 4734 751
rect 4710 732 4713 738
rect 4670 672 4673 688
rect 4702 682 4705 698
rect 4710 672 4713 708
rect 4730 688 4734 691
rect 4742 682 4745 748
rect 4782 742 4785 758
rect 4790 752 4793 758
rect 4798 742 4801 778
rect 4750 692 4753 738
rect 4814 732 4817 768
rect 4846 748 4854 751
rect 4758 682 4761 698
rect 4766 672 4769 698
rect 4798 692 4801 728
rect 4814 672 4817 708
rect 4846 692 4849 748
rect 4862 722 4865 868
rect 4870 822 4873 868
rect 4894 862 4897 868
rect 4902 862 4905 868
rect 4882 848 4886 851
rect 4894 842 4897 858
rect 4918 852 4921 858
rect 4906 848 4910 851
rect 4926 842 4929 868
rect 4934 862 4937 868
rect 4950 832 4953 848
rect 4990 842 4993 868
rect 5014 862 5017 868
rect 5030 852 5033 858
rect 5002 848 5006 851
rect 4950 772 4953 828
rect 4982 792 4985 818
rect 5014 792 5017 848
rect 5038 842 5041 938
rect 5046 932 5049 938
rect 5070 932 5073 938
rect 5118 922 5121 1018
rect 5194 948 5198 951
rect 5126 942 5129 948
rect 5110 892 5113 918
rect 5142 892 5145 928
rect 5174 922 5177 948
rect 5150 878 5153 908
rect 5222 892 5225 1018
rect 5238 952 5241 968
rect 5258 958 5262 961
rect 5262 932 5265 938
rect 5270 892 5273 1008
rect 5278 942 5281 948
rect 5286 892 5289 948
rect 5182 888 5190 891
rect 5202 888 5206 891
rect 5174 872 5177 888
rect 5182 872 5185 888
rect 5262 882 5265 888
rect 5250 879 5257 881
rect 5246 878 5257 879
rect 5050 868 5054 871
rect 5030 792 5033 838
rect 4974 762 4977 768
rect 4930 748 4934 751
rect 4870 732 4873 738
rect 4854 682 4857 698
rect 4622 652 4625 658
rect 4654 642 4657 648
rect 4694 642 4697 668
rect 4862 662 4865 668
rect 4886 662 4889 748
rect 4910 742 4913 748
rect 4946 738 4950 741
rect 4902 712 4905 728
rect 4950 721 4953 728
rect 4942 718 4953 721
rect 4926 692 4929 718
rect 4902 672 4905 688
rect 4942 682 4945 718
rect 4952 703 4954 707
rect 4958 703 4961 707
rect 4965 703 4968 707
rect 4974 692 4977 758
rect 4982 752 4985 758
rect 4990 692 4993 768
rect 5002 758 5006 761
rect 5014 752 5017 788
rect 5022 772 5025 778
rect 5038 732 5041 748
rect 5046 712 5049 718
rect 5054 712 5057 728
rect 4910 662 4913 668
rect 4826 658 4830 661
rect 4718 642 4721 658
rect 4742 642 4745 658
rect 4886 652 4889 658
rect 4918 652 4921 668
rect 4942 662 4945 678
rect 5030 672 5033 708
rect 5042 678 5046 681
rect 5062 671 5065 718
rect 5058 668 5065 671
rect 5070 672 5073 858
rect 5110 782 5113 818
rect 5230 802 5233 868
rect 5254 862 5257 878
rect 5274 868 5278 871
rect 5282 858 5286 861
rect 5262 792 5265 858
rect 5130 788 5134 791
rect 5138 768 5142 771
rect 5126 762 5129 768
rect 5150 762 5153 768
rect 5106 758 5110 761
rect 5078 752 5081 758
rect 5078 732 5081 748
rect 5110 742 5113 748
rect 5094 722 5097 738
rect 5086 682 5089 688
rect 5118 682 5121 748
rect 5126 742 5129 748
rect 5098 678 5102 681
rect 4974 662 4977 668
rect 5022 662 5025 668
rect 5158 662 5161 718
rect 5166 682 5169 768
rect 5182 752 5185 778
rect 5202 748 5206 751
rect 5246 732 5249 738
rect 5202 688 5206 691
rect 5230 662 5233 668
rect 5254 662 5257 678
rect 4982 652 4985 658
rect 4878 642 4881 648
rect 4966 642 4969 648
rect 5102 642 5105 658
rect 4440 603 4442 607
rect 4446 603 4449 607
rect 4453 603 4456 607
rect 4378 568 4385 571
rect 4162 548 4166 551
rect 4274 548 4278 551
rect 4314 548 4318 551
rect 4354 548 4358 551
rect 4142 538 4150 541
rect 4086 528 4094 531
rect 4006 502 4009 528
rect 4054 522 4057 528
rect 4138 528 4142 531
rect 4170 528 4174 531
rect 4042 518 4046 521
rect 3990 482 3993 498
rect 3998 482 4001 488
rect 4046 472 4049 488
rect 4054 472 4057 478
rect 3974 452 3977 458
rect 4006 452 4009 468
rect 4014 442 4017 458
rect 3978 438 3982 441
rect 3974 352 3977 368
rect 4006 352 4009 358
rect 3978 338 3982 341
rect 3990 332 3993 348
rect 3998 332 4001 338
rect 4014 322 4017 438
rect 4022 402 4025 468
rect 4054 462 4057 468
rect 4070 462 4073 488
rect 4102 472 4105 488
rect 4110 482 4113 498
rect 4134 492 4137 528
rect 4094 462 4097 468
rect 4082 458 4086 461
rect 4126 452 4129 468
rect 4134 462 4137 468
rect 4142 452 4145 498
rect 4190 472 4193 538
rect 4198 532 4201 548
rect 4262 542 4265 548
rect 4210 538 4214 541
rect 4270 532 4273 538
rect 4278 532 4281 538
rect 4302 532 4305 548
rect 4382 542 4385 568
rect 4414 568 4422 571
rect 4222 502 4225 528
rect 4246 512 4249 518
rect 4294 512 4297 528
rect 4326 522 4329 538
rect 4334 522 4337 538
rect 4338 518 4342 521
rect 4390 502 4393 548
rect 4414 542 4417 568
rect 4462 542 4465 608
rect 5270 592 5273 618
rect 4546 568 4550 571
rect 4518 562 4521 568
rect 4566 562 4569 568
rect 4522 548 4526 551
rect 4494 531 4497 538
rect 4490 528 4497 531
rect 4198 482 4201 498
rect 4222 472 4225 488
rect 4242 479 4249 481
rect 4238 478 4249 479
rect 4154 458 4158 461
rect 4206 452 4209 468
rect 4246 462 4249 478
rect 4438 472 4441 478
rect 4446 472 4449 518
rect 4486 512 4489 528
rect 4518 522 4521 538
rect 4534 502 4537 558
rect 4554 548 4558 551
rect 4590 542 4593 548
rect 4598 532 4601 568
rect 4626 548 4630 551
rect 4674 548 4678 551
rect 4698 548 4702 551
rect 4638 542 4641 548
rect 4726 541 4729 548
rect 4726 538 4734 541
rect 4750 541 4753 548
rect 4746 538 4753 541
rect 4606 532 4609 538
rect 4650 528 4654 531
rect 4482 478 4486 481
rect 4218 458 4222 461
rect 4062 442 4065 448
rect 4078 392 4081 448
rect 4174 442 4177 448
rect 4162 438 4166 441
rect 4150 432 4153 438
rect 4270 422 4273 458
rect 4278 412 4281 458
rect 4302 452 4305 468
rect 4358 442 4361 468
rect 4382 462 4385 468
rect 4446 452 4449 468
rect 4502 462 4505 488
rect 4518 472 4521 478
rect 4534 472 4537 488
rect 4378 448 4382 451
rect 4454 442 4457 458
rect 4494 442 4497 458
rect 4518 452 4521 458
rect 4550 452 4553 498
rect 4558 462 4561 518
rect 4590 512 4593 528
rect 4614 492 4617 518
rect 4662 492 4665 518
rect 4734 502 4737 538
rect 4590 462 4593 478
rect 4602 468 4606 471
rect 4574 452 4577 458
rect 4550 442 4553 448
rect 4566 442 4569 448
rect 4322 418 4326 421
rect 4390 392 4393 438
rect 4406 412 4409 418
rect 4440 403 4442 407
rect 4446 403 4449 407
rect 4453 403 4456 407
rect 4166 368 4174 371
rect 4022 342 4025 348
rect 4030 342 4033 368
rect 4086 362 4089 368
rect 4034 338 4038 341
rect 3986 318 3990 321
rect 4038 312 4041 328
rect 4054 322 4057 348
rect 4062 342 4065 348
rect 4078 322 4081 348
rect 4166 342 4169 368
rect 4214 342 4217 388
rect 4426 378 4430 381
rect 4266 368 4273 371
rect 4322 368 4329 371
rect 4242 348 4246 351
rect 4270 342 4273 368
rect 4278 342 4281 348
rect 4326 342 4329 368
rect 4382 342 4385 368
rect 4406 342 4409 348
rect 4454 342 4457 378
rect 4478 362 4481 418
rect 4502 382 4505 418
rect 4498 368 4502 371
rect 4514 358 4518 361
rect 4526 352 4529 378
rect 4542 362 4545 398
rect 4506 348 4510 351
rect 4486 342 4489 348
rect 4542 342 4545 348
rect 4558 342 4561 418
rect 4582 362 4585 458
rect 4602 448 4606 451
rect 4614 442 4617 458
rect 4622 442 4625 488
rect 4638 462 4641 488
rect 4654 462 4657 478
rect 4666 468 4670 471
rect 4666 458 4670 461
rect 4638 452 4641 458
rect 4566 342 4569 358
rect 4598 352 4601 378
rect 4614 371 4617 418
rect 4646 402 4649 458
rect 4678 452 4681 468
rect 4614 368 4625 371
rect 4610 358 4614 361
rect 4622 342 4625 368
rect 4638 352 4641 378
rect 4570 338 4574 341
rect 3928 303 3930 307
rect 3934 303 3937 307
rect 3941 303 3944 307
rect 4086 302 4089 338
rect 4102 332 4105 338
rect 4006 292 4009 298
rect 4110 291 4113 338
rect 4106 288 4113 291
rect 4138 318 4142 321
rect 4222 321 4225 338
rect 4334 332 4337 338
rect 4222 318 4230 321
rect 4354 318 4358 321
rect 4102 272 4105 288
rect 4118 272 4121 318
rect 4182 312 4185 318
rect 4134 292 4137 298
rect 4182 282 4185 298
rect 4210 288 4214 291
rect 4250 288 4254 291
rect 4294 282 4297 318
rect 4182 272 4185 278
rect 3578 268 3582 271
rect 3634 268 3638 271
rect 3722 268 3726 271
rect 4002 268 4006 271
rect 4170 268 4174 271
rect 4242 268 4246 271
rect 3526 252 3529 268
rect 3670 262 3673 268
rect 3750 262 3753 268
rect 3758 262 3761 268
rect 3830 262 3833 268
rect 3866 258 3870 261
rect 3938 258 3942 261
rect 4106 258 4110 261
rect 3646 252 3649 258
rect 3726 252 3729 258
rect 3626 248 3630 251
rect 3750 241 3753 258
rect 3814 252 3817 258
rect 3910 242 3913 258
rect 4038 252 4041 258
rect 3750 238 3761 241
rect 3358 171 3361 218
rect 3416 203 3418 207
rect 3422 203 3425 207
rect 3429 203 3432 207
rect 3350 168 3361 171
rect 3310 162 3313 168
rect 3326 162 3329 168
rect 3278 112 3281 158
rect 3350 152 3353 168
rect 3362 158 3366 161
rect 3458 158 3462 161
rect 3302 82 3305 148
rect 3350 142 3353 148
rect 3358 142 3361 158
rect 3406 142 3409 158
rect 3486 152 3489 218
rect 3570 168 3574 171
rect 3438 142 3441 148
rect 3486 142 3489 148
rect 3526 142 3529 168
rect 3622 162 3625 188
rect 3638 172 3641 188
rect 3686 182 3689 218
rect 3654 162 3657 168
rect 3710 162 3713 168
rect 3570 158 3574 161
rect 3698 158 3702 161
rect 3378 138 3382 141
rect 3522 138 3526 141
rect 3310 92 3313 138
rect 3326 122 3329 138
rect 3462 132 3465 138
rect 3370 128 3374 131
rect 3386 128 3390 131
rect 3402 128 3406 131
rect 3390 102 3393 128
rect 3382 92 3385 98
rect 3290 78 3294 81
rect 3154 68 3158 71
rect 3134 62 3137 68
rect 3174 62 3177 68
rect 3190 62 3193 68
rect 3278 62 3281 78
rect 3358 72 3361 78
rect 3366 72 3369 78
rect 3322 68 3326 71
rect 3418 68 3422 71
rect 3218 58 3222 61
rect 3002 38 3006 41
rect 3138 38 3142 41
rect 3286 32 3289 68
rect 3326 52 3329 68
rect 3342 62 3345 68
rect 3430 62 3433 98
rect 3438 72 3441 88
rect 3454 82 3457 118
rect 3462 72 3465 128
rect 3470 122 3473 128
rect 3478 122 3481 138
rect 3558 132 3561 138
rect 3582 132 3585 148
rect 3590 142 3593 158
rect 3598 132 3601 158
rect 3630 152 3633 158
rect 3698 148 3702 151
rect 3638 142 3641 148
rect 3654 142 3657 148
rect 3710 142 3713 148
rect 3618 138 3622 141
rect 3490 128 3494 131
rect 3522 128 3526 131
rect 3562 128 3569 131
rect 3534 122 3537 128
rect 3502 112 3505 118
rect 3502 92 3505 108
rect 3526 72 3529 78
rect 3462 52 3465 68
rect 3550 62 3553 68
rect 3566 52 3569 128
rect 3686 122 3689 138
rect 3718 132 3721 218
rect 3758 192 3761 238
rect 3786 188 3790 191
rect 3742 172 3745 178
rect 3746 168 3750 171
rect 3734 142 3737 148
rect 3742 132 3745 158
rect 3766 142 3769 178
rect 3794 168 3798 171
rect 3818 168 3822 171
rect 3774 162 3777 168
rect 3826 158 3830 161
rect 3886 152 3889 228
rect 3946 178 3950 181
rect 3786 148 3790 151
rect 3822 142 3825 148
rect 3602 118 3606 121
rect 3718 102 3721 128
rect 3774 92 3777 118
rect 3574 72 3577 78
rect 3606 62 3609 88
rect 3630 82 3633 88
rect 3646 82 3649 88
rect 3614 72 3617 78
rect 3626 68 3630 71
rect 3650 68 3654 71
rect 3662 62 3665 78
rect 3706 68 3710 71
rect 3642 58 3646 61
rect 3698 58 3702 61
rect 3590 52 3593 58
rect 3598 52 3601 58
rect 3306 48 3310 51
rect 3350 42 3353 48
rect 3678 42 3681 48
rect 3702 42 3705 48
rect 3718 42 3721 78
rect 3758 72 3761 78
rect 3730 68 3734 71
rect 3734 42 3737 48
rect 3742 42 3745 58
rect 3766 52 3769 78
rect 3782 70 3785 138
rect 3822 122 3825 128
rect 3798 72 3801 98
rect 3822 92 3825 118
rect 3886 92 3889 138
rect 3810 88 3814 91
rect 3822 72 3825 78
rect 3846 72 3849 88
rect 3874 78 3878 81
rect 3786 66 3790 69
rect 3822 52 3825 58
rect 3854 52 3857 78
rect 3886 52 3889 58
rect 3754 48 3758 51
rect 3810 48 3814 51
rect 3874 48 3878 51
rect 3490 38 3494 41
rect 3006 22 3009 28
rect 3902 12 3905 147
rect 3918 132 3921 138
rect 3982 132 3985 138
rect 3910 82 3913 98
rect 3918 72 3921 118
rect 3928 103 3930 107
rect 3934 103 3937 107
rect 3941 103 3944 107
rect 3938 88 3942 91
rect 3918 62 3921 68
rect 3958 62 3961 108
rect 3982 92 3985 98
rect 2982 -18 2985 8
rect 3006 -18 3009 8
rect 3086 -18 3089 8
rect 3182 -18 3185 8
rect 3342 -18 3345 8
rect 3416 3 3418 7
rect 3422 3 3425 7
rect 3429 3 3432 7
rect 3502 -18 3505 8
rect 3558 -18 3561 8
rect 3718 -18 3721 8
rect 3878 -18 3881 8
rect 3990 -18 3993 148
rect 4046 131 4049 148
rect 4054 142 4057 258
rect 4118 252 4121 268
rect 4130 258 4134 261
rect 4246 252 4249 258
rect 4294 252 4297 278
rect 4274 248 4278 251
rect 4094 152 4097 198
rect 4102 152 4105 248
rect 4134 192 4137 248
rect 4146 238 4158 241
rect 4302 192 4305 268
rect 4310 242 4313 318
rect 4346 288 4350 291
rect 4398 282 4401 338
rect 4534 332 4537 338
rect 4622 332 4625 338
rect 4578 328 4582 331
rect 4510 322 4513 328
rect 4614 292 4617 318
rect 4578 279 4585 281
rect 4574 278 4585 279
rect 4494 272 4497 278
rect 4322 258 4326 261
rect 4374 252 4377 268
rect 4462 262 4465 268
rect 4582 262 4585 278
rect 4590 272 4593 278
rect 4638 272 4641 278
rect 4646 272 4649 378
rect 4662 342 4665 348
rect 4670 332 4673 418
rect 4686 412 4689 458
rect 4694 422 4697 478
rect 4710 472 4713 488
rect 4738 478 4742 481
rect 4766 472 4769 518
rect 4774 512 4777 528
rect 4790 522 4793 548
rect 4814 532 4817 558
rect 4842 548 4846 551
rect 4854 542 4857 568
rect 4866 558 4870 561
rect 4866 548 4870 551
rect 4878 542 4881 558
rect 4890 548 4894 551
rect 5010 548 5014 551
rect 4902 542 4905 548
rect 4834 538 4838 541
rect 4954 538 4958 541
rect 4894 522 4897 538
rect 5022 532 5025 558
rect 5046 552 5049 578
rect 5078 572 5081 578
rect 5114 548 5118 551
rect 5142 551 5145 578
rect 5278 572 5281 588
rect 5174 562 5177 568
rect 5294 562 5297 1488
rect 5302 1272 5305 1278
rect 5302 1122 5305 1148
rect 5302 742 5305 868
rect 5038 522 5041 548
rect 5210 548 5214 551
rect 5238 551 5241 558
rect 4782 472 4785 518
rect 4798 482 4801 518
rect 4822 482 4825 518
rect 4862 502 4865 518
rect 4846 482 4849 488
rect 4862 481 4865 498
rect 4862 478 4870 481
rect 4702 382 4705 418
rect 4682 368 4686 371
rect 4710 362 4713 468
rect 4718 462 4721 468
rect 4790 462 4793 468
rect 4722 458 4726 461
rect 4798 452 4801 478
rect 4806 462 4809 468
rect 4746 448 4750 451
rect 4718 442 4721 448
rect 4758 432 4761 438
rect 4854 412 4857 468
rect 4862 462 4865 468
rect 4886 432 4889 468
rect 4894 462 4897 468
rect 4870 422 4873 428
rect 4902 401 4905 478
rect 4910 472 4913 508
rect 4952 503 4954 507
rect 4958 503 4961 507
rect 4965 503 4968 507
rect 5030 492 5033 518
rect 5054 501 5057 540
rect 5070 502 5073 518
rect 5050 498 5065 501
rect 4950 462 4953 468
rect 4982 462 4985 478
rect 5054 472 5057 478
rect 4958 452 4961 458
rect 4926 442 4929 448
rect 4998 442 5001 468
rect 5006 462 5009 468
rect 5030 462 5033 468
rect 5038 442 5041 448
rect 4938 438 4942 441
rect 5018 438 5022 441
rect 5046 432 5049 468
rect 5062 452 5065 498
rect 5074 478 5078 481
rect 5086 462 5089 488
rect 5094 472 5097 498
rect 5122 468 5126 471
rect 5174 462 5177 468
rect 5214 462 5217 548
rect 5282 548 5286 551
rect 5294 542 5297 558
rect 5278 482 5281 538
rect 5070 452 5073 458
rect 5130 448 5134 451
rect 5142 442 5145 458
rect 5170 448 5174 451
rect 4934 422 4937 428
rect 4902 398 4910 401
rect 4746 388 4750 391
rect 4966 382 4969 418
rect 5014 412 5017 418
rect 5054 392 5057 438
rect 5142 382 5145 418
rect 5150 392 5153 438
rect 4910 372 4913 378
rect 4938 368 4942 371
rect 4894 362 4897 368
rect 4962 358 4966 361
rect 4686 352 4689 358
rect 4694 342 4697 348
rect 4726 342 4729 348
rect 4682 338 4686 341
rect 4554 258 4558 261
rect 4162 188 4166 191
rect 4198 152 4201 158
rect 4102 142 4105 148
rect 4046 128 4054 131
rect 4014 72 4017 128
rect 4162 118 4166 121
rect 4102 63 4105 88
rect 4166 82 4169 88
rect 4214 72 4217 168
rect 4122 68 4126 71
rect 4022 -18 4025 58
rect 4046 -18 4049 8
rect 4094 -18 4097 8
rect 4118 -18 4121 58
rect 4190 -18 4193 8
rect 4214 -18 4217 58
rect 4230 -18 4233 147
rect 4310 142 4313 238
rect 4342 182 4345 188
rect 4398 172 4401 238
rect 4414 168 4422 171
rect 4338 148 4342 151
rect 4358 142 4361 148
rect 4414 142 4417 168
rect 4430 162 4433 258
rect 4440 203 4442 207
rect 4446 203 4449 207
rect 4453 203 4456 207
rect 4462 142 4465 208
rect 4502 192 4505 248
rect 4614 242 4617 258
rect 4646 252 4649 268
rect 4662 262 4665 268
rect 4662 242 4665 248
rect 4678 242 4681 288
rect 4686 262 4689 288
rect 4702 272 4705 328
rect 4710 302 4713 318
rect 4698 268 4702 271
rect 4718 271 4721 328
rect 4774 322 4777 338
rect 4782 332 4785 338
rect 4790 332 4793 348
rect 4798 342 4801 348
rect 4806 342 4809 358
rect 4862 352 4865 358
rect 4902 352 4905 358
rect 4914 348 4918 351
rect 4826 340 4830 343
rect 4838 342 4841 348
rect 4850 338 4854 341
rect 4718 268 4726 271
rect 4710 262 4713 268
rect 4726 262 4729 268
rect 4690 248 4694 251
rect 4542 142 4545 208
rect 4590 142 4593 148
rect 4598 142 4601 208
rect 4686 182 4689 218
rect 4706 168 4710 171
rect 4678 152 4681 168
rect 4718 162 4721 258
rect 4734 252 4737 278
rect 4758 272 4761 298
rect 4798 292 4801 318
rect 4794 268 4798 271
rect 4750 262 4753 268
rect 4806 262 4809 338
rect 4862 322 4865 328
rect 4814 282 4817 318
rect 4862 282 4865 318
rect 4870 312 4873 328
rect 4878 302 4881 338
rect 4926 332 4929 358
rect 4938 348 4942 351
rect 4954 348 4966 351
rect 4970 348 4974 351
rect 4982 342 4985 378
rect 5042 368 5046 371
rect 4990 342 4993 368
rect 5006 342 5009 358
rect 5018 348 5022 351
rect 4952 303 4954 307
rect 4958 303 4961 307
rect 4965 303 4968 307
rect 4870 282 4873 298
rect 4890 288 4894 291
rect 4982 282 4985 338
rect 5006 332 5009 338
rect 5014 322 5017 338
rect 4990 282 4993 288
rect 4882 278 4886 281
rect 4998 281 5001 318
rect 5030 292 5033 358
rect 5214 352 5217 458
rect 5246 452 5249 459
rect 5270 352 5273 358
rect 5050 348 5054 351
rect 5106 348 5110 351
rect 5130 348 5134 351
rect 5078 332 5081 338
rect 5110 332 5113 338
rect 5086 322 5089 328
rect 5118 322 5121 348
rect 5174 342 5177 348
rect 5142 332 5145 338
rect 4998 278 5009 281
rect 4770 258 4774 261
rect 4826 258 4830 261
rect 4838 252 4841 278
rect 4958 272 4961 278
rect 4906 268 4910 271
rect 4994 268 4998 271
rect 4778 248 4782 251
rect 4834 248 4838 251
rect 4726 242 4729 248
rect 4702 152 4705 158
rect 4726 152 4729 238
rect 4646 142 4649 148
rect 4262 122 4265 138
rect 4294 112 4297 118
rect 4326 98 4334 101
rect 4258 88 4262 91
rect 4318 82 4321 88
rect 4270 72 4273 78
rect 4302 72 4305 78
rect 4314 68 4318 71
rect 4286 62 4289 68
rect 4298 58 4302 61
rect 4326 52 4329 98
rect 4334 82 4337 98
rect 4350 92 4353 128
rect 4406 122 4409 138
rect 4374 102 4377 118
rect 4438 72 4441 108
rect 4486 72 4489 108
rect 4534 102 4537 138
rect 4618 118 4622 121
rect 4558 112 4561 118
rect 4654 102 4657 148
rect 4734 142 4737 178
rect 4758 172 4761 248
rect 4858 238 4862 241
rect 4894 232 4897 268
rect 4926 262 4929 268
rect 4906 258 4910 261
rect 4910 232 4913 248
rect 4926 242 4929 248
rect 4950 242 4953 268
rect 5006 262 5009 278
rect 5006 242 5009 258
rect 5030 242 5033 258
rect 5038 252 5041 278
rect 5062 272 5065 278
rect 5046 262 5049 268
rect 5078 262 5081 268
rect 5086 251 5089 318
rect 5134 312 5137 328
rect 5190 292 5193 328
rect 5214 302 5217 348
rect 5134 282 5137 288
rect 5182 282 5185 288
rect 5166 272 5169 278
rect 5106 268 5110 271
rect 5130 268 5134 271
rect 5154 268 5158 271
rect 5182 262 5185 278
rect 5206 262 5209 288
rect 5214 272 5217 288
rect 5222 262 5225 268
rect 5098 258 5102 261
rect 5122 258 5126 261
rect 5154 258 5158 261
rect 5082 248 5089 251
rect 5094 248 5102 251
rect 5018 238 5022 241
rect 5014 222 5017 228
rect 4766 172 4769 218
rect 5046 202 5049 248
rect 5086 232 5089 238
rect 5070 192 5073 198
rect 4878 182 4881 188
rect 4778 158 4782 161
rect 4798 152 4801 178
rect 5062 172 5065 178
rect 4850 168 4854 171
rect 5074 168 5078 171
rect 5094 162 5097 248
rect 5102 192 5105 238
rect 5134 192 5137 248
rect 5106 168 5110 171
rect 4810 158 4814 161
rect 4874 158 4878 161
rect 4922 158 4926 161
rect 4946 158 4950 161
rect 5098 158 5105 161
rect 4838 152 4841 158
rect 4778 148 4782 151
rect 4866 148 4873 151
rect 4790 142 4793 148
rect 4862 142 4865 148
rect 4682 138 4686 141
rect 4802 138 4806 141
rect 4742 132 4745 138
rect 4838 132 4841 138
rect 4706 128 4710 131
rect 4762 128 4766 131
rect 4718 122 4721 128
rect 4770 118 4774 121
rect 4494 92 4497 98
rect 4606 92 4609 98
rect 4870 92 4873 148
rect 4886 132 4889 158
rect 4894 102 4897 148
rect 4978 138 4982 141
rect 4918 132 4921 138
rect 4934 132 4937 138
rect 4952 103 4954 107
rect 4958 103 4961 107
rect 4965 103 4968 107
rect 4982 92 4985 128
rect 4990 92 4993 158
rect 5090 148 5094 151
rect 5002 138 5006 141
rect 5030 131 5033 148
rect 5102 142 5105 158
rect 5142 152 5145 158
rect 5122 148 5126 151
rect 5074 138 5078 141
rect 5030 128 5038 131
rect 5046 131 5049 138
rect 5042 128 5049 131
rect 5142 132 5145 138
rect 4998 122 5001 128
rect 5038 112 5041 128
rect 5098 108 5105 111
rect 4842 88 4849 91
rect 4922 88 4926 91
rect 5026 88 5030 91
rect 5082 88 5086 91
rect 4558 82 4561 88
rect 4558 72 4561 78
rect 4638 72 4641 88
rect 4654 72 4657 78
rect 4846 72 4849 88
rect 5006 72 5009 78
rect 5038 72 5041 88
rect 5062 72 5065 78
rect 4338 68 4342 71
rect 4414 62 4417 68
rect 4358 52 4361 58
rect 4470 52 4473 58
rect 4290 48 4294 51
rect 4386 38 4390 41
rect 4422 -18 4425 8
rect 4440 3 4442 7
rect 4446 3 4449 7
rect 4453 3 4456 7
rect 4486 -18 4489 8
rect 4534 -18 4537 58
rect 4590 41 4593 68
rect 4762 58 4766 61
rect 4590 38 4598 41
rect 4686 -18 4689 58
rect 4790 41 4793 68
rect 4798 62 4801 68
rect 4902 52 4905 68
rect 4786 38 4793 41
rect 4974 -18 4977 58
rect 5038 52 5041 58
rect 5070 52 5073 78
rect 5094 72 5097 78
rect 5102 72 5105 108
rect 5150 111 5153 158
rect 5210 148 5214 151
rect 5166 122 5169 138
rect 5174 132 5177 138
rect 5146 108 5153 111
rect 5126 78 5129 108
rect 5158 82 5161 88
rect 5206 72 5209 78
rect 5118 52 5121 58
rect 5026 48 5030 51
rect 5082 48 5086 51
rect 5214 -18 5217 58
rect 5230 -18 5233 348
rect 5270 332 5273 338
rect 5278 332 5281 478
rect 5286 372 5289 418
rect 5310 392 5313 2128
rect 5358 592 5361 2898
rect 5262 272 5265 279
rect 5238 270 5246 271
rect 5242 268 5246 270
rect 5266 268 5273 271
rect 5246 262 5249 268
rect 5270 262 5273 268
rect 5286 262 5289 348
rect 5294 332 5297 338
rect 5298 328 5305 331
rect 5294 292 5297 318
rect 5282 238 5286 241
rect 5270 162 5273 188
rect 5294 172 5297 258
rect 5302 252 5305 328
rect 5238 142 5241 147
rect 5238 82 5241 128
rect 5270 92 5273 148
rect 5286 122 5289 138
rect 5294 72 5297 78
rect 5290 58 5294 61
rect 5270 52 5273 58
rect 5246 -18 5249 8
rect 2326 -19 2330 -18
rect 2318 -22 2330 -19
rect 2358 -22 2362 -18
rect 2446 -22 2450 -18
rect 2510 -22 2514 -18
rect 2558 -22 2562 -18
rect 2926 -22 2930 -18
rect 2942 -22 2946 -18
rect 2982 -22 2986 -18
rect 3006 -22 3010 -18
rect 3086 -22 3090 -18
rect 3182 -22 3186 -18
rect 3342 -22 3346 -18
rect 3502 -22 3506 -18
rect 3558 -22 3562 -18
rect 3718 -22 3722 -18
rect 3878 -22 3882 -18
rect 3990 -22 3994 -18
rect 4022 -22 4026 -18
rect 4046 -22 4050 -18
rect 4094 -22 4098 -18
rect 4118 -22 4122 -18
rect 4190 -22 4194 -18
rect 4214 -22 4218 -18
rect 4230 -22 4234 -18
rect 4422 -22 4426 -18
rect 4486 -22 4490 -18
rect 4534 -22 4538 -18
rect 4686 -22 4690 -18
rect 4974 -22 4978 -18
rect 5214 -22 5218 -18
rect 5230 -22 5234 -18
rect 5246 -22 5250 -18
<< m3contact >>
rect 858 3703 862 3707
rect 865 3703 869 3707
rect 1874 3703 1878 3707
rect 1881 3703 1885 3707
rect 518 3698 522 3702
rect 558 3698 562 3702
rect 694 3698 698 3702
rect 1950 3698 1954 3702
rect 1982 3698 1986 3702
rect 2206 3698 2210 3702
rect 294 3688 298 3692
rect 486 3688 490 3692
rect 422 3678 426 3682
rect 446 3678 450 3682
rect 454 3678 458 3682
rect 478 3678 482 3682
rect 254 3648 258 3652
rect 174 3638 178 3642
rect 262 3638 266 3642
rect 222 3608 226 3612
rect 14 3568 18 3572
rect 174 3568 178 3572
rect 246 3568 250 3572
rect 86 3558 90 3562
rect 174 3558 178 3562
rect 214 3558 218 3562
rect 262 3558 266 3562
rect 118 3548 122 3552
rect 134 3548 138 3552
rect 198 3548 202 3552
rect 214 3548 218 3552
rect 54 3538 58 3542
rect 126 3538 130 3542
rect 78 3528 82 3532
rect 86 3528 90 3532
rect 118 3528 122 3532
rect 230 3528 234 3532
rect 262 3528 266 3532
rect 30 3458 34 3462
rect 62 3458 66 3462
rect 150 3518 154 3522
rect 94 3478 98 3482
rect 110 3478 114 3482
rect 126 3478 130 3482
rect 102 3458 106 3462
rect 230 3518 234 3522
rect 246 3518 250 3522
rect 198 3498 202 3502
rect 118 3458 122 3462
rect 150 3458 154 3462
rect 94 3448 98 3452
rect 134 3448 138 3452
rect 54 3388 58 3392
rect 54 3368 58 3372
rect 246 3498 250 3502
rect 310 3658 314 3662
rect 286 3638 290 3642
rect 318 3628 322 3632
rect 286 3618 290 3622
rect 350 3628 354 3632
rect 542 3678 546 3682
rect 1078 3688 1082 3692
rect 1102 3688 1106 3692
rect 566 3678 570 3682
rect 622 3678 626 3682
rect 734 3678 738 3682
rect 830 3678 834 3682
rect 950 3678 954 3682
rect 982 3678 986 3682
rect 1046 3678 1050 3682
rect 606 3668 610 3672
rect 414 3658 418 3662
rect 462 3658 466 3662
rect 614 3658 618 3662
rect 406 3628 410 3632
rect 342 3618 346 3622
rect 374 3618 378 3622
rect 334 3608 338 3612
rect 346 3603 350 3607
rect 353 3603 357 3607
rect 294 3558 298 3562
rect 278 3528 282 3532
rect 270 3478 274 3482
rect 182 3468 186 3472
rect 198 3458 202 3462
rect 222 3438 226 3442
rect 126 3388 130 3392
rect 142 3368 146 3372
rect 158 3368 162 3372
rect 78 3358 82 3362
rect 190 3368 194 3372
rect 14 3348 18 3352
rect 62 3348 66 3352
rect 150 3348 154 3352
rect 22 3258 26 3262
rect 54 3338 58 3342
rect 94 3338 98 3342
rect 158 3338 162 3342
rect 126 3328 130 3332
rect 54 3278 58 3282
rect 70 3278 74 3282
rect 86 3278 90 3282
rect 54 3268 58 3272
rect 78 3268 82 3272
rect 38 3248 42 3252
rect 62 3248 66 3252
rect 126 3288 130 3292
rect 102 3278 106 3282
rect 110 3278 114 3282
rect 166 3298 170 3302
rect 142 3278 146 3282
rect 118 3268 122 3272
rect 134 3268 138 3272
rect 150 3268 154 3272
rect 206 3308 210 3312
rect 206 3278 210 3282
rect 190 3258 194 3262
rect 238 3458 242 3462
rect 262 3458 266 3462
rect 334 3588 338 3592
rect 430 3558 434 3562
rect 286 3518 290 3522
rect 302 3528 306 3532
rect 318 3528 322 3532
rect 342 3518 346 3522
rect 294 3498 298 3502
rect 302 3468 306 3472
rect 310 3468 314 3472
rect 326 3468 330 3472
rect 286 3458 290 3462
rect 270 3378 274 3382
rect 246 3348 250 3352
rect 222 3298 226 3302
rect 230 3298 234 3302
rect 294 3438 298 3442
rect 286 3388 290 3392
rect 278 3358 282 3362
rect 358 3458 362 3462
rect 318 3448 322 3452
rect 422 3548 426 3552
rect 590 3638 594 3642
rect 726 3668 730 3672
rect 654 3658 658 3662
rect 670 3658 674 3662
rect 630 3648 634 3652
rect 654 3648 658 3652
rect 606 3628 610 3632
rect 622 3628 626 3632
rect 638 3628 642 3632
rect 646 3628 650 3632
rect 574 3618 578 3622
rect 542 3588 546 3592
rect 550 3578 554 3582
rect 454 3548 458 3552
rect 646 3588 650 3592
rect 782 3668 786 3672
rect 910 3668 914 3672
rect 798 3658 802 3662
rect 822 3658 826 3662
rect 846 3658 850 3662
rect 878 3658 882 3662
rect 758 3648 762 3652
rect 774 3648 778 3652
rect 790 3638 794 3642
rect 806 3638 810 3642
rect 742 3618 746 3622
rect 694 3568 698 3572
rect 742 3568 746 3572
rect 774 3608 778 3612
rect 774 3588 778 3592
rect 822 3628 826 3632
rect 830 3608 834 3612
rect 814 3598 818 3602
rect 838 3588 842 3592
rect 558 3558 562 3562
rect 630 3558 634 3562
rect 646 3558 650 3562
rect 686 3558 690 3562
rect 758 3558 762 3562
rect 398 3538 402 3542
rect 470 3538 474 3542
rect 534 3538 538 3542
rect 542 3538 546 3542
rect 558 3538 562 3542
rect 478 3528 482 3532
rect 390 3518 394 3522
rect 494 3518 498 3522
rect 502 3518 506 3522
rect 414 3498 418 3502
rect 390 3468 394 3472
rect 566 3528 570 3532
rect 526 3498 530 3502
rect 590 3498 594 3502
rect 622 3528 626 3532
rect 614 3488 618 3492
rect 718 3548 722 3552
rect 750 3548 754 3552
rect 646 3528 650 3532
rect 718 3528 722 3532
rect 446 3478 450 3482
rect 454 3478 458 3482
rect 542 3478 546 3482
rect 574 3478 578 3482
rect 582 3478 586 3482
rect 606 3478 610 3482
rect 446 3468 450 3472
rect 406 3458 410 3462
rect 454 3458 458 3462
rect 374 3428 378 3432
rect 346 3403 350 3407
rect 353 3403 357 3407
rect 310 3378 314 3382
rect 358 3368 362 3372
rect 382 3368 386 3372
rect 302 3338 306 3342
rect 262 3328 266 3332
rect 294 3328 298 3332
rect 310 3328 314 3332
rect 262 3318 266 3322
rect 254 3288 258 3292
rect 278 3308 282 3312
rect 246 3258 250 3262
rect 262 3258 266 3262
rect 102 3248 106 3252
rect 30 3238 34 3242
rect 94 3238 98 3242
rect 6 3178 10 3182
rect 38 3178 42 3182
rect 110 3178 114 3182
rect 22 3168 26 3172
rect 94 3168 98 3172
rect 182 3238 186 3242
rect 270 3228 274 3232
rect 166 3178 170 3182
rect 134 3168 138 3172
rect 270 3168 274 3172
rect 54 3158 58 3162
rect 78 3158 82 3162
rect 54 3148 58 3152
rect 94 3148 98 3152
rect 30 3138 34 3142
rect 54 3138 58 3142
rect 38 3128 42 3132
rect 70 3128 74 3132
rect 62 3118 66 3122
rect 14 3098 18 3102
rect 54 3098 58 3102
rect 86 3118 90 3122
rect 78 3078 82 3082
rect 54 3048 58 3052
rect 86 3058 90 3062
rect 102 3058 106 3062
rect 118 3148 122 3152
rect 206 3158 210 3162
rect 238 3158 242 3162
rect 142 3148 146 3152
rect 398 3408 402 3412
rect 518 3468 522 3472
rect 494 3458 498 3462
rect 478 3418 482 3422
rect 422 3408 426 3412
rect 446 3388 450 3392
rect 510 3438 514 3442
rect 494 3418 498 3422
rect 398 3378 402 3382
rect 406 3378 410 3382
rect 486 3378 490 3382
rect 414 3368 418 3372
rect 478 3368 482 3372
rect 390 3338 394 3342
rect 414 3338 418 3342
rect 406 3318 410 3322
rect 358 3298 362 3302
rect 382 3298 386 3302
rect 630 3478 634 3482
rect 654 3478 658 3482
rect 678 3478 682 3482
rect 550 3468 554 3472
rect 558 3468 562 3472
rect 590 3468 594 3472
rect 638 3468 642 3472
rect 798 3538 802 3542
rect 782 3498 786 3502
rect 686 3468 690 3472
rect 534 3458 538 3462
rect 566 3458 570 3462
rect 630 3458 634 3462
rect 670 3458 674 3462
rect 590 3448 594 3452
rect 614 3448 618 3452
rect 526 3438 530 3442
rect 526 3428 530 3432
rect 582 3418 586 3422
rect 606 3388 610 3392
rect 534 3378 538 3382
rect 566 3378 570 3382
rect 526 3368 530 3372
rect 550 3368 554 3372
rect 574 3368 578 3372
rect 454 3338 458 3342
rect 550 3338 554 3342
rect 574 3338 578 3342
rect 598 3338 602 3342
rect 430 3328 434 3332
rect 422 3298 426 3302
rect 326 3288 330 3292
rect 494 3328 498 3332
rect 478 3318 482 3322
rect 486 3318 490 3322
rect 390 3278 394 3282
rect 310 3268 314 3272
rect 326 3268 330 3272
rect 334 3258 338 3262
rect 286 3218 290 3222
rect 302 3168 306 3172
rect 318 3168 322 3172
rect 318 3158 322 3162
rect 126 3138 130 3142
rect 150 3118 154 3122
rect 174 3108 178 3112
rect 286 3128 290 3132
rect 302 3128 306 3132
rect 422 3268 426 3272
rect 446 3258 450 3262
rect 470 3258 474 3262
rect 366 3238 370 3242
rect 350 3218 354 3222
rect 346 3203 350 3207
rect 353 3203 357 3207
rect 398 3248 402 3252
rect 422 3188 426 3192
rect 366 3178 370 3182
rect 398 3178 402 3182
rect 374 3158 378 3162
rect 454 3158 458 3162
rect 414 3138 418 3142
rect 350 3128 354 3132
rect 374 3128 378 3132
rect 422 3128 426 3132
rect 438 3128 442 3132
rect 414 3118 418 3122
rect 254 3088 258 3092
rect 286 3088 290 3092
rect 206 3078 210 3082
rect 254 3078 258 3082
rect 294 3078 298 3082
rect 118 3058 122 3062
rect 134 3058 138 3062
rect 78 3048 82 3052
rect 110 3048 114 3052
rect 70 3038 74 3042
rect 94 3038 98 3042
rect 46 3008 50 3012
rect 62 3008 66 3012
rect 62 2968 66 2972
rect 46 2958 50 2962
rect 86 2958 90 2962
rect 70 2948 74 2952
rect 86 2948 90 2952
rect 78 2928 82 2932
rect 22 2908 26 2912
rect 238 3058 242 3062
rect 126 3048 130 3052
rect 158 3048 162 3052
rect 198 3048 202 3052
rect 222 3048 226 3052
rect 230 3048 234 3052
rect 174 3038 178 3042
rect 238 3038 242 3042
rect 246 3038 250 3042
rect 222 3028 226 3032
rect 230 3028 234 3032
rect 206 3018 210 3022
rect 158 2968 162 2972
rect 190 2968 194 2972
rect 406 3078 410 3082
rect 446 3078 450 3082
rect 390 3068 394 3072
rect 422 3068 426 3072
rect 510 3318 514 3322
rect 574 3288 578 3292
rect 502 3278 506 3282
rect 558 3268 562 3272
rect 550 3258 554 3262
rect 582 3258 586 3262
rect 574 3248 578 3252
rect 750 3458 754 3462
rect 758 3418 762 3422
rect 630 3408 634 3412
rect 670 3408 674 3412
rect 662 3398 666 3402
rect 686 3388 690 3392
rect 630 3378 634 3382
rect 654 3348 658 3352
rect 766 3408 770 3412
rect 710 3368 714 3372
rect 718 3368 722 3372
rect 630 3338 634 3342
rect 646 3338 650 3342
rect 894 3628 898 3632
rect 878 3588 882 3592
rect 854 3578 858 3582
rect 822 3558 826 3562
rect 846 3558 850 3562
rect 870 3558 874 3562
rect 878 3508 882 3512
rect 858 3503 862 3507
rect 865 3503 869 3507
rect 822 3488 826 3492
rect 838 3478 842 3482
rect 838 3468 842 3472
rect 798 3458 802 3462
rect 830 3448 834 3452
rect 814 3438 818 3442
rect 854 3458 858 3462
rect 846 3418 850 3422
rect 782 3368 786 3372
rect 798 3368 802 3372
rect 814 3368 818 3372
rect 902 3598 906 3602
rect 918 3558 922 3562
rect 902 3548 906 3552
rect 1214 3688 1218 3692
rect 1222 3688 1226 3692
rect 1742 3688 1746 3692
rect 1774 3688 1778 3692
rect 958 3668 962 3672
rect 990 3668 994 3672
rect 950 3658 954 3662
rect 942 3638 946 3642
rect 998 3658 1002 3662
rect 1046 3658 1050 3662
rect 974 3648 978 3652
rect 1030 3648 1034 3652
rect 1238 3668 1242 3672
rect 1214 3658 1218 3662
rect 1150 3648 1154 3652
rect 1158 3648 1162 3652
rect 1230 3648 1234 3652
rect 1126 3628 1130 3632
rect 966 3618 970 3622
rect 910 3528 914 3532
rect 982 3558 986 3562
rect 1222 3628 1226 3632
rect 1230 3618 1234 3622
rect 1190 3588 1194 3592
rect 1070 3568 1074 3572
rect 1238 3598 1242 3602
rect 950 3548 954 3552
rect 966 3548 970 3552
rect 998 3548 1002 3552
rect 1038 3538 1042 3542
rect 934 3528 938 3532
rect 942 3528 946 3532
rect 926 3508 930 3512
rect 1094 3558 1098 3562
rect 1126 3558 1130 3562
rect 1142 3558 1146 3562
rect 1054 3538 1058 3542
rect 1094 3548 1098 3552
rect 1118 3548 1122 3552
rect 1166 3548 1170 3552
rect 1086 3538 1090 3542
rect 1062 3528 1066 3532
rect 1118 3528 1122 3532
rect 950 3508 954 3512
rect 1014 3508 1018 3512
rect 1006 3498 1010 3502
rect 918 3478 922 3482
rect 926 3478 930 3482
rect 902 3468 906 3472
rect 942 3458 946 3462
rect 910 3448 914 3452
rect 1270 3638 1274 3642
rect 1294 3678 1298 3682
rect 1302 3658 1306 3662
rect 1286 3648 1290 3652
rect 1294 3638 1298 3642
rect 1598 3678 1602 3682
rect 1622 3678 1626 3682
rect 1670 3678 1674 3682
rect 1694 3678 1698 3682
rect 1822 3678 1826 3682
rect 1478 3668 1482 3672
rect 1502 3668 1506 3672
rect 1630 3668 1634 3672
rect 1646 3668 1650 3672
rect 1742 3668 1746 3672
rect 1334 3658 1338 3662
rect 1422 3658 1426 3662
rect 1430 3658 1434 3662
rect 1518 3658 1522 3662
rect 1566 3658 1570 3662
rect 1582 3658 1586 3662
rect 1398 3648 1402 3652
rect 1430 3648 1434 3652
rect 1326 3638 1330 3642
rect 1318 3618 1322 3622
rect 1270 3608 1274 3612
rect 1278 3608 1282 3612
rect 1278 3558 1282 3562
rect 1318 3578 1322 3582
rect 1438 3638 1442 3642
rect 1358 3608 1362 3612
rect 1370 3603 1374 3607
rect 1377 3603 1381 3607
rect 1654 3658 1658 3662
rect 1518 3648 1522 3652
rect 1550 3648 1554 3652
rect 1606 3648 1610 3652
rect 1622 3648 1626 3652
rect 1526 3638 1530 3642
rect 1446 3588 1450 3592
rect 1302 3568 1306 3572
rect 1326 3568 1330 3572
rect 1342 3568 1346 3572
rect 1374 3568 1378 3572
rect 1414 3568 1418 3572
rect 1294 3548 1298 3552
rect 1182 3538 1186 3542
rect 1326 3558 1330 3562
rect 1342 3558 1346 3562
rect 1406 3558 1410 3562
rect 1318 3548 1322 3552
rect 1166 3528 1170 3532
rect 1190 3528 1194 3532
rect 1158 3498 1162 3502
rect 1150 3488 1154 3492
rect 1126 3478 1130 3482
rect 1030 3468 1034 3472
rect 1054 3468 1058 3472
rect 1014 3458 1018 3462
rect 1174 3488 1178 3492
rect 1062 3458 1066 3462
rect 1094 3458 1098 3462
rect 1118 3458 1122 3462
rect 1134 3458 1138 3462
rect 1038 3448 1042 3452
rect 1318 3518 1322 3522
rect 1294 3508 1298 3512
rect 1222 3488 1226 3492
rect 1302 3498 1306 3502
rect 1278 3488 1282 3492
rect 1198 3458 1202 3462
rect 1062 3438 1066 3442
rect 958 3428 962 3432
rect 950 3418 954 3422
rect 1182 3388 1186 3392
rect 1142 3378 1146 3382
rect 1006 3368 1010 3372
rect 1062 3368 1066 3372
rect 1094 3368 1098 3372
rect 1110 3368 1114 3372
rect 950 3358 954 3362
rect 1038 3358 1042 3362
rect 1078 3358 1082 3362
rect 694 3338 698 3342
rect 702 3338 706 3342
rect 734 3340 738 3344
rect 758 3338 762 3342
rect 774 3338 778 3342
rect 878 3338 882 3342
rect 718 3328 722 3332
rect 798 3328 802 3332
rect 814 3328 818 3332
rect 646 3318 650 3322
rect 614 3308 618 3312
rect 718 3288 722 3292
rect 858 3303 862 3307
rect 865 3303 869 3307
rect 782 3298 786 3302
rect 750 3288 754 3292
rect 614 3278 618 3282
rect 670 3278 674 3282
rect 606 3258 610 3262
rect 486 3238 490 3242
rect 494 3238 498 3242
rect 598 3238 602 3242
rect 678 3248 682 3252
rect 686 3238 690 3242
rect 710 3228 714 3232
rect 662 3218 666 3222
rect 470 3208 474 3212
rect 534 3208 538 3212
rect 470 3178 474 3182
rect 478 3168 482 3172
rect 526 3168 530 3172
rect 470 3158 474 3162
rect 566 3198 570 3202
rect 542 3158 546 3162
rect 550 3158 554 3162
rect 710 3158 714 3162
rect 478 3138 482 3142
rect 494 3138 498 3142
rect 526 3138 530 3142
rect 470 3128 474 3132
rect 510 3128 514 3132
rect 462 3108 466 3112
rect 478 3098 482 3102
rect 494 3068 498 3072
rect 350 3058 354 3062
rect 398 3058 402 3062
rect 430 3058 434 3062
rect 446 3058 450 3062
rect 278 3048 282 3052
rect 270 3038 274 3042
rect 254 3028 258 3032
rect 270 2978 274 2982
rect 254 2968 258 2972
rect 134 2958 138 2962
rect 222 2958 226 2962
rect 270 2958 274 2962
rect 150 2948 154 2952
rect 118 2938 122 2942
rect 142 2938 146 2942
rect 158 2938 162 2942
rect 534 3118 538 3122
rect 582 3148 586 3152
rect 630 3148 634 3152
rect 574 3128 578 3132
rect 638 3128 642 3132
rect 686 3128 690 3132
rect 574 3108 578 3112
rect 670 3108 674 3112
rect 830 3288 834 3292
rect 798 3278 802 3282
rect 806 3278 810 3282
rect 830 3278 834 3282
rect 870 3278 874 3282
rect 790 3268 794 3272
rect 726 3258 730 3262
rect 734 3218 738 3222
rect 798 3248 802 3252
rect 814 3248 818 3252
rect 838 3258 842 3262
rect 878 3258 882 3262
rect 854 3238 858 3242
rect 886 3238 890 3242
rect 1006 3338 1010 3342
rect 918 3328 922 3332
rect 966 3328 970 3332
rect 990 3328 994 3332
rect 974 3308 978 3312
rect 902 3298 906 3302
rect 942 3298 946 3302
rect 966 3298 970 3302
rect 982 3298 986 3302
rect 910 3278 914 3282
rect 958 3278 962 3282
rect 1326 3468 1330 3472
rect 1382 3548 1386 3552
rect 1510 3588 1514 3592
rect 1502 3558 1506 3562
rect 1526 3568 1530 3572
rect 1550 3568 1554 3572
rect 1574 3568 1578 3572
rect 1622 3568 1626 3572
rect 1470 3548 1474 3552
rect 1486 3548 1490 3552
rect 1550 3548 1554 3552
rect 1350 3538 1354 3542
rect 1398 3538 1402 3542
rect 1430 3538 1434 3542
rect 1414 3508 1418 3512
rect 1398 3478 1402 3482
rect 1406 3468 1410 3472
rect 1342 3458 1346 3462
rect 1302 3418 1306 3422
rect 1302 3398 1306 3402
rect 1166 3368 1170 3372
rect 1190 3368 1194 3372
rect 1030 3338 1034 3342
rect 1046 3338 1050 3342
rect 1110 3338 1114 3342
rect 1110 3328 1114 3332
rect 1014 3318 1018 3322
rect 1046 3318 1050 3322
rect 1094 3318 1098 3322
rect 1102 3318 1106 3322
rect 1214 3358 1218 3362
rect 1254 3358 1258 3362
rect 1246 3348 1250 3352
rect 1270 3348 1274 3352
rect 1198 3338 1202 3342
rect 1214 3338 1218 3342
rect 1166 3328 1170 3332
rect 1574 3548 1578 3552
rect 1598 3548 1602 3552
rect 1614 3548 1618 3552
rect 1582 3538 1586 3542
rect 1590 3538 1594 3542
rect 1454 3528 1458 3532
rect 1534 3528 1538 3532
rect 1566 3528 1570 3532
rect 1606 3528 1610 3532
rect 1478 3518 1482 3522
rect 1510 3508 1514 3512
rect 1446 3478 1450 3482
rect 1486 3478 1490 3482
rect 1494 3468 1498 3472
rect 1326 3448 1330 3452
rect 1350 3448 1354 3452
rect 1430 3448 1434 3452
rect 1318 3388 1322 3392
rect 1366 3438 1370 3442
rect 1390 3438 1394 3442
rect 1446 3438 1450 3442
rect 1382 3428 1386 3432
rect 1646 3648 1650 3652
rect 1654 3598 1658 3602
rect 1686 3598 1690 3602
rect 1646 3588 1650 3592
rect 2718 3698 2722 3702
rect 2906 3703 2910 3707
rect 2913 3703 2917 3707
rect 3286 3698 3290 3702
rect 2230 3688 2234 3692
rect 2254 3688 2258 3692
rect 2278 3688 2282 3692
rect 2310 3688 2314 3692
rect 2550 3688 2554 3692
rect 2638 3688 2642 3692
rect 2686 3688 2690 3692
rect 1966 3678 1970 3682
rect 1886 3668 1890 3672
rect 1910 3668 1914 3672
rect 1742 3658 1746 3662
rect 1798 3658 1802 3662
rect 1846 3658 1850 3662
rect 1862 3658 1866 3662
rect 1982 3668 1986 3672
rect 1934 3658 1938 3662
rect 1958 3658 1962 3662
rect 1726 3648 1730 3652
rect 1822 3648 1826 3652
rect 1838 3648 1842 3652
rect 1854 3648 1858 3652
rect 1902 3648 1906 3652
rect 2254 3678 2258 3682
rect 2286 3678 2290 3682
rect 2294 3678 2298 3682
rect 2454 3678 2458 3682
rect 2470 3678 2474 3682
rect 3062 3678 3066 3682
rect 3110 3678 3114 3682
rect 3214 3678 3218 3682
rect 3318 3678 3322 3682
rect 3726 3678 3730 3682
rect 1998 3658 2002 3662
rect 1726 3638 1730 3642
rect 1806 3638 1810 3642
rect 1830 3638 1834 3642
rect 1854 3638 1858 3642
rect 1694 3578 1698 3582
rect 1686 3568 1690 3572
rect 1742 3588 1746 3592
rect 1750 3568 1754 3572
rect 1806 3568 1810 3572
rect 1662 3558 1666 3562
rect 1726 3558 1730 3562
rect 1718 3548 1722 3552
rect 1766 3558 1770 3562
rect 1790 3548 1794 3552
rect 1710 3538 1714 3542
rect 1758 3538 1762 3542
rect 1742 3528 1746 3532
rect 1758 3518 1762 3522
rect 1662 3508 1666 3512
rect 1518 3478 1522 3482
rect 1622 3478 1626 3482
rect 1582 3468 1586 3472
rect 1598 3468 1602 3472
rect 1590 3458 1594 3462
rect 1462 3428 1466 3432
rect 1486 3428 1490 3432
rect 1430 3418 1434 3422
rect 1454 3418 1458 3422
rect 1390 3408 1394 3412
rect 1370 3403 1374 3407
rect 1377 3403 1381 3407
rect 1334 3378 1338 3382
rect 1422 3358 1426 3362
rect 1462 3408 1466 3412
rect 1550 3438 1554 3442
rect 1558 3428 1562 3432
rect 1494 3398 1498 3402
rect 1446 3388 1450 3392
rect 1486 3388 1490 3392
rect 1518 3388 1522 3392
rect 1454 3358 1458 3362
rect 1534 3358 1538 3362
rect 1566 3358 1570 3362
rect 1574 3358 1578 3362
rect 1478 3348 1482 3352
rect 1494 3348 1498 3352
rect 1358 3338 1362 3342
rect 1366 3338 1370 3342
rect 1430 3338 1434 3342
rect 1550 3348 1554 3352
rect 1662 3488 1666 3492
rect 1686 3488 1690 3492
rect 1678 3478 1682 3482
rect 1686 3478 1690 3482
rect 1710 3478 1714 3482
rect 1670 3468 1674 3472
rect 1694 3468 1698 3472
rect 1734 3468 1738 3472
rect 1654 3458 1658 3462
rect 1678 3458 1682 3462
rect 1710 3458 1714 3462
rect 1726 3458 1730 3462
rect 1750 3458 1754 3462
rect 1606 3448 1610 3452
rect 1766 3508 1770 3512
rect 1790 3498 1794 3502
rect 1782 3478 1786 3482
rect 1902 3568 1906 3572
rect 1894 3558 1898 3562
rect 1846 3548 1850 3552
rect 1854 3548 1858 3552
rect 1934 3568 1938 3572
rect 1958 3558 1962 3562
rect 1910 3548 1914 3552
rect 1926 3548 1930 3552
rect 1950 3548 1954 3552
rect 1814 3538 1818 3542
rect 1838 3538 1842 3542
rect 1862 3538 1866 3542
rect 1814 3528 1818 3532
rect 1822 3528 1826 3532
rect 1830 3498 1834 3502
rect 1918 3528 1922 3532
rect 1874 3503 1878 3507
rect 1881 3503 1885 3507
rect 1854 3488 1858 3492
rect 1942 3528 1946 3532
rect 1966 3518 1970 3522
rect 2094 3668 2098 3672
rect 2190 3668 2194 3672
rect 2214 3668 2218 3672
rect 2246 3668 2250 3672
rect 2102 3658 2106 3662
rect 2118 3658 2122 3662
rect 2142 3658 2146 3662
rect 2062 3648 2066 3652
rect 2174 3648 2178 3652
rect 2110 3638 2114 3642
rect 2134 3638 2138 3642
rect 2054 3628 2058 3632
rect 2006 3618 2010 3622
rect 2134 3598 2138 3602
rect 2126 3578 2130 3582
rect 2014 3558 2018 3562
rect 2030 3548 2034 3552
rect 2070 3548 2074 3552
rect 2046 3538 2050 3542
rect 2158 3588 2162 3592
rect 2174 3568 2178 3572
rect 2006 3528 2010 3532
rect 1990 3498 1994 3502
rect 2062 3498 2066 3502
rect 1966 3488 1970 3492
rect 2022 3488 2026 3492
rect 1862 3478 1866 3482
rect 1902 3478 1906 3482
rect 1870 3468 1874 3472
rect 1854 3458 1858 3462
rect 1782 3448 1786 3452
rect 1814 3448 1818 3452
rect 1718 3438 1722 3442
rect 1598 3398 1602 3402
rect 1662 3378 1666 3382
rect 1782 3378 1786 3382
rect 1734 3368 1738 3372
rect 1622 3348 1626 3352
rect 1718 3348 1722 3352
rect 1774 3358 1778 3362
rect 1798 3348 1802 3352
rect 1958 3468 1962 3472
rect 1894 3458 1898 3462
rect 1942 3448 1946 3452
rect 1958 3378 1962 3382
rect 2086 3458 2090 3462
rect 2030 3398 2034 3402
rect 2190 3628 2194 3632
rect 2182 3558 2186 3562
rect 2206 3558 2210 3562
rect 2150 3548 2154 3552
rect 2190 3548 2194 3552
rect 2158 3528 2162 3532
rect 2142 3518 2146 3522
rect 2166 3518 2170 3522
rect 2118 3508 2122 3512
rect 2158 3508 2162 3512
rect 2238 3648 2242 3652
rect 2270 3668 2274 3672
rect 2358 3668 2362 3672
rect 2438 3668 2442 3672
rect 2270 3658 2274 3662
rect 2294 3658 2298 3662
rect 2302 3658 2306 3662
rect 2318 3658 2322 3662
rect 2398 3658 2402 3662
rect 2342 3648 2346 3652
rect 2358 3648 2362 3652
rect 2390 3648 2394 3652
rect 2422 3648 2426 3652
rect 2318 3638 2322 3642
rect 2326 3638 2330 3642
rect 2374 3638 2378 3642
rect 2246 3618 2250 3622
rect 2342 3618 2346 3622
rect 2398 3618 2402 3622
rect 2270 3598 2274 3602
rect 2238 3588 2242 3592
rect 2394 3603 2398 3607
rect 2401 3603 2405 3607
rect 2302 3588 2306 3592
rect 2446 3648 2450 3652
rect 2510 3658 2514 3662
rect 2542 3658 2546 3662
rect 2494 3648 2498 3652
rect 2534 3648 2538 3652
rect 2478 3638 2482 3642
rect 2486 3638 2490 3642
rect 2430 3628 2434 3632
rect 2462 3628 2466 3632
rect 2486 3628 2490 3632
rect 2654 3668 2658 3672
rect 2678 3668 2682 3672
rect 2918 3668 2922 3672
rect 2646 3658 2650 3662
rect 2558 3648 2562 3652
rect 2510 3618 2514 3622
rect 2550 3618 2554 3622
rect 2518 3608 2522 3612
rect 2662 3628 2666 3632
rect 2678 3608 2682 3612
rect 2662 3598 2666 3602
rect 2558 3588 2562 3592
rect 2278 3578 2282 3582
rect 2286 3578 2290 3582
rect 2422 3578 2426 3582
rect 2686 3578 2690 3582
rect 2366 3568 2370 3572
rect 2534 3568 2538 3572
rect 2550 3568 2554 3572
rect 2590 3568 2594 3572
rect 2622 3568 2626 3572
rect 2654 3568 2658 3572
rect 2662 3568 2666 3572
rect 2246 3558 2250 3562
rect 2278 3558 2282 3562
rect 2318 3558 2322 3562
rect 2414 3558 2418 3562
rect 2446 3558 2450 3562
rect 2230 3548 2234 3552
rect 2262 3548 2266 3552
rect 2190 3528 2194 3532
rect 2270 3528 2274 3532
rect 2294 3528 2298 3532
rect 2334 3548 2338 3552
rect 2358 3548 2362 3552
rect 2398 3548 2402 3552
rect 2238 3518 2242 3522
rect 2310 3518 2314 3522
rect 2438 3548 2442 3552
rect 2510 3558 2514 3562
rect 2486 3548 2490 3552
rect 2494 3548 2498 3552
rect 2350 3528 2354 3532
rect 2398 3528 2402 3532
rect 2422 3528 2426 3532
rect 2454 3528 2458 3532
rect 2214 3508 2218 3512
rect 2198 3488 2202 3492
rect 2214 3488 2218 3492
rect 2254 3488 2258 3492
rect 2142 3478 2146 3482
rect 2110 3468 2114 3472
rect 2134 3468 2138 3472
rect 2102 3458 2106 3462
rect 2110 3448 2114 3452
rect 2126 3448 2130 3452
rect 2134 3448 2138 3452
rect 2094 3398 2098 3402
rect 1838 3368 1842 3372
rect 2006 3368 2010 3372
rect 2142 3368 2146 3372
rect 2150 3368 2154 3372
rect 1822 3358 1826 3362
rect 1862 3358 1866 3362
rect 1902 3358 1906 3362
rect 2070 3358 2074 3362
rect 1894 3348 1898 3352
rect 2054 3348 2058 3352
rect 2070 3348 2074 3352
rect 1542 3338 1546 3342
rect 1558 3338 1562 3342
rect 1630 3338 1634 3342
rect 1734 3338 1738 3342
rect 1742 3338 1746 3342
rect 1774 3338 1778 3342
rect 1814 3338 1818 3342
rect 1238 3328 1242 3332
rect 1262 3328 1266 3332
rect 1270 3328 1274 3332
rect 1470 3328 1474 3332
rect 1510 3328 1514 3332
rect 1606 3328 1610 3332
rect 1190 3318 1194 3322
rect 1230 3318 1234 3322
rect 1046 3308 1050 3312
rect 1134 3308 1138 3312
rect 1158 3308 1162 3312
rect 1134 3298 1138 3302
rect 1006 3288 1010 3292
rect 1030 3288 1034 3292
rect 1078 3288 1082 3292
rect 998 3278 1002 3282
rect 1014 3278 1018 3282
rect 1118 3278 1122 3282
rect 902 3258 906 3262
rect 910 3258 914 3262
rect 1022 3258 1026 3262
rect 1046 3258 1050 3262
rect 1070 3258 1074 3262
rect 1102 3258 1106 3262
rect 982 3248 986 3252
rect 926 3238 930 3242
rect 966 3238 970 3242
rect 894 3198 898 3202
rect 798 3188 802 3192
rect 830 3188 834 3192
rect 854 3188 858 3192
rect 782 3148 786 3152
rect 942 3168 946 3172
rect 950 3168 954 3172
rect 774 3138 778 3142
rect 878 3138 882 3142
rect 614 3088 618 3092
rect 614 3078 618 3082
rect 678 3068 682 3072
rect 686 3068 690 3072
rect 750 3068 754 3072
rect 422 3048 426 3052
rect 438 3048 442 3052
rect 478 3048 482 3052
rect 502 3048 506 3052
rect 510 3048 514 3052
rect 406 3038 410 3042
rect 398 3028 402 3032
rect 346 3003 350 3007
rect 353 3003 357 3007
rect 382 2968 386 2972
rect 294 2958 298 2962
rect 198 2948 202 2952
rect 230 2948 234 2952
rect 246 2948 250 2952
rect 334 2948 338 2952
rect 382 2948 386 2952
rect 198 2928 202 2932
rect 150 2918 154 2922
rect 206 2918 210 2922
rect 102 2888 106 2892
rect 166 2888 170 2892
rect 190 2888 194 2892
rect 86 2878 90 2882
rect 150 2878 154 2882
rect 158 2878 162 2882
rect 54 2858 58 2862
rect 102 2858 106 2862
rect 134 2848 138 2852
rect 102 2828 106 2832
rect 54 2768 58 2772
rect 86 2768 90 2772
rect 94 2768 98 2772
rect 30 2748 34 2752
rect 62 2748 66 2752
rect 46 2738 50 2742
rect 70 2738 74 2742
rect 62 2728 66 2732
rect 6 2608 10 2612
rect 30 2568 34 2572
rect 142 2758 146 2762
rect 110 2748 114 2752
rect 86 2738 90 2742
rect 102 2738 106 2742
rect 78 2728 82 2732
rect 166 2858 170 2862
rect 174 2848 178 2852
rect 174 2758 178 2762
rect 190 2818 194 2822
rect 174 2738 178 2742
rect 150 2728 154 2732
rect 118 2688 122 2692
rect 70 2678 74 2682
rect 110 2678 114 2682
rect 166 2678 170 2682
rect 118 2668 122 2672
rect 134 2668 138 2672
rect 46 2658 50 2662
rect 78 2658 82 2662
rect 94 2658 98 2662
rect 54 2648 58 2652
rect 158 2658 162 2662
rect 214 2738 218 2742
rect 182 2728 186 2732
rect 222 2708 226 2712
rect 294 2938 298 2942
rect 278 2928 282 2932
rect 278 2888 282 2892
rect 318 2928 322 2932
rect 406 2958 410 2962
rect 446 2958 450 2962
rect 382 2928 386 2932
rect 390 2928 394 2932
rect 342 2918 346 2922
rect 310 2898 314 2902
rect 398 2908 402 2912
rect 550 3058 554 3062
rect 574 3048 578 3052
rect 558 3028 562 3032
rect 590 2988 594 2992
rect 558 2958 562 2962
rect 582 2958 586 2962
rect 478 2948 482 2952
rect 526 2948 530 2952
rect 422 2938 426 2942
rect 446 2928 450 2932
rect 422 2908 426 2912
rect 438 2908 442 2912
rect 294 2878 298 2882
rect 422 2878 426 2882
rect 254 2848 258 2852
rect 278 2858 282 2862
rect 342 2858 346 2862
rect 262 2778 266 2782
rect 238 2768 242 2772
rect 262 2748 266 2752
rect 246 2738 250 2742
rect 254 2708 258 2712
rect 198 2658 202 2662
rect 166 2648 170 2652
rect 190 2648 194 2652
rect 126 2638 130 2642
rect 142 2638 146 2642
rect 150 2638 154 2642
rect 166 2628 170 2632
rect 118 2618 122 2622
rect 94 2608 98 2612
rect 118 2568 122 2572
rect 62 2558 66 2562
rect 22 2548 26 2552
rect 46 2548 50 2552
rect 118 2548 122 2552
rect 54 2528 58 2532
rect 118 2528 122 2532
rect 134 2528 138 2532
rect 110 2518 114 2522
rect 262 2648 266 2652
rect 254 2628 258 2632
rect 206 2608 210 2612
rect 438 2858 442 2862
rect 550 2938 554 2942
rect 486 2918 490 2922
rect 542 2928 546 2932
rect 494 2908 498 2912
rect 510 2908 514 2912
rect 454 2868 458 2872
rect 374 2818 378 2822
rect 346 2803 350 2807
rect 353 2803 357 2807
rect 446 2798 450 2802
rect 302 2778 306 2782
rect 350 2768 354 2772
rect 414 2768 418 2772
rect 278 2758 282 2762
rect 342 2748 346 2752
rect 366 2748 370 2752
rect 302 2728 306 2732
rect 430 2748 434 2752
rect 326 2728 330 2732
rect 342 2728 346 2732
rect 390 2728 394 2732
rect 422 2728 426 2732
rect 310 2718 314 2722
rect 358 2718 362 2722
rect 326 2688 330 2692
rect 302 2668 306 2672
rect 294 2658 298 2662
rect 310 2658 314 2662
rect 278 2648 282 2652
rect 302 2648 306 2652
rect 390 2708 394 2712
rect 470 2818 474 2822
rect 566 2948 570 2952
rect 670 3058 674 3062
rect 670 3038 674 3042
rect 742 3058 746 3062
rect 702 3038 706 3042
rect 750 3038 754 3042
rect 790 3128 794 3132
rect 822 3118 826 3122
rect 798 3078 802 3082
rect 782 3068 786 3072
rect 774 3058 778 3062
rect 858 3103 862 3107
rect 865 3103 869 3107
rect 830 3098 834 3102
rect 902 3128 906 3132
rect 990 3238 994 3242
rect 1006 3238 1010 3242
rect 1142 3238 1146 3242
rect 1038 3218 1042 3222
rect 1134 3218 1138 3222
rect 1158 3258 1162 3262
rect 1702 3328 1706 3332
rect 1710 3328 1714 3332
rect 1326 3318 1330 3322
rect 1470 3318 1474 3322
rect 1534 3318 1538 3322
rect 1654 3318 1658 3322
rect 1350 3298 1354 3302
rect 1254 3288 1258 3292
rect 1286 3288 1290 3292
rect 1390 3288 1394 3292
rect 1246 3278 1250 3282
rect 1350 3278 1354 3282
rect 1190 3248 1194 3252
rect 1438 3278 1442 3282
rect 1454 3278 1458 3282
rect 1486 3268 1490 3272
rect 1206 3238 1210 3242
rect 1198 3228 1202 3232
rect 1150 3218 1154 3222
rect 1254 3248 1258 3252
rect 1262 3248 1266 3252
rect 1278 3248 1282 3252
rect 1318 3258 1322 3262
rect 1294 3248 1298 3252
rect 1286 3238 1290 3242
rect 1294 3228 1298 3232
rect 1270 3218 1274 3222
rect 1390 3248 1394 3252
rect 1370 3203 1374 3207
rect 1377 3203 1381 3207
rect 1230 3188 1234 3192
rect 1310 3188 1314 3192
rect 1222 3178 1226 3182
rect 1238 3178 1242 3182
rect 998 3168 1002 3172
rect 1182 3168 1186 3172
rect 1198 3168 1202 3172
rect 1206 3168 1210 3172
rect 1062 3158 1066 3162
rect 1142 3158 1146 3162
rect 1190 3158 1194 3162
rect 1214 3158 1218 3162
rect 1006 3148 1010 3152
rect 926 3138 930 3142
rect 966 3138 970 3142
rect 990 3138 994 3142
rect 918 3118 922 3122
rect 974 3118 978 3122
rect 1006 3128 1010 3132
rect 910 3098 914 3102
rect 942 3098 946 3102
rect 958 3098 962 3102
rect 990 3098 994 3102
rect 1078 3118 1082 3122
rect 1038 3098 1042 3102
rect 926 3088 930 3092
rect 950 3088 954 3092
rect 974 3088 978 3092
rect 1038 3088 1042 3092
rect 918 3078 922 3082
rect 806 3068 810 3072
rect 838 3068 842 3072
rect 806 3058 810 3062
rect 958 3068 962 3072
rect 1166 3138 1170 3142
rect 1278 3168 1282 3172
rect 1286 3168 1290 3172
rect 1246 3158 1250 3162
rect 1246 3148 1250 3152
rect 1270 3148 1274 3152
rect 1206 3138 1210 3142
rect 1158 3128 1162 3132
rect 1182 3128 1186 3132
rect 1134 3118 1138 3122
rect 1030 3078 1034 3082
rect 1094 3078 1098 3082
rect 990 3068 994 3072
rect 1094 3068 1098 3072
rect 1110 3068 1114 3072
rect 958 3058 962 3062
rect 1006 3058 1010 3062
rect 1038 3058 1042 3062
rect 1054 3058 1058 3062
rect 838 3048 842 3052
rect 846 3048 850 3052
rect 910 3048 914 3052
rect 998 3048 1002 3052
rect 1006 3048 1010 3052
rect 886 3038 890 3042
rect 902 3018 906 3022
rect 742 2988 746 2992
rect 766 2988 770 2992
rect 782 2988 786 2992
rect 686 2968 690 2972
rect 694 2948 698 2952
rect 662 2938 666 2942
rect 606 2918 610 2922
rect 686 2918 690 2922
rect 694 2918 698 2922
rect 590 2888 594 2892
rect 630 2888 634 2892
rect 662 2868 666 2872
rect 574 2818 578 2822
rect 486 2768 490 2772
rect 534 2768 538 2772
rect 494 2758 498 2762
rect 462 2718 466 2722
rect 414 2688 418 2692
rect 454 2688 458 2692
rect 374 2678 378 2682
rect 414 2678 418 2682
rect 430 2678 434 2682
rect 486 2738 490 2742
rect 518 2740 522 2744
rect 630 2858 634 2862
rect 654 2858 658 2862
rect 678 2838 682 2842
rect 606 2828 610 2832
rect 638 2788 642 2792
rect 678 2758 682 2762
rect 590 2748 594 2752
rect 550 2738 554 2742
rect 470 2698 474 2702
rect 518 2728 522 2732
rect 526 2728 530 2732
rect 606 2728 610 2732
rect 558 2698 562 2702
rect 654 2738 658 2742
rect 638 2718 642 2722
rect 582 2688 586 2692
rect 478 2678 482 2682
rect 342 2668 346 2672
rect 382 2668 386 2672
rect 446 2668 450 2672
rect 406 2658 410 2662
rect 438 2658 442 2662
rect 470 2658 474 2662
rect 534 2668 538 2672
rect 574 2668 578 2672
rect 582 2668 586 2672
rect 550 2658 554 2662
rect 398 2648 402 2652
rect 422 2648 426 2652
rect 446 2648 450 2652
rect 454 2648 458 2652
rect 502 2648 506 2652
rect 542 2648 546 2652
rect 270 2578 274 2582
rect 278 2568 282 2572
rect 310 2568 314 2572
rect 270 2558 274 2562
rect 158 2548 162 2552
rect 150 2538 154 2542
rect 166 2538 170 2542
rect 346 2603 350 2607
rect 353 2603 357 2607
rect 342 2588 346 2592
rect 414 2558 418 2562
rect 478 2638 482 2642
rect 558 2648 562 2652
rect 486 2588 490 2592
rect 558 2558 562 2562
rect 582 2558 586 2562
rect 302 2548 306 2552
rect 318 2548 322 2552
rect 518 2548 522 2552
rect 550 2548 554 2552
rect 198 2538 202 2542
rect 262 2538 266 2542
rect 310 2538 314 2542
rect 190 2528 194 2532
rect 206 2528 210 2532
rect 30 2478 34 2482
rect 86 2478 90 2482
rect 110 2478 114 2482
rect 78 2468 82 2472
rect 62 2458 66 2462
rect 78 2458 82 2462
rect 38 2438 42 2442
rect 62 2438 66 2442
rect 150 2478 154 2482
rect 142 2458 146 2462
rect 118 2448 122 2452
rect 22 2408 26 2412
rect 14 2368 18 2372
rect 14 2338 18 2342
rect 166 2468 170 2472
rect 190 2458 194 2462
rect 158 2448 162 2452
rect 134 2438 138 2442
rect 166 2438 170 2442
rect 30 2378 34 2382
rect 294 2488 298 2492
rect 374 2488 378 2492
rect 214 2478 218 2482
rect 310 2478 314 2482
rect 358 2478 362 2482
rect 246 2468 250 2472
rect 278 2468 282 2472
rect 318 2468 322 2472
rect 198 2418 202 2422
rect 270 2448 274 2452
rect 310 2458 314 2462
rect 334 2448 338 2452
rect 294 2438 298 2442
rect 310 2438 314 2442
rect 198 2408 202 2412
rect 222 2408 226 2412
rect 302 2418 306 2422
rect 382 2428 386 2432
rect 326 2418 330 2422
rect 342 2418 346 2422
rect 198 2368 202 2372
rect 38 2358 42 2362
rect 118 2358 122 2362
rect 166 2358 170 2362
rect 150 2348 154 2352
rect 86 2338 90 2342
rect 118 2338 122 2342
rect 54 2308 58 2312
rect 62 2288 66 2292
rect 158 2328 162 2332
rect 142 2318 146 2322
rect 110 2288 114 2292
rect 174 2308 178 2312
rect 254 2358 258 2362
rect 278 2358 282 2362
rect 206 2348 210 2352
rect 230 2348 234 2352
rect 222 2338 226 2342
rect 206 2308 210 2312
rect 190 2278 194 2282
rect 382 2408 386 2412
rect 346 2403 350 2407
rect 353 2403 357 2407
rect 454 2518 458 2522
rect 454 2508 458 2512
rect 502 2538 506 2542
rect 502 2528 506 2532
rect 518 2518 522 2522
rect 510 2488 514 2492
rect 486 2458 490 2462
rect 494 2458 498 2462
rect 526 2458 530 2462
rect 414 2438 418 2442
rect 502 2418 506 2422
rect 398 2408 402 2412
rect 350 2388 354 2392
rect 390 2388 394 2392
rect 478 2388 482 2392
rect 486 2388 490 2392
rect 318 2348 322 2352
rect 270 2338 274 2342
rect 302 2338 306 2342
rect 326 2338 330 2342
rect 254 2308 258 2312
rect 214 2298 218 2302
rect 230 2298 234 2302
rect 246 2298 250 2302
rect 214 2278 218 2282
rect 270 2298 274 2302
rect 422 2368 426 2372
rect 486 2368 490 2372
rect 374 2348 378 2352
rect 414 2348 418 2352
rect 430 2348 434 2352
rect 366 2338 370 2342
rect 374 2318 378 2322
rect 422 2338 426 2342
rect 406 2318 410 2322
rect 502 2348 506 2352
rect 518 2348 522 2352
rect 510 2338 514 2342
rect 454 2318 458 2322
rect 262 2288 266 2292
rect 286 2288 290 2292
rect 310 2278 314 2282
rect 382 2278 386 2282
rect 398 2278 402 2282
rect 518 2318 522 2322
rect 566 2548 570 2552
rect 598 2528 602 2532
rect 710 2978 714 2982
rect 766 2978 770 2982
rect 726 2948 730 2952
rect 734 2948 738 2952
rect 758 2948 762 2952
rect 718 2938 722 2942
rect 766 2938 770 2942
rect 870 2948 874 2952
rect 854 2938 858 2942
rect 758 2928 762 2932
rect 782 2928 786 2932
rect 822 2918 826 2922
rect 858 2903 862 2907
rect 865 2903 869 2907
rect 1014 3038 1018 3042
rect 1046 3038 1050 3042
rect 1062 3038 1066 3042
rect 934 2938 938 2942
rect 1014 2998 1018 3002
rect 966 2958 970 2962
rect 1078 3038 1082 3042
rect 1118 3038 1122 3042
rect 1190 3098 1194 3102
rect 1150 3078 1154 3082
rect 1174 3058 1178 3062
rect 1102 3028 1106 3032
rect 1118 3028 1122 3032
rect 1134 3028 1138 3032
rect 1142 2958 1146 2962
rect 1126 2948 1130 2952
rect 1142 2948 1146 2952
rect 1190 3048 1194 3052
rect 1166 2958 1170 2962
rect 1158 2948 1162 2952
rect 998 2938 1002 2942
rect 1070 2938 1074 2942
rect 1078 2938 1082 2942
rect 942 2928 946 2932
rect 982 2908 986 2912
rect 1038 2908 1042 2912
rect 838 2898 842 2902
rect 910 2898 914 2902
rect 934 2898 938 2902
rect 734 2888 738 2892
rect 766 2888 770 2892
rect 1070 2888 1074 2892
rect 1222 3138 1226 3142
rect 1262 3138 1266 3142
rect 1302 3138 1306 3142
rect 1270 3128 1274 3132
rect 1334 3128 1338 3132
rect 1214 3118 1218 3122
rect 1294 3118 1298 3122
rect 1214 3108 1218 3112
rect 1238 3098 1242 3102
rect 1270 3098 1274 3102
rect 1222 3058 1226 3062
rect 1254 3058 1258 3062
rect 1230 3048 1234 3052
rect 1286 3048 1290 3052
rect 1430 3188 1434 3192
rect 1422 3158 1426 3162
rect 1350 3138 1354 3142
rect 1350 3128 1354 3132
rect 1342 3108 1346 3112
rect 1390 3128 1394 3132
rect 1374 3118 1378 3122
rect 1366 3108 1370 3112
rect 1406 3148 1410 3152
rect 1366 3078 1370 3082
rect 1430 3138 1434 3142
rect 1414 3118 1418 3122
rect 1446 3258 1450 3262
rect 1462 3248 1466 3252
rect 1494 3248 1498 3252
rect 1510 3248 1514 3252
rect 1470 3218 1474 3222
rect 1686 3308 1690 3312
rect 1734 3318 1738 3322
rect 1646 3278 1650 3282
rect 1678 3278 1682 3282
rect 1694 3278 1698 3282
rect 1542 3268 1546 3272
rect 1566 3268 1570 3272
rect 1574 3268 1578 3272
rect 1670 3268 1674 3272
rect 1686 3268 1690 3272
rect 1638 3258 1642 3262
rect 1558 3248 1562 3252
rect 1582 3248 1586 3252
rect 1654 3248 1658 3252
rect 1614 3238 1618 3242
rect 1526 3228 1530 3232
rect 1558 3228 1562 3232
rect 1694 3258 1698 3262
rect 1718 3258 1722 3262
rect 1734 3258 1738 3262
rect 1718 3248 1722 3252
rect 1646 3178 1650 3182
rect 1454 3148 1458 3152
rect 1446 3118 1450 3122
rect 1590 3158 1594 3162
rect 1486 3148 1490 3152
rect 1534 3148 1538 3152
rect 1582 3148 1586 3152
rect 1518 3138 1522 3142
rect 1518 3128 1522 3132
rect 1510 3118 1514 3122
rect 1470 3108 1474 3112
rect 1478 3108 1482 3112
rect 1438 3098 1442 3102
rect 1534 3128 1538 3132
rect 1574 3138 1578 3142
rect 1630 3148 1634 3152
rect 1614 3138 1618 3142
rect 1550 3118 1554 3122
rect 1582 3108 1586 3112
rect 1550 3088 1554 3092
rect 1422 3078 1426 3082
rect 1526 3078 1530 3082
rect 1542 3078 1546 3082
rect 1414 3068 1418 3072
rect 1438 3068 1442 3072
rect 1462 3068 1466 3072
rect 1302 3058 1306 3062
rect 1310 3058 1314 3062
rect 1382 3058 1386 3062
rect 1446 3058 1450 3062
rect 1318 3048 1322 3052
rect 1390 3048 1394 3052
rect 1238 3038 1242 3042
rect 1294 3038 1298 3042
rect 1326 3038 1330 3042
rect 1230 3018 1234 3022
rect 1370 3003 1374 3007
rect 1377 3003 1381 3007
rect 1486 3066 1490 3070
rect 1534 3068 1538 3072
rect 1622 3118 1626 3122
rect 1630 3108 1634 3112
rect 1718 3168 1722 3172
rect 1662 3158 1666 3162
rect 1782 3258 1786 3262
rect 1774 3248 1778 3252
rect 1862 3338 1866 3342
rect 1814 3328 1818 3332
rect 1838 3328 1842 3332
rect 1874 3303 1878 3307
rect 1881 3303 1885 3307
rect 1830 3298 1834 3302
rect 1838 3278 1842 3282
rect 1806 3258 1810 3262
rect 1758 3238 1762 3242
rect 1886 3258 1890 3262
rect 1838 3248 1842 3252
rect 1870 3248 1874 3252
rect 1870 3178 1874 3182
rect 1862 3158 1866 3162
rect 1710 3148 1714 3152
rect 1742 3148 1746 3152
rect 1750 3148 1754 3152
rect 1782 3148 1786 3152
rect 1830 3148 1834 3152
rect 1694 3138 1698 3142
rect 1726 3140 1730 3144
rect 1926 3288 1930 3292
rect 1990 3288 1994 3292
rect 2006 3318 2010 3322
rect 1982 3278 1986 3282
rect 1966 3258 1970 3262
rect 2038 3308 2042 3312
rect 2054 3328 2058 3332
rect 2014 3288 2018 3292
rect 2022 3288 2026 3292
rect 2030 3288 2034 3292
rect 1934 3248 1938 3252
rect 1982 3248 1986 3252
rect 1998 3238 2002 3242
rect 1926 3178 1930 3182
rect 1918 3168 1922 3172
rect 1966 3168 1970 3172
rect 1926 3158 1930 3162
rect 1942 3158 1946 3162
rect 1958 3148 1962 3152
rect 2078 3338 2082 3342
rect 2150 3358 2154 3362
rect 2094 3348 2098 3352
rect 2110 3338 2114 3342
rect 2142 3348 2146 3352
rect 2126 3328 2130 3332
rect 2094 3318 2098 3322
rect 2078 3268 2082 3272
rect 2022 3258 2026 3262
rect 2054 3258 2058 3262
rect 2062 3258 2066 3262
rect 2046 3248 2050 3252
rect 2086 3248 2090 3252
rect 2166 3348 2170 3352
rect 2158 3338 2162 3342
rect 2198 3478 2202 3482
rect 2222 3478 2226 3482
rect 2310 3478 2314 3482
rect 2326 3478 2330 3482
rect 2358 3478 2362 3482
rect 2286 3468 2290 3472
rect 2302 3468 2306 3472
rect 2214 3458 2218 3462
rect 2294 3458 2298 3462
rect 2230 3448 2234 3452
rect 2254 3448 2258 3452
rect 2278 3448 2282 3452
rect 2318 3448 2322 3452
rect 2350 3448 2354 3452
rect 2206 3428 2210 3432
rect 2206 3378 2210 3382
rect 2190 3338 2194 3342
rect 2174 3328 2178 3332
rect 2182 3328 2186 3332
rect 2198 3288 2202 3292
rect 2118 3268 2122 3272
rect 2110 3258 2114 3262
rect 2102 3248 2106 3252
rect 2142 3248 2146 3252
rect 2174 3238 2178 3242
rect 2150 3218 2154 3222
rect 1766 3138 1770 3142
rect 1806 3138 1810 3142
rect 1902 3138 1906 3142
rect 1670 3128 1674 3132
rect 1782 3108 1786 3112
rect 1874 3103 1878 3107
rect 1881 3103 1885 3107
rect 1830 3098 1834 3102
rect 1654 3088 1658 3092
rect 1750 3088 1754 3092
rect 1990 3088 1994 3092
rect 1998 3088 2002 3092
rect 1990 3078 1994 3082
rect 1654 3068 1658 3072
rect 1742 3068 1746 3072
rect 2006 3068 2010 3072
rect 1470 3048 1474 3052
rect 1718 3048 1722 3052
rect 1726 3048 1730 3052
rect 1790 3048 1794 3052
rect 1518 3038 1522 3042
rect 1470 3028 1474 3032
rect 1478 2988 1482 2992
rect 1574 2988 1578 2992
rect 1430 2968 1434 2972
rect 1454 2968 1458 2972
rect 1222 2958 1226 2962
rect 1342 2958 1346 2962
rect 1406 2958 1410 2962
rect 1198 2948 1202 2952
rect 1206 2938 1210 2942
rect 1294 2938 1298 2942
rect 1438 2938 1442 2942
rect 1094 2888 1098 2892
rect 1230 2888 1234 2892
rect 742 2878 746 2882
rect 918 2878 922 2882
rect 1014 2878 1018 2882
rect 1078 2878 1082 2882
rect 1182 2878 1186 2882
rect 806 2868 810 2872
rect 1254 2868 1258 2872
rect 1374 2868 1378 2872
rect 774 2848 778 2852
rect 734 2768 738 2772
rect 750 2748 754 2752
rect 766 2748 770 2752
rect 710 2738 714 2742
rect 742 2718 746 2722
rect 766 2708 770 2712
rect 798 2858 802 2862
rect 902 2848 906 2852
rect 998 2848 1002 2852
rect 1214 2858 1218 2862
rect 1230 2858 1234 2862
rect 1302 2858 1306 2862
rect 1166 2848 1170 2852
rect 918 2838 922 2842
rect 1094 2838 1098 2842
rect 1174 2818 1178 2822
rect 798 2758 802 2762
rect 846 2758 850 2762
rect 1118 2758 1122 2762
rect 902 2748 906 2752
rect 950 2748 954 2752
rect 982 2748 986 2752
rect 1086 2748 1090 2752
rect 806 2738 810 2742
rect 806 2728 810 2732
rect 814 2728 818 2732
rect 830 2728 834 2732
rect 790 2718 794 2722
rect 902 2728 906 2732
rect 846 2718 850 2722
rect 870 2718 874 2722
rect 926 2718 930 2722
rect 782 2688 786 2692
rect 858 2703 862 2707
rect 865 2703 869 2707
rect 894 2698 898 2702
rect 894 2688 898 2692
rect 646 2678 650 2682
rect 654 2678 658 2682
rect 734 2678 738 2682
rect 934 2708 938 2712
rect 966 2728 970 2732
rect 974 2718 978 2722
rect 982 2718 986 2722
rect 950 2688 954 2692
rect 662 2668 666 2672
rect 822 2668 826 2672
rect 838 2668 842 2672
rect 918 2668 922 2672
rect 646 2628 650 2632
rect 622 2608 626 2612
rect 638 2558 642 2562
rect 622 2548 626 2552
rect 614 2528 618 2532
rect 670 2658 674 2662
rect 694 2658 698 2662
rect 718 2658 722 2662
rect 806 2648 810 2652
rect 718 2598 722 2602
rect 742 2598 746 2602
rect 798 2598 802 2602
rect 742 2578 746 2582
rect 758 2578 762 2582
rect 790 2578 794 2582
rect 1006 2698 1010 2702
rect 1006 2678 1010 2682
rect 1094 2728 1098 2732
rect 1046 2688 1050 2692
rect 1158 2738 1162 2742
rect 1118 2728 1122 2732
rect 1142 2728 1146 2732
rect 1166 2728 1170 2732
rect 1118 2688 1122 2692
rect 1054 2678 1058 2682
rect 1110 2678 1114 2682
rect 1182 2758 1186 2762
rect 1206 2758 1210 2762
rect 1182 2738 1186 2742
rect 1182 2708 1186 2712
rect 1222 2748 1226 2752
rect 1246 2748 1250 2752
rect 1262 2748 1266 2752
rect 1206 2738 1210 2742
rect 1246 2738 1250 2742
rect 1270 2728 1274 2732
rect 1262 2708 1266 2712
rect 1198 2688 1202 2692
rect 1022 2668 1026 2672
rect 1038 2668 1042 2672
rect 1054 2668 1058 2672
rect 1086 2668 1090 2672
rect 1110 2668 1114 2672
rect 1158 2668 1162 2672
rect 1166 2668 1170 2672
rect 830 2658 834 2662
rect 894 2658 898 2662
rect 942 2658 946 2662
rect 958 2658 962 2662
rect 990 2658 994 2662
rect 886 2628 890 2632
rect 846 2598 850 2602
rect 710 2568 714 2572
rect 798 2568 802 2572
rect 670 2548 674 2552
rect 686 2538 690 2542
rect 678 2528 682 2532
rect 654 2498 658 2502
rect 742 2558 746 2562
rect 782 2558 786 2562
rect 806 2558 810 2562
rect 854 2558 858 2562
rect 774 2548 778 2552
rect 742 2538 746 2542
rect 782 2538 786 2542
rect 702 2508 706 2512
rect 766 2508 770 2512
rect 630 2488 634 2492
rect 734 2478 738 2482
rect 678 2468 682 2472
rect 574 2458 578 2462
rect 702 2458 706 2462
rect 710 2458 714 2462
rect 638 2438 642 2442
rect 686 2438 690 2442
rect 678 2428 682 2432
rect 598 2368 602 2372
rect 622 2368 626 2372
rect 678 2368 682 2372
rect 614 2348 618 2352
rect 630 2348 634 2352
rect 646 2348 650 2352
rect 694 2358 698 2362
rect 718 2448 722 2452
rect 774 2468 778 2472
rect 734 2448 738 2452
rect 750 2448 754 2452
rect 726 2438 730 2442
rect 718 2368 722 2372
rect 814 2548 818 2552
rect 862 2548 866 2552
rect 902 2548 906 2552
rect 790 2528 794 2532
rect 806 2528 810 2532
rect 838 2538 842 2542
rect 910 2538 914 2542
rect 910 2528 914 2532
rect 858 2503 862 2507
rect 865 2503 869 2507
rect 814 2488 818 2492
rect 830 2488 834 2492
rect 814 2478 818 2482
rect 854 2478 858 2482
rect 798 2468 802 2472
rect 774 2448 778 2452
rect 806 2438 810 2442
rect 838 2468 842 2472
rect 894 2468 898 2472
rect 822 2448 826 2452
rect 758 2428 762 2432
rect 790 2428 794 2432
rect 814 2428 818 2432
rect 766 2388 770 2392
rect 798 2378 802 2382
rect 766 2368 770 2372
rect 790 2368 794 2372
rect 742 2358 746 2362
rect 750 2358 754 2362
rect 726 2348 730 2352
rect 638 2338 642 2342
rect 654 2338 658 2342
rect 678 2338 682 2342
rect 534 2328 538 2332
rect 630 2328 634 2332
rect 614 2318 618 2322
rect 590 2308 594 2312
rect 678 2318 682 2322
rect 742 2338 746 2342
rect 782 2348 786 2352
rect 894 2448 898 2452
rect 1046 2658 1050 2662
rect 966 2648 970 2652
rect 950 2628 954 2632
rect 966 2628 970 2632
rect 950 2578 954 2582
rect 1006 2608 1010 2612
rect 1022 2588 1026 2592
rect 982 2558 986 2562
rect 990 2548 994 2552
rect 966 2518 970 2522
rect 934 2478 938 2482
rect 950 2478 954 2482
rect 894 2438 898 2442
rect 918 2438 922 2442
rect 862 2368 866 2372
rect 814 2348 818 2352
rect 734 2328 738 2332
rect 758 2328 762 2332
rect 926 2418 930 2422
rect 942 2448 946 2452
rect 958 2428 962 2432
rect 934 2378 938 2382
rect 910 2358 914 2362
rect 998 2518 1002 2522
rect 1078 2658 1082 2662
rect 1062 2648 1066 2652
rect 1078 2608 1082 2612
rect 1134 2658 1138 2662
rect 1142 2648 1146 2652
rect 1118 2628 1122 2632
rect 1110 2608 1114 2612
rect 1134 2608 1138 2612
rect 1254 2678 1258 2682
rect 1214 2668 1218 2672
rect 1230 2668 1234 2672
rect 1246 2668 1250 2672
rect 1214 2658 1218 2662
rect 1254 2658 1258 2662
rect 1262 2658 1266 2662
rect 1206 2648 1210 2652
rect 1198 2588 1202 2592
rect 1078 2578 1082 2582
rect 1110 2578 1114 2582
rect 1102 2558 1106 2562
rect 1078 2548 1082 2552
rect 1078 2538 1082 2542
rect 1054 2528 1058 2532
rect 1022 2518 1026 2522
rect 1038 2518 1042 2522
rect 1094 2538 1098 2542
rect 1086 2508 1090 2512
rect 1214 2618 1218 2622
rect 1270 2628 1274 2632
rect 1566 2958 1570 2962
rect 2022 3058 2026 3062
rect 2078 3098 2082 3102
rect 2062 3078 2066 3082
rect 2054 3058 2058 3062
rect 2094 3098 2098 3102
rect 2086 3068 2090 3072
rect 2174 3168 2178 3172
rect 2158 3158 2162 3162
rect 2238 3298 2242 3302
rect 2222 3288 2226 3292
rect 2238 3288 2242 3292
rect 2334 3438 2338 3442
rect 2422 3508 2426 3512
rect 2398 3468 2402 3472
rect 2406 3458 2410 3462
rect 2382 3448 2386 3452
rect 2606 3558 2610 3562
rect 2630 3558 2634 3562
rect 2742 3658 2746 3662
rect 2726 3578 2730 3582
rect 2838 3648 2842 3652
rect 3118 3668 3122 3672
rect 2870 3658 2874 3662
rect 2910 3658 2914 3662
rect 2902 3648 2906 3652
rect 2854 3638 2858 3642
rect 2782 3628 2786 3632
rect 2966 3618 2970 3622
rect 3326 3668 3330 3672
rect 3462 3668 3466 3672
rect 3670 3668 3674 3672
rect 3742 3668 3746 3672
rect 3094 3658 3098 3662
rect 3110 3658 3114 3662
rect 3150 3658 3154 3662
rect 3078 3638 3082 3642
rect 3078 3628 3082 3632
rect 3006 3618 3010 3622
rect 2862 3608 2866 3612
rect 2990 3608 2994 3612
rect 2774 3598 2778 3602
rect 2798 3598 2802 3602
rect 2742 3568 2746 3572
rect 2582 3548 2586 3552
rect 2542 3538 2546 3542
rect 2558 3538 2562 3542
rect 2534 3528 2538 3532
rect 2510 3518 2514 3522
rect 2494 3508 2498 3512
rect 2470 3498 2474 3502
rect 2462 3468 2466 3472
rect 2470 3458 2474 3462
rect 2326 3418 2330 3422
rect 2318 3388 2322 3392
rect 2278 3378 2282 3382
rect 2394 3403 2398 3407
rect 2401 3403 2405 3407
rect 2334 3368 2338 3372
rect 2350 3368 2354 3372
rect 2382 3368 2386 3372
rect 2318 3358 2322 3362
rect 2342 3358 2346 3362
rect 2302 3348 2306 3352
rect 2294 3338 2298 3342
rect 2302 3328 2306 3332
rect 2318 3328 2322 3332
rect 2358 3328 2362 3332
rect 2262 3318 2266 3322
rect 2318 3318 2322 3322
rect 2310 3308 2314 3312
rect 2358 3308 2362 3312
rect 2270 3288 2274 3292
rect 2302 3288 2306 3292
rect 2254 3268 2258 3272
rect 2214 3258 2218 3262
rect 2230 3258 2234 3262
rect 2206 3158 2210 3162
rect 2358 3298 2362 3302
rect 2278 3258 2282 3262
rect 2278 3248 2282 3252
rect 2318 3248 2322 3252
rect 2326 3248 2330 3252
rect 2350 3248 2354 3252
rect 2270 3188 2274 3192
rect 2262 3148 2266 3152
rect 2166 3128 2170 3132
rect 2206 3118 2210 3122
rect 2086 3058 2090 3062
rect 1902 3048 1906 3052
rect 1918 3048 1922 3052
rect 2038 3048 2042 3052
rect 2046 3048 2050 3052
rect 2110 3048 2114 3052
rect 1822 3038 1826 3042
rect 1838 3038 1842 3042
rect 1870 3038 1874 3042
rect 1902 3038 1906 3042
rect 1814 2968 1818 2972
rect 1790 2958 1794 2962
rect 1846 2968 1850 2972
rect 1862 2968 1866 2972
rect 1550 2948 1554 2952
rect 1398 2918 1402 2922
rect 1326 2858 1330 2862
rect 1390 2858 1394 2862
rect 1318 2838 1322 2842
rect 1286 2828 1290 2832
rect 1370 2803 1374 2807
rect 1377 2803 1381 2807
rect 1350 2788 1354 2792
rect 1318 2728 1322 2732
rect 1414 2888 1418 2892
rect 1438 2868 1442 2872
rect 1446 2858 1450 2862
rect 1806 2948 1810 2952
rect 1846 2948 1850 2952
rect 2038 3028 2042 3032
rect 1998 3018 2002 3022
rect 2022 2998 2026 3002
rect 1974 2968 1978 2972
rect 1958 2958 1962 2962
rect 1614 2938 1618 2942
rect 1646 2938 1650 2942
rect 1710 2938 1714 2942
rect 1774 2938 1778 2942
rect 1854 2938 1858 2942
rect 1790 2928 1794 2932
rect 1574 2888 1578 2892
rect 1646 2888 1650 2892
rect 1678 2888 1682 2892
rect 1590 2868 1594 2872
rect 1638 2868 1642 2872
rect 1502 2858 1506 2862
rect 1470 2818 1474 2822
rect 1454 2758 1458 2762
rect 1494 2758 1498 2762
rect 1438 2748 1442 2752
rect 1454 2748 1458 2752
rect 1302 2688 1306 2692
rect 1326 2678 1330 2682
rect 1342 2668 1346 2672
rect 1366 2668 1370 2672
rect 1286 2648 1290 2652
rect 1310 2648 1314 2652
rect 1302 2628 1306 2632
rect 1278 2618 1282 2622
rect 1310 2618 1314 2622
rect 1366 2648 1370 2652
rect 1350 2638 1354 2642
rect 1246 2588 1250 2592
rect 1294 2548 1298 2552
rect 1102 2508 1106 2512
rect 1094 2488 1098 2492
rect 1190 2518 1194 2522
rect 1174 2508 1178 2512
rect 1158 2498 1162 2502
rect 1134 2488 1138 2492
rect 1126 2478 1130 2482
rect 1254 2528 1258 2532
rect 1326 2538 1330 2542
rect 1278 2508 1282 2512
rect 1318 2498 1322 2502
rect 1206 2488 1210 2492
rect 1246 2488 1250 2492
rect 1142 2478 1146 2482
rect 1198 2478 1202 2482
rect 1014 2438 1018 2442
rect 1038 2398 1042 2402
rect 1030 2388 1034 2392
rect 982 2368 986 2372
rect 1014 2368 1018 2372
rect 1022 2368 1026 2372
rect 942 2348 946 2352
rect 966 2348 970 2352
rect 894 2338 898 2342
rect 974 2338 978 2342
rect 694 2308 698 2312
rect 806 2308 810 2312
rect 526 2288 530 2292
rect 662 2288 666 2292
rect 654 2278 658 2282
rect 102 2268 106 2272
rect 158 2268 162 2272
rect 342 2268 346 2272
rect 422 2268 426 2272
rect 478 2268 482 2272
rect 542 2268 546 2272
rect 558 2268 562 2272
rect 598 2268 602 2272
rect 54 2258 58 2262
rect 110 2258 114 2262
rect 6 2198 10 2202
rect 174 2258 178 2262
rect 190 2258 194 2262
rect 238 2258 242 2262
rect 318 2258 322 2262
rect 206 2248 210 2252
rect 366 2238 370 2242
rect 326 2228 330 2232
rect 366 2218 370 2222
rect 346 2203 350 2207
rect 353 2203 357 2207
rect 430 2258 434 2262
rect 454 2258 458 2262
rect 406 2248 410 2252
rect 414 2238 418 2242
rect 374 2208 378 2212
rect 158 2178 162 2182
rect 534 2228 538 2232
rect 550 2258 554 2262
rect 590 2258 594 2262
rect 858 2303 862 2307
rect 865 2303 869 2307
rect 790 2298 794 2302
rect 1014 2358 1018 2362
rect 998 2348 1002 2352
rect 958 2328 962 2332
rect 926 2318 930 2322
rect 990 2308 994 2312
rect 926 2278 930 2282
rect 798 2268 802 2272
rect 710 2258 714 2262
rect 646 2248 650 2252
rect 758 2248 762 2252
rect 550 2238 554 2242
rect 678 2238 682 2242
rect 542 2218 546 2222
rect 566 2208 570 2212
rect 486 2188 490 2192
rect 462 2178 466 2182
rect 534 2178 538 2182
rect 638 2178 642 2182
rect 694 2178 698 2182
rect 126 2168 130 2172
rect 158 2168 162 2172
rect 166 2168 170 2172
rect 278 2168 282 2172
rect 414 2168 418 2172
rect 54 2158 58 2162
rect 62 2158 66 2162
rect 110 2148 114 2152
rect 78 2138 82 2142
rect 102 2138 106 2142
rect 174 2158 178 2162
rect 214 2158 218 2162
rect 134 2148 138 2152
rect 158 2148 162 2152
rect 206 2148 210 2152
rect 54 2128 58 2132
rect 70 2128 74 2132
rect 78 2128 82 2132
rect 94 2128 98 2132
rect 110 2128 114 2132
rect 22 2108 26 2112
rect 46 2108 50 2112
rect 30 2098 34 2102
rect 110 2108 114 2112
rect 142 2138 146 2142
rect 134 2098 138 2102
rect 174 2098 178 2102
rect 86 2078 90 2082
rect 142 2078 146 2082
rect 62 2068 66 2072
rect 6 1978 10 1982
rect 14 1898 18 1902
rect 38 2048 42 2052
rect 78 2048 82 2052
rect 110 2038 114 2042
rect 134 2038 138 2042
rect 158 2068 162 2072
rect 150 2058 154 2062
rect 238 2138 242 2142
rect 206 2128 210 2132
rect 174 2078 178 2082
rect 206 2078 210 2082
rect 262 2128 266 2132
rect 230 2088 234 2092
rect 398 2158 402 2162
rect 390 2148 394 2152
rect 286 2138 290 2142
rect 350 2138 354 2142
rect 382 2138 386 2142
rect 342 2128 346 2132
rect 366 2128 370 2132
rect 270 2108 274 2112
rect 318 2108 322 2112
rect 254 2088 258 2092
rect 350 2118 354 2122
rect 454 2158 458 2162
rect 478 2158 482 2162
rect 422 2148 426 2152
rect 406 2108 410 2112
rect 446 2148 450 2152
rect 438 2128 442 2132
rect 438 2098 442 2102
rect 398 2088 402 2092
rect 422 2088 426 2092
rect 454 2088 458 2092
rect 246 2078 250 2082
rect 430 2078 434 2082
rect 438 2078 442 2082
rect 622 2158 626 2162
rect 518 2148 522 2152
rect 558 2148 562 2152
rect 662 2168 666 2172
rect 678 2168 682 2172
rect 686 2168 690 2172
rect 662 2158 666 2162
rect 606 2148 610 2152
rect 622 2148 626 2152
rect 646 2148 650 2152
rect 542 2138 546 2142
rect 582 2138 586 2142
rect 598 2138 602 2142
rect 566 2128 570 2132
rect 494 2108 498 2112
rect 486 2088 490 2092
rect 742 2168 746 2172
rect 798 2228 802 2232
rect 854 2228 858 2232
rect 766 2188 770 2192
rect 774 2188 778 2192
rect 702 2148 706 2152
rect 758 2148 762 2152
rect 662 2128 666 2132
rect 606 2118 610 2122
rect 622 2118 626 2122
rect 582 2088 586 2092
rect 566 2078 570 2082
rect 646 2078 650 2082
rect 262 2068 266 2072
rect 246 2058 250 2062
rect 270 2058 274 2062
rect 286 2058 290 2062
rect 302 2058 306 2062
rect 214 2048 218 2052
rect 294 2048 298 2052
rect 318 2048 322 2052
rect 158 2038 162 2042
rect 222 2038 226 2042
rect 230 2038 234 2042
rect 390 2038 394 2042
rect 30 1978 34 1982
rect 86 1978 90 1982
rect 38 1968 42 1972
rect 54 1958 58 1962
rect 78 1958 82 1962
rect 54 1948 58 1952
rect 94 1948 98 1952
rect 174 2028 178 2032
rect 206 1988 210 1992
rect 214 1978 218 1982
rect 254 1978 258 1982
rect 134 1968 138 1972
rect 230 1968 234 1972
rect 238 1968 242 1972
rect 270 1968 274 1972
rect 142 1958 146 1962
rect 454 2058 458 2062
rect 414 2048 418 2052
rect 422 2038 426 2042
rect 470 2038 474 2042
rect 454 2018 458 2022
rect 470 2018 474 2022
rect 494 2018 498 2022
rect 406 2008 410 2012
rect 346 2003 350 2007
rect 353 2003 357 2007
rect 398 1998 402 2002
rect 398 1968 402 1972
rect 302 1958 306 1962
rect 318 1958 322 1962
rect 390 1958 394 1962
rect 38 1938 42 1942
rect 62 1938 66 1942
rect 78 1938 82 1942
rect 30 1928 34 1932
rect 46 1928 50 1932
rect 70 1928 74 1932
rect 78 1928 82 1932
rect 62 1898 66 1902
rect 38 1838 42 1842
rect 110 1868 114 1872
rect 118 1868 122 1872
rect 62 1848 66 1852
rect 86 1858 90 1862
rect 102 1858 106 1862
rect 78 1838 82 1842
rect 6 1778 10 1782
rect 14 1778 18 1782
rect 22 1768 26 1772
rect 38 1768 42 1772
rect 30 1758 34 1762
rect 262 1948 266 1952
rect 206 1938 210 1942
rect 158 1908 162 1912
rect 166 1898 170 1902
rect 214 1928 218 1932
rect 206 1918 210 1922
rect 222 1918 226 1922
rect 198 1898 202 1902
rect 110 1848 114 1852
rect 158 1848 162 1852
rect 94 1838 98 1842
rect 150 1818 154 1822
rect 86 1788 90 1792
rect 126 1788 130 1792
rect 70 1778 74 1782
rect 94 1768 98 1772
rect 134 1768 138 1772
rect 94 1758 98 1762
rect 94 1748 98 1752
rect 126 1748 130 1752
rect 142 1748 146 1752
rect 62 1738 66 1742
rect 46 1688 50 1692
rect 134 1738 138 1742
rect 326 1948 330 1952
rect 350 1948 354 1952
rect 294 1938 298 1942
rect 334 1938 338 1942
rect 262 1928 266 1932
rect 310 1918 314 1922
rect 254 1908 258 1912
rect 238 1898 242 1902
rect 342 1908 346 1912
rect 238 1888 242 1892
rect 334 1888 338 1892
rect 222 1878 226 1882
rect 214 1868 218 1872
rect 270 1878 274 1882
rect 326 1878 330 1882
rect 342 1878 346 1882
rect 254 1868 258 1872
rect 294 1868 298 1872
rect 302 1868 306 1872
rect 198 1838 202 1842
rect 206 1838 210 1842
rect 182 1828 186 1832
rect 214 1828 218 1832
rect 174 1778 178 1782
rect 366 1948 370 1952
rect 382 1948 386 1952
rect 358 1908 362 1912
rect 446 1968 450 1972
rect 438 1958 442 1962
rect 430 1918 434 1922
rect 518 2058 522 2062
rect 518 2048 522 2052
rect 582 2068 586 2072
rect 574 2048 578 2052
rect 782 2158 786 2162
rect 774 2148 778 2152
rect 830 2148 834 2152
rect 1006 2338 1010 2342
rect 1006 2328 1010 2332
rect 1110 2458 1114 2462
rect 1118 2458 1122 2462
rect 1294 2478 1298 2482
rect 1302 2478 1306 2482
rect 1158 2458 1162 2462
rect 1206 2458 1210 2462
rect 1246 2458 1250 2462
rect 1262 2458 1266 2462
rect 1294 2458 1298 2462
rect 1206 2448 1210 2452
rect 1230 2448 1234 2452
rect 1294 2448 1298 2452
rect 1174 2438 1178 2442
rect 1278 2438 1282 2442
rect 1126 2398 1130 2402
rect 1062 2378 1066 2382
rect 1102 2378 1106 2382
rect 1118 2378 1122 2382
rect 1454 2708 1458 2712
rect 1430 2618 1434 2622
rect 1370 2603 1374 2607
rect 1377 2603 1381 2607
rect 1390 2548 1394 2552
rect 1382 2438 1386 2442
rect 1350 2428 1354 2432
rect 1326 2418 1330 2422
rect 1318 2378 1322 2382
rect 1182 2368 1186 2372
rect 1078 2358 1082 2362
rect 1062 2348 1066 2352
rect 1078 2348 1082 2352
rect 1174 2348 1178 2352
rect 1054 2338 1058 2342
rect 1126 2338 1130 2342
rect 1102 2328 1106 2332
rect 1046 2318 1050 2322
rect 1030 2308 1034 2312
rect 1030 2288 1034 2292
rect 1030 2248 1034 2252
rect 1014 2238 1018 2242
rect 990 2218 994 2222
rect 926 2178 930 2182
rect 950 2178 954 2182
rect 894 2148 898 2152
rect 934 2148 938 2152
rect 806 2138 810 2142
rect 830 2138 834 2142
rect 854 2138 858 2142
rect 910 2138 914 2142
rect 926 2138 930 2142
rect 942 2138 946 2142
rect 854 2128 858 2132
rect 858 2103 862 2107
rect 865 2103 869 2107
rect 806 2078 810 2082
rect 526 2008 530 2012
rect 502 1998 506 2002
rect 574 1998 578 2002
rect 462 1988 466 1992
rect 494 1988 498 1992
rect 502 1988 506 1992
rect 470 1958 474 1962
rect 470 1928 474 1932
rect 742 2038 746 2042
rect 694 2028 698 2032
rect 726 1988 730 1992
rect 582 1968 586 1972
rect 638 1968 642 1972
rect 526 1958 530 1962
rect 534 1958 538 1962
rect 574 1948 578 1952
rect 590 1948 594 1952
rect 518 1938 522 1942
rect 590 1938 594 1942
rect 510 1928 514 1932
rect 550 1928 554 1932
rect 614 1928 618 1932
rect 382 1888 386 1892
rect 366 1878 370 1882
rect 758 2028 762 2032
rect 782 1948 786 1952
rect 638 1938 642 1942
rect 646 1938 650 1942
rect 598 1918 602 1922
rect 630 1918 634 1922
rect 662 1908 666 1912
rect 526 1878 530 1882
rect 558 1878 562 1882
rect 694 1878 698 1882
rect 358 1868 362 1872
rect 446 1868 450 1872
rect 462 1868 466 1872
rect 670 1868 674 1872
rect 262 1858 266 1862
rect 286 1858 290 1862
rect 326 1858 330 1862
rect 438 1858 442 1862
rect 278 1848 282 1852
rect 246 1838 250 1842
rect 350 1838 354 1842
rect 346 1803 350 1807
rect 353 1803 357 1807
rect 334 1788 338 1792
rect 278 1768 282 1772
rect 294 1768 298 1772
rect 390 1768 394 1772
rect 414 1768 418 1772
rect 150 1738 154 1742
rect 182 1728 186 1732
rect 222 1718 226 1722
rect 198 1708 202 1712
rect 286 1758 290 1762
rect 310 1758 314 1762
rect 390 1758 394 1762
rect 398 1758 402 1762
rect 286 1748 290 1752
rect 334 1748 338 1752
rect 374 1748 378 1752
rect 262 1738 266 1742
rect 254 1708 258 1712
rect 110 1678 114 1682
rect 166 1678 170 1682
rect 22 1618 26 1622
rect 86 1568 90 1572
rect 62 1558 66 1562
rect 46 1548 50 1552
rect 14 1538 18 1542
rect 38 1518 42 1522
rect 38 1498 42 1502
rect 6 1458 10 1462
rect 46 1448 50 1452
rect 22 1428 26 1432
rect 22 1408 26 1412
rect 46 1408 50 1412
rect 46 1368 50 1372
rect 78 1538 82 1542
rect 166 1648 170 1652
rect 238 1648 242 1652
rect 158 1628 162 1632
rect 110 1588 114 1592
rect 158 1588 162 1592
rect 134 1568 138 1572
rect 158 1558 162 1562
rect 110 1538 114 1542
rect 134 1518 138 1522
rect 102 1508 106 1512
rect 158 1508 162 1512
rect 94 1488 98 1492
rect 70 1478 74 1482
rect 70 1458 74 1462
rect 102 1458 106 1462
rect 134 1458 138 1462
rect 62 1378 66 1382
rect 94 1378 98 1382
rect 126 1388 130 1392
rect 118 1378 122 1382
rect 46 1358 50 1362
rect 54 1358 58 1362
rect 86 1358 90 1362
rect 110 1358 114 1362
rect 70 1338 74 1342
rect 94 1338 98 1342
rect 62 1328 66 1332
rect 78 1328 82 1332
rect 118 1278 122 1282
rect 302 1678 306 1682
rect 654 1858 658 1862
rect 550 1848 554 1852
rect 638 1848 642 1852
rect 582 1838 586 1842
rect 782 1918 786 1922
rect 774 1878 778 1882
rect 726 1858 730 1862
rect 574 1778 578 1782
rect 462 1768 466 1772
rect 550 1768 554 1772
rect 406 1738 410 1742
rect 422 1738 426 1742
rect 438 1738 442 1742
rect 702 1798 706 1802
rect 742 1818 746 1822
rect 734 1808 738 1812
rect 726 1778 730 1782
rect 758 1788 762 1792
rect 742 1778 746 1782
rect 750 1778 754 1782
rect 686 1748 690 1752
rect 902 2058 906 2062
rect 926 2008 930 2012
rect 990 2118 994 2122
rect 1270 2348 1274 2352
rect 1166 2338 1170 2342
rect 1198 2338 1202 2342
rect 1182 2328 1186 2332
rect 1150 2308 1154 2312
rect 1126 2288 1130 2292
rect 1118 2278 1122 2282
rect 1166 2268 1170 2272
rect 1102 2248 1106 2252
rect 1278 2308 1282 2312
rect 1254 2288 1258 2292
rect 1246 2278 1250 2282
rect 1462 2598 1466 2602
rect 1518 2728 1522 2732
rect 1566 2858 1570 2862
rect 1614 2858 1618 2862
rect 1558 2848 1562 2852
rect 1630 2848 1634 2852
rect 1654 2878 1658 2882
rect 1806 2918 1810 2922
rect 1798 2888 1802 2892
rect 1694 2878 1698 2882
rect 1662 2868 1666 2872
rect 1710 2868 1714 2872
rect 1662 2858 1666 2862
rect 1718 2858 1722 2862
rect 1678 2848 1682 2852
rect 1734 2848 1738 2852
rect 1542 2768 1546 2772
rect 1654 2828 1658 2832
rect 1582 2758 1586 2762
rect 1646 2798 1650 2802
rect 1806 2868 1810 2872
rect 1874 2903 1878 2907
rect 1881 2903 1885 2907
rect 1870 2888 1874 2892
rect 1918 2928 1922 2932
rect 2006 2958 2010 2962
rect 2030 2968 2034 2972
rect 2038 2958 2042 2962
rect 1982 2948 1986 2952
rect 2030 2948 2034 2952
rect 2046 2948 2050 2952
rect 1950 2938 1954 2942
rect 1942 2928 1946 2932
rect 1926 2918 1930 2922
rect 1990 2918 1994 2922
rect 2230 3108 2234 3112
rect 2246 3108 2250 3112
rect 2126 3078 2130 3082
rect 2182 3078 2186 3082
rect 2222 3078 2226 3082
rect 2350 3178 2354 3182
rect 2326 3158 2330 3162
rect 2342 3158 2346 3162
rect 2318 3148 2322 3152
rect 2302 3138 2306 3142
rect 2294 3128 2298 3132
rect 2302 3108 2306 3112
rect 2374 3278 2378 3282
rect 2414 3348 2418 3352
rect 2430 3348 2434 3352
rect 2494 3448 2498 3452
rect 2526 3508 2530 3512
rect 2670 3548 2674 3552
rect 2638 3538 2642 3542
rect 2678 3538 2682 3542
rect 2590 3528 2594 3532
rect 2630 3528 2634 3532
rect 2574 3488 2578 3492
rect 2598 3518 2602 3522
rect 2622 3498 2626 3502
rect 2614 3478 2618 3482
rect 2518 3438 2522 3442
rect 2510 3408 2514 3412
rect 2478 3398 2482 3402
rect 2486 3358 2490 3362
rect 2462 3348 2466 3352
rect 2526 3388 2530 3392
rect 2582 3458 2586 3462
rect 2542 3448 2546 3452
rect 2558 3438 2562 3442
rect 2534 3378 2538 3382
rect 2654 3528 2658 3532
rect 2694 3528 2698 3532
rect 2646 3488 2650 3492
rect 2614 3458 2618 3462
rect 2638 3458 2642 3462
rect 2662 3518 2666 3522
rect 2718 3548 2722 3552
rect 2782 3558 2786 3562
rect 2734 3518 2738 3522
rect 2822 3548 2826 3552
rect 2854 3548 2858 3552
rect 3022 3588 3026 3592
rect 2950 3568 2954 3572
rect 2966 3548 2970 3552
rect 3014 3548 3018 3552
rect 2830 3538 2834 3542
rect 2846 3538 2850 3542
rect 2918 3538 2922 3542
rect 2766 3528 2770 3532
rect 2822 3528 2826 3532
rect 2958 3528 2962 3532
rect 2990 3528 2994 3532
rect 2750 3518 2754 3522
rect 2726 3508 2730 3512
rect 2742 3508 2746 3512
rect 2702 3488 2706 3492
rect 2814 3508 2818 3512
rect 2766 3498 2770 3502
rect 2726 3478 2730 3482
rect 2886 3518 2890 3522
rect 2906 3503 2910 3507
rect 2913 3503 2917 3507
rect 2878 3498 2882 3502
rect 2910 3488 2914 3492
rect 2950 3488 2954 3492
rect 2966 3488 2970 3492
rect 2870 3478 2874 3482
rect 2902 3478 2906 3482
rect 2958 3478 2962 3482
rect 2694 3468 2698 3472
rect 2726 3468 2730 3472
rect 2630 3408 2634 3412
rect 2622 3398 2626 3402
rect 2590 3378 2594 3382
rect 2750 3448 2754 3452
rect 2686 3428 2690 3432
rect 2726 3428 2730 3432
rect 2726 3398 2730 3402
rect 2678 3388 2682 3392
rect 2662 3378 2666 3382
rect 2574 3368 2578 3372
rect 2582 3368 2586 3372
rect 2526 3348 2530 3352
rect 2574 3348 2578 3352
rect 2390 3338 2394 3342
rect 2502 3338 2506 3342
rect 2518 3338 2522 3342
rect 2550 3338 2554 3342
rect 2566 3338 2570 3342
rect 2486 3328 2490 3332
rect 2502 3328 2506 3332
rect 2598 3348 2602 3352
rect 2590 3328 2594 3332
rect 2606 3328 2610 3332
rect 2446 3278 2450 3282
rect 2406 3258 2410 3262
rect 2430 3248 2434 3252
rect 2390 3238 2394 3242
rect 2462 3288 2466 3292
rect 2534 3278 2538 3282
rect 2718 3368 2722 3372
rect 2622 3358 2626 3362
rect 2638 3358 2642 3362
rect 2702 3358 2706 3362
rect 2654 3348 2658 3352
rect 2702 3348 2706 3352
rect 2646 3338 2650 3342
rect 2686 3338 2690 3342
rect 2742 3368 2746 3372
rect 2974 3468 2978 3472
rect 3006 3528 3010 3532
rect 3038 3558 3042 3562
rect 3062 3558 3066 3562
rect 3118 3648 3122 3652
rect 3118 3558 3122 3562
rect 3046 3538 3050 3542
rect 3078 3538 3082 3542
rect 2918 3458 2922 3462
rect 2958 3458 2962 3462
rect 2966 3458 2970 3462
rect 2982 3458 2986 3462
rect 2998 3458 3002 3462
rect 2790 3438 2794 3442
rect 2830 3438 2834 3442
rect 2766 3378 2770 3382
rect 2758 3358 2762 3362
rect 2814 3358 2818 3362
rect 2846 3428 2850 3432
rect 2846 3368 2850 3372
rect 2862 3368 2866 3372
rect 2830 3348 2834 3352
rect 2726 3338 2730 3342
rect 2646 3328 2650 3332
rect 2678 3328 2682 3332
rect 2726 3288 2730 3292
rect 2622 3278 2626 3282
rect 2686 3278 2690 3282
rect 2558 3268 2562 3272
rect 2590 3268 2594 3272
rect 2614 3268 2618 3272
rect 2630 3268 2634 3272
rect 2670 3268 2674 3272
rect 2478 3258 2482 3262
rect 2510 3258 2514 3262
rect 2494 3248 2498 3252
rect 2518 3248 2522 3252
rect 2550 3238 2554 3242
rect 2454 3228 2458 3232
rect 2478 3218 2482 3222
rect 2394 3203 2398 3207
rect 2401 3203 2405 3207
rect 2446 3188 2450 3192
rect 2374 3178 2378 3182
rect 2390 3158 2394 3162
rect 2382 3148 2386 3152
rect 2390 3148 2394 3152
rect 2358 3128 2362 3132
rect 2486 3168 2490 3172
rect 2398 3108 2402 3112
rect 2446 3108 2450 3112
rect 2550 3158 2554 3162
rect 2502 3148 2506 3152
rect 2526 3148 2530 3152
rect 2566 3258 2570 3262
rect 2646 3258 2650 3262
rect 2654 3258 2658 3262
rect 2614 3228 2618 3232
rect 2718 3268 2722 3272
rect 2710 3248 2714 3252
rect 2742 3248 2746 3252
rect 2678 3228 2682 3232
rect 2670 3208 2674 3212
rect 2654 3178 2658 3182
rect 2494 3138 2498 3142
rect 2622 3138 2626 3142
rect 2510 3118 2514 3122
rect 2334 3088 2338 3092
rect 2358 3088 2362 3092
rect 2326 3078 2330 3082
rect 2342 3068 2346 3072
rect 2366 3078 2370 3082
rect 2518 3078 2522 3082
rect 2638 3128 2642 3132
rect 2702 3208 2706 3212
rect 2710 3188 2714 3192
rect 2670 3158 2674 3162
rect 2686 3158 2690 3162
rect 2774 3338 2778 3342
rect 2838 3338 2842 3342
rect 2782 3328 2786 3332
rect 2830 3328 2834 3332
rect 2774 3318 2778 3322
rect 2790 3268 2794 3272
rect 2814 3268 2818 3272
rect 2926 3448 2930 3452
rect 3118 3538 3122 3542
rect 3110 3498 3114 3502
rect 3086 3488 3090 3492
rect 3110 3488 3114 3492
rect 3078 3468 3082 3472
rect 3014 3448 3018 3452
rect 2958 3398 2962 3402
rect 2862 3358 2866 3362
rect 2886 3358 2890 3362
rect 2894 3358 2898 3362
rect 2950 3358 2954 3362
rect 2990 3358 2994 3362
rect 2870 3288 2874 3292
rect 2846 3268 2850 3272
rect 2854 3268 2858 3272
rect 2766 3258 2770 3262
rect 2790 3248 2794 3252
rect 2822 3248 2826 3252
rect 2766 3228 2770 3232
rect 2814 3198 2818 3202
rect 2894 3338 2898 3342
rect 2974 3338 2978 3342
rect 2982 3338 2986 3342
rect 3006 3338 3010 3342
rect 2966 3318 2970 3322
rect 3014 3318 3018 3322
rect 2906 3303 2910 3307
rect 2913 3303 2917 3307
rect 3038 3458 3042 3462
rect 3054 3438 3058 3442
rect 3158 3618 3162 3622
rect 3142 3538 3146 3542
rect 3134 3528 3138 3532
rect 3126 3488 3130 3492
rect 3222 3638 3226 3642
rect 3278 3618 3282 3622
rect 3302 3618 3306 3622
rect 3190 3568 3194 3572
rect 3198 3568 3202 3572
rect 3198 3558 3202 3562
rect 3374 3658 3378 3662
rect 3326 3648 3330 3652
rect 3438 3618 3442 3622
rect 3398 3608 3402 3612
rect 3350 3558 3354 3562
rect 3418 3603 3422 3607
rect 3425 3603 3429 3607
rect 3326 3548 3330 3552
rect 3446 3548 3450 3552
rect 3454 3548 3458 3552
rect 3182 3528 3186 3532
rect 3174 3508 3178 3512
rect 3158 3488 3162 3492
rect 3142 3458 3146 3462
rect 3118 3448 3122 3452
rect 3126 3448 3130 3452
rect 3190 3498 3194 3502
rect 3270 3478 3274 3482
rect 3166 3468 3170 3472
rect 3150 3438 3154 3442
rect 3030 3428 3034 3432
rect 3046 3428 3050 3432
rect 3062 3428 3066 3432
rect 3102 3428 3106 3432
rect 3134 3418 3138 3422
rect 3046 3378 3050 3382
rect 3062 3378 3066 3382
rect 3030 3368 3034 3372
rect 3046 3348 3050 3352
rect 2974 3288 2978 3292
rect 3022 3288 3026 3292
rect 2950 3278 2954 3282
rect 2998 3278 3002 3282
rect 3022 3278 3026 3282
rect 2894 3268 2898 3272
rect 2934 3268 2938 3272
rect 2966 3268 2970 3272
rect 3022 3268 3026 3272
rect 2918 3258 2922 3262
rect 2902 3228 2906 3232
rect 2894 3218 2898 3222
rect 2822 3188 2826 3192
rect 2838 3188 2842 3192
rect 2798 3168 2802 3172
rect 2806 3168 2810 3172
rect 2838 3168 2842 3172
rect 2854 3168 2858 3172
rect 2886 3168 2890 3172
rect 2766 3158 2770 3162
rect 2758 3148 2762 3152
rect 2678 3138 2682 3142
rect 2702 3138 2706 3142
rect 2734 3138 2738 3142
rect 2774 3148 2778 3152
rect 2814 3138 2818 3142
rect 2718 3128 2722 3132
rect 2742 3128 2746 3132
rect 3078 3348 3082 3352
rect 3094 3338 3098 3342
rect 3126 3338 3130 3342
rect 3062 3328 3066 3332
rect 3110 3328 3114 3332
rect 3126 3328 3130 3332
rect 3094 3298 3098 3302
rect 3062 3288 3066 3292
rect 3102 3288 3106 3292
rect 3110 3278 3114 3282
rect 3086 3268 3090 3272
rect 2934 3248 2938 3252
rect 2958 3248 2962 3252
rect 2998 3258 3002 3262
rect 3030 3258 3034 3262
rect 2966 3168 2970 3172
rect 2942 3158 2946 3162
rect 3142 3268 3146 3272
rect 3126 3258 3130 3262
rect 3054 3248 3058 3252
rect 3062 3248 3066 3252
rect 3038 3238 3042 3242
rect 3078 3238 3082 3242
rect 3094 3238 3098 3242
rect 3006 3178 3010 3182
rect 2982 3148 2986 3152
rect 2662 3118 2666 3122
rect 2710 3118 2714 3122
rect 2718 3108 2722 3112
rect 2830 3118 2834 3122
rect 2750 3088 2754 3092
rect 2798 3088 2802 3092
rect 2446 3068 2450 3072
rect 2622 3068 2626 3072
rect 2678 3068 2682 3072
rect 2710 3068 2714 3072
rect 2718 3068 2722 3072
rect 2158 3058 2162 3062
rect 2198 3058 2202 3062
rect 2246 3058 2250 3062
rect 2350 3058 2354 3062
rect 2382 3058 2386 3062
rect 2566 3058 2570 3062
rect 2598 3058 2602 3062
rect 2654 3058 2658 3062
rect 2694 3058 2698 3062
rect 2230 3048 2234 3052
rect 2254 3048 2258 3052
rect 2422 3048 2426 3052
rect 2646 3048 2650 3052
rect 2118 3038 2122 3042
rect 2366 3038 2370 3042
rect 2582 3038 2586 3042
rect 2070 2998 2074 3002
rect 2062 2988 2066 2992
rect 2062 2958 2066 2962
rect 2150 2998 2154 3002
rect 2078 2988 2082 2992
rect 2118 2988 2122 2992
rect 2086 2978 2090 2982
rect 2166 2978 2170 2982
rect 2110 2958 2114 2962
rect 2126 2958 2130 2962
rect 2230 2978 2234 2982
rect 2158 2958 2162 2962
rect 2198 2958 2202 2962
rect 2214 2958 2218 2962
rect 2086 2948 2090 2952
rect 2110 2948 2114 2952
rect 2150 2948 2154 2952
rect 2182 2948 2186 2952
rect 2134 2938 2138 2942
rect 2158 2938 2162 2942
rect 2222 2948 2226 2952
rect 2158 2928 2162 2932
rect 2414 3018 2418 3022
rect 2394 3003 2398 3007
rect 2401 3003 2405 3007
rect 2390 2988 2394 2992
rect 2286 2978 2290 2982
rect 2262 2968 2266 2972
rect 2310 2968 2314 2972
rect 2286 2958 2290 2962
rect 2294 2958 2298 2962
rect 2238 2948 2242 2952
rect 2246 2938 2250 2942
rect 2278 2938 2282 2942
rect 2906 3103 2910 3107
rect 2913 3103 2917 3107
rect 2950 3098 2954 3102
rect 2982 3098 2986 3102
rect 2950 3078 2954 3082
rect 2974 3078 2978 3082
rect 2846 3068 2850 3072
rect 2862 3068 2866 3072
rect 2966 3068 2970 3072
rect 2806 3058 2810 3062
rect 2774 3028 2778 3032
rect 2902 3058 2906 3062
rect 2862 3048 2866 3052
rect 2878 3048 2882 3052
rect 2758 3008 2762 3012
rect 2838 3008 2842 3012
rect 2854 3008 2858 3012
rect 2638 2978 2642 2982
rect 2558 2968 2562 2972
rect 2462 2958 2466 2962
rect 2526 2958 2530 2962
rect 2582 2958 2586 2962
rect 2614 2958 2618 2962
rect 2622 2958 2626 2962
rect 2422 2938 2426 2942
rect 2318 2928 2322 2932
rect 2294 2908 2298 2912
rect 2070 2898 2074 2902
rect 2126 2898 2130 2902
rect 2142 2898 2146 2902
rect 1918 2888 1922 2892
rect 1950 2888 1954 2892
rect 2030 2888 2034 2892
rect 2038 2888 2042 2892
rect 2054 2888 2058 2892
rect 2102 2888 2106 2892
rect 1894 2878 1898 2882
rect 1830 2868 1834 2872
rect 1846 2868 1850 2872
rect 1982 2868 1986 2872
rect 1758 2858 1762 2862
rect 1798 2858 1802 2862
rect 1774 2848 1778 2852
rect 1766 2838 1770 2842
rect 1742 2828 1746 2832
rect 1654 2778 1658 2782
rect 1702 2768 1706 2772
rect 1758 2768 1762 2772
rect 1542 2748 1546 2752
rect 1566 2748 1570 2752
rect 1606 2748 1610 2752
rect 1550 2738 1554 2742
rect 1526 2688 1530 2692
rect 1502 2588 1506 2592
rect 1518 2558 1522 2562
rect 1542 2518 1546 2522
rect 1526 2498 1530 2502
rect 1438 2488 1442 2492
rect 1422 2408 1426 2412
rect 1370 2403 1374 2407
rect 1377 2403 1381 2407
rect 1390 2368 1394 2372
rect 1350 2338 1354 2342
rect 1390 2318 1394 2322
rect 1342 2298 1346 2302
rect 1390 2298 1394 2302
rect 1286 2278 1290 2282
rect 1446 2478 1450 2482
rect 1518 2468 1522 2472
rect 1518 2438 1522 2442
rect 1462 2358 1466 2362
rect 1478 2358 1482 2362
rect 1502 2348 1506 2352
rect 1518 2318 1522 2322
rect 1590 2698 1594 2702
rect 1670 2758 1674 2762
rect 1726 2748 1730 2752
rect 1846 2848 1850 2852
rect 1942 2858 1946 2862
rect 1974 2858 1978 2862
rect 1862 2848 1866 2852
rect 1902 2848 1906 2852
rect 1814 2838 1818 2842
rect 1854 2838 1858 2842
rect 1790 2818 1794 2822
rect 1782 2798 1786 2802
rect 1998 2838 2002 2842
rect 2006 2838 2010 2842
rect 1926 2828 1930 2832
rect 1878 2798 1882 2802
rect 1838 2788 1842 2792
rect 1822 2778 1826 2782
rect 1838 2778 1842 2782
rect 1830 2768 1834 2772
rect 1830 2758 1834 2762
rect 1838 2758 1842 2762
rect 1774 2748 1778 2752
rect 1710 2738 1714 2742
rect 1782 2738 1786 2742
rect 1814 2738 1818 2742
rect 1670 2728 1674 2732
rect 1726 2728 1730 2732
rect 1902 2788 1906 2792
rect 1918 2778 1922 2782
rect 1910 2748 1914 2752
rect 1934 2798 1938 2802
rect 2062 2878 2066 2882
rect 2078 2868 2082 2872
rect 2262 2888 2266 2892
rect 2142 2878 2146 2882
rect 2166 2878 2170 2882
rect 2174 2878 2178 2882
rect 2110 2868 2114 2872
rect 2158 2868 2162 2872
rect 2046 2858 2050 2862
rect 2094 2858 2098 2862
rect 2126 2858 2130 2862
rect 2038 2838 2042 2842
rect 2054 2838 2058 2842
rect 2062 2838 2066 2842
rect 2174 2868 2178 2872
rect 2342 2908 2346 2912
rect 2302 2898 2306 2902
rect 2302 2878 2306 2882
rect 2334 2878 2338 2882
rect 2334 2868 2338 2872
rect 2510 2948 2514 2952
rect 2422 2878 2426 2882
rect 2382 2868 2386 2872
rect 2198 2858 2202 2862
rect 2246 2858 2250 2862
rect 2286 2858 2290 2862
rect 2358 2858 2362 2862
rect 2318 2848 2322 2852
rect 2334 2848 2338 2852
rect 2150 2838 2154 2842
rect 2190 2838 2194 2842
rect 2094 2828 2098 2832
rect 2022 2818 2026 2822
rect 2182 2818 2186 2822
rect 2230 2818 2234 2822
rect 2054 2798 2058 2802
rect 2118 2788 2122 2792
rect 1974 2778 1978 2782
rect 2222 2778 2226 2782
rect 1958 2768 1962 2772
rect 1950 2758 1954 2762
rect 1942 2748 1946 2752
rect 1934 2738 1938 2742
rect 1910 2728 1914 2732
rect 1958 2728 1962 2732
rect 1710 2718 1714 2722
rect 1742 2718 1746 2722
rect 1630 2678 1634 2682
rect 1598 2668 1602 2672
rect 1654 2658 1658 2662
rect 1614 2538 1618 2542
rect 1798 2718 1802 2722
rect 1998 2768 2002 2772
rect 2022 2768 2026 2772
rect 1998 2758 2002 2762
rect 2006 2758 2010 2762
rect 2142 2758 2146 2762
rect 2070 2748 2074 2752
rect 2046 2738 2050 2742
rect 1782 2708 1786 2712
rect 1934 2708 1938 2712
rect 1966 2708 1970 2712
rect 2038 2708 2042 2712
rect 1758 2688 1762 2692
rect 1718 2678 1722 2682
rect 1670 2648 1674 2652
rect 1702 2648 1706 2652
rect 1702 2638 1706 2642
rect 1694 2628 1698 2632
rect 1662 2568 1666 2572
rect 1686 2538 1690 2542
rect 1734 2598 1738 2602
rect 1750 2598 1754 2602
rect 1678 2528 1682 2532
rect 1646 2518 1650 2522
rect 1606 2478 1610 2482
rect 1678 2468 1682 2472
rect 1678 2458 1682 2462
rect 1550 2438 1554 2442
rect 1574 2438 1578 2442
rect 1566 2428 1570 2432
rect 1598 2428 1602 2432
rect 1614 2428 1618 2432
rect 1566 2378 1570 2382
rect 1662 2358 1666 2362
rect 1582 2348 1586 2352
rect 1670 2348 1674 2352
rect 1750 2528 1754 2532
rect 1718 2508 1722 2512
rect 1718 2468 1722 2472
rect 1734 2459 1738 2463
rect 1758 2458 1762 2462
rect 1710 2408 1714 2412
rect 1774 2428 1778 2432
rect 1758 2398 1762 2402
rect 1710 2378 1714 2382
rect 1726 2378 1730 2382
rect 1750 2378 1754 2382
rect 1694 2368 1698 2372
rect 1742 2368 1746 2372
rect 1726 2358 1730 2362
rect 1766 2358 1770 2362
rect 1718 2348 1722 2352
rect 1638 2338 1642 2342
rect 1558 2318 1562 2322
rect 1526 2308 1530 2312
rect 1478 2298 1482 2302
rect 1494 2298 1498 2302
rect 1502 2298 1506 2302
rect 1518 2298 1522 2302
rect 1350 2268 1354 2272
rect 1542 2268 1546 2272
rect 1558 2268 1562 2272
rect 1566 2268 1570 2272
rect 1286 2258 1290 2262
rect 1198 2248 1202 2252
rect 1182 2218 1186 2222
rect 1182 2188 1186 2192
rect 1342 2258 1346 2262
rect 1062 2158 1066 2162
rect 1158 2158 1162 2162
rect 1286 2158 1290 2162
rect 1334 2158 1338 2162
rect 1382 2258 1386 2262
rect 1398 2258 1402 2262
rect 1406 2238 1410 2242
rect 1370 2203 1374 2207
rect 1377 2203 1381 2207
rect 1430 2258 1434 2262
rect 1438 2218 1442 2222
rect 1414 2198 1418 2202
rect 1510 2258 1514 2262
rect 1550 2258 1554 2262
rect 1566 2248 1570 2252
rect 1470 2238 1474 2242
rect 1462 2198 1466 2202
rect 1526 2218 1530 2222
rect 1542 2208 1546 2212
rect 1470 2178 1474 2182
rect 1542 2178 1546 2182
rect 1566 2178 1570 2182
rect 1542 2158 1546 2162
rect 1246 2147 1250 2151
rect 1358 2148 1362 2152
rect 1390 2148 1394 2152
rect 1422 2148 1426 2152
rect 1486 2148 1490 2152
rect 1502 2148 1506 2152
rect 1150 2138 1154 2142
rect 1222 2138 1226 2142
rect 1078 2128 1082 2132
rect 1094 2128 1098 2132
rect 1046 2108 1050 2112
rect 1086 2098 1090 2102
rect 1022 2078 1026 2082
rect 1030 2078 1034 2082
rect 1214 2108 1218 2112
rect 1054 2078 1058 2082
rect 1070 2078 1074 2082
rect 950 2068 954 2072
rect 1014 2068 1018 2072
rect 958 2058 962 2062
rect 1022 2058 1026 2062
rect 1270 2088 1274 2092
rect 1262 2078 1266 2082
rect 1070 2048 1074 2052
rect 1078 2048 1082 2052
rect 1118 2038 1122 2042
rect 942 1978 946 1982
rect 870 1968 874 1972
rect 902 1968 906 1972
rect 934 1968 938 1972
rect 990 1968 994 1972
rect 822 1958 826 1962
rect 830 1948 834 1952
rect 838 1938 842 1942
rect 910 1958 914 1962
rect 934 1958 938 1962
rect 942 1958 946 1962
rect 990 1958 994 1962
rect 918 1948 922 1952
rect 886 1938 890 1942
rect 926 1938 930 1942
rect 858 1903 862 1907
rect 865 1903 869 1907
rect 822 1888 826 1892
rect 838 1888 842 1892
rect 870 1888 874 1892
rect 886 1888 890 1892
rect 918 1888 922 1892
rect 798 1828 802 1832
rect 790 1818 794 1822
rect 814 1818 818 1822
rect 798 1808 802 1812
rect 918 1868 922 1872
rect 886 1858 890 1862
rect 846 1798 850 1802
rect 894 1778 898 1782
rect 958 1928 962 1932
rect 1182 2048 1186 2052
rect 1246 2048 1250 2052
rect 1278 2048 1282 2052
rect 1150 2028 1154 2032
rect 1358 2138 1362 2142
rect 1334 2118 1338 2122
rect 1502 2128 1506 2132
rect 1486 2118 1490 2122
rect 1470 2108 1474 2112
rect 1494 2098 1498 2102
rect 1414 2088 1418 2092
rect 1478 2088 1482 2092
rect 1310 2068 1314 2072
rect 1334 2068 1338 2072
rect 1342 2068 1346 2072
rect 1302 2018 1306 2022
rect 1150 1988 1154 1992
rect 1294 1988 1298 1992
rect 1206 1978 1210 1982
rect 1054 1968 1058 1972
rect 1078 1968 1082 1972
rect 1118 1968 1122 1972
rect 1150 1968 1154 1972
rect 1022 1948 1026 1952
rect 1038 1948 1042 1952
rect 1062 1948 1066 1952
rect 990 1938 994 1942
rect 1006 1938 1010 1942
rect 1046 1938 1050 1942
rect 1110 1958 1114 1962
rect 1134 1948 1138 1952
rect 1166 1948 1170 1952
rect 1086 1938 1090 1942
rect 1102 1938 1106 1942
rect 974 1928 978 1932
rect 1014 1928 1018 1932
rect 1158 1928 1162 1932
rect 1262 1968 1266 1972
rect 1222 1958 1226 1962
rect 1254 1958 1258 1962
rect 998 1878 1002 1882
rect 1054 1878 1058 1882
rect 1286 1958 1290 1962
rect 1318 1958 1322 1962
rect 1286 1948 1290 1952
rect 1310 1948 1314 1952
rect 1278 1938 1282 1942
rect 1294 1938 1298 1942
rect 1318 1938 1322 1942
rect 1334 1938 1338 1942
rect 1438 2058 1442 2062
rect 1390 2018 1394 2022
rect 1370 2003 1374 2007
rect 1377 2003 1381 2007
rect 1534 2088 1538 2092
rect 1518 2078 1522 2082
rect 1462 2058 1466 2062
rect 1478 2038 1482 2042
rect 1350 1988 1354 1992
rect 1446 1988 1450 1992
rect 1414 1978 1418 1982
rect 1558 2148 1562 2152
rect 1574 2138 1578 2142
rect 1630 2308 1634 2312
rect 1622 2298 1626 2302
rect 1598 2288 1602 2292
rect 1606 2288 1610 2292
rect 1598 2278 1602 2282
rect 1598 2268 1602 2272
rect 1590 2258 1594 2262
rect 1614 2168 1618 2172
rect 1590 2148 1594 2152
rect 1558 2078 1562 2082
rect 1566 2068 1570 2072
rect 1558 2058 1562 2062
rect 1566 2058 1570 2062
rect 1558 2018 1562 2022
rect 1502 1968 1506 1972
rect 1582 2088 1586 2092
rect 1590 2078 1594 2082
rect 1582 2068 1586 2072
rect 1582 2058 1586 2062
rect 1574 2048 1578 2052
rect 1566 1988 1570 1992
rect 1574 1978 1578 1982
rect 1638 2248 1642 2252
rect 1742 2328 1746 2332
rect 1710 2308 1714 2312
rect 1734 2298 1738 2302
rect 1718 2278 1722 2282
rect 1874 2703 1878 2707
rect 1881 2703 1885 2707
rect 1798 2698 1802 2702
rect 1894 2698 1898 2702
rect 1934 2688 1938 2692
rect 2054 2728 2058 2732
rect 2118 2728 2122 2732
rect 2126 2718 2130 2722
rect 2078 2708 2082 2712
rect 2102 2698 2106 2702
rect 2070 2688 2074 2692
rect 1814 2678 1818 2682
rect 1926 2678 1930 2682
rect 2046 2678 2050 2682
rect 1830 2668 1834 2672
rect 1982 2668 1986 2672
rect 1918 2658 1922 2662
rect 1934 2658 1938 2662
rect 1958 2658 1962 2662
rect 1990 2658 1994 2662
rect 2014 2666 2018 2670
rect 2062 2668 2066 2672
rect 2174 2748 2178 2752
rect 2254 2788 2258 2792
rect 2302 2788 2306 2792
rect 2342 2838 2346 2842
rect 2366 2838 2370 2842
rect 2366 2828 2370 2832
rect 2394 2803 2398 2807
rect 2401 2803 2405 2807
rect 2374 2798 2378 2802
rect 2342 2768 2346 2772
rect 2374 2768 2378 2772
rect 2246 2758 2250 2762
rect 2310 2758 2314 2762
rect 2326 2758 2330 2762
rect 2342 2758 2346 2762
rect 2374 2758 2378 2762
rect 2398 2758 2402 2762
rect 2350 2748 2354 2752
rect 2366 2748 2370 2752
rect 2414 2748 2418 2752
rect 2214 2678 2218 2682
rect 2094 2668 2098 2672
rect 2086 2658 2090 2662
rect 2126 2658 2130 2662
rect 2166 2668 2170 2672
rect 2174 2658 2178 2662
rect 2238 2658 2242 2662
rect 1990 2648 1994 2652
rect 1998 2648 2002 2652
rect 2038 2648 2042 2652
rect 2134 2648 2138 2652
rect 2206 2648 2210 2652
rect 2342 2708 2346 2712
rect 2454 2848 2458 2852
rect 2518 2938 2522 2942
rect 2590 2938 2594 2942
rect 2614 2938 2618 2942
rect 2630 2938 2634 2942
rect 2590 2928 2594 2932
rect 2614 2908 2618 2912
rect 2566 2888 2570 2892
rect 2934 3008 2938 3012
rect 3158 3428 3162 3432
rect 3254 3448 3258 3452
rect 3286 3428 3290 3432
rect 3182 3408 3186 3412
rect 3206 3388 3210 3392
rect 3214 3378 3218 3382
rect 3270 3378 3274 3382
rect 3198 3368 3202 3372
rect 3174 3358 3178 3362
rect 3198 3358 3202 3362
rect 3190 3348 3194 3352
rect 3166 3328 3170 3332
rect 3190 3338 3194 3342
rect 3158 3288 3162 3292
rect 3166 3248 3170 3252
rect 3230 3358 3234 3362
rect 3246 3358 3250 3362
rect 3318 3408 3322 3412
rect 3262 3338 3266 3342
rect 3302 3338 3306 3342
rect 3222 3328 3226 3332
rect 3206 3278 3210 3282
rect 3198 3258 3202 3262
rect 3182 3238 3186 3242
rect 3166 3218 3170 3222
rect 3102 3208 3106 3212
rect 3150 3208 3154 3212
rect 3174 3208 3178 3212
rect 3030 3158 3034 3162
rect 3014 3148 3018 3152
rect 3094 3148 3098 3152
rect 3294 3288 3298 3292
rect 3286 3278 3290 3282
rect 3342 3498 3346 3502
rect 3422 3538 3426 3542
rect 3358 3488 3362 3492
rect 3366 3488 3370 3492
rect 3358 3478 3362 3482
rect 3342 3398 3346 3402
rect 3334 3388 3338 3392
rect 3654 3658 3658 3662
rect 3694 3658 3698 3662
rect 3558 3648 3562 3652
rect 3582 3638 3586 3642
rect 3494 3628 3498 3632
rect 3654 3628 3658 3632
rect 3598 3618 3602 3622
rect 3622 3618 3626 3622
rect 3638 3618 3642 3622
rect 3638 3558 3642 3562
rect 3622 3548 3626 3552
rect 3646 3548 3650 3552
rect 3446 3468 3450 3472
rect 3502 3508 3506 3512
rect 3582 3528 3586 3532
rect 3614 3528 3618 3532
rect 3566 3518 3570 3522
rect 3630 3518 3634 3522
rect 3662 3528 3666 3532
rect 3670 3518 3674 3522
rect 3678 3518 3682 3522
rect 3478 3498 3482 3502
rect 3534 3498 3538 3502
rect 3606 3498 3610 3502
rect 3462 3478 3466 3482
rect 3670 3508 3674 3512
rect 3694 3508 3698 3512
rect 3638 3478 3642 3482
rect 3638 3468 3642 3472
rect 3398 3458 3402 3462
rect 3630 3458 3634 3462
rect 3574 3448 3578 3452
rect 3590 3448 3594 3452
rect 3542 3408 3546 3412
rect 3418 3403 3422 3407
rect 3425 3403 3429 3407
rect 3566 3388 3570 3392
rect 3542 3368 3546 3372
rect 3630 3368 3634 3372
rect 3750 3648 3754 3652
rect 3758 3648 3762 3652
rect 3758 3618 3762 3622
rect 3710 3538 3714 3542
rect 3702 3498 3706 3502
rect 3686 3488 3690 3492
rect 3734 3538 3738 3542
rect 3758 3538 3762 3542
rect 3726 3528 3730 3532
rect 3718 3518 3722 3522
rect 3718 3478 3722 3482
rect 3686 3458 3690 3462
rect 3702 3448 3706 3452
rect 3930 3703 3934 3707
rect 3937 3703 3941 3707
rect 3958 3698 3962 3702
rect 3998 3698 4002 3702
rect 4078 3698 4082 3702
rect 3806 3688 3810 3692
rect 3862 3688 3866 3692
rect 4086 3688 4090 3692
rect 3854 3678 3858 3682
rect 4054 3678 4058 3682
rect 4102 3678 4106 3682
rect 3958 3668 3962 3672
rect 3846 3658 3850 3662
rect 3822 3648 3826 3652
rect 3862 3638 3866 3642
rect 3806 3568 3810 3572
rect 3886 3558 3890 3562
rect 4006 3648 4010 3652
rect 4094 3668 4098 3672
rect 4086 3658 4090 3662
rect 4110 3648 4114 3652
rect 3950 3638 3954 3642
rect 3966 3638 3970 3642
rect 3982 3638 3986 3642
rect 4070 3638 4074 3642
rect 3910 3628 3914 3632
rect 3910 3568 3914 3572
rect 3822 3548 3826 3552
rect 3886 3548 3890 3552
rect 3902 3548 3906 3552
rect 3846 3538 3850 3542
rect 3886 3518 3890 3522
rect 3814 3508 3818 3512
rect 3870 3508 3874 3512
rect 3782 3478 3786 3482
rect 3838 3478 3842 3482
rect 3774 3438 3778 3442
rect 3726 3398 3730 3402
rect 3766 3398 3770 3402
rect 3718 3348 3722 3352
rect 3438 3338 3442 3342
rect 3478 3338 3482 3342
rect 3358 3298 3362 3302
rect 3310 3288 3314 3292
rect 3326 3288 3330 3292
rect 3358 3278 3362 3282
rect 3294 3268 3298 3272
rect 3254 3258 3258 3262
rect 3286 3258 3290 3262
rect 3270 3248 3274 3252
rect 3198 3238 3202 3242
rect 3214 3238 3218 3242
rect 3246 3238 3250 3242
rect 3222 3208 3226 3212
rect 3286 3218 3290 3222
rect 3190 3188 3194 3192
rect 3278 3188 3282 3192
rect 3254 3178 3258 3182
rect 3134 3158 3138 3162
rect 3174 3158 3178 3162
rect 3230 3158 3234 3162
rect 3190 3148 3194 3152
rect 3158 3138 3162 3142
rect 3262 3138 3266 3142
rect 3278 3138 3282 3142
rect 3038 3108 3042 3112
rect 3046 3088 3050 3092
rect 2990 3078 2994 3082
rect 3054 3078 3058 3082
rect 2974 3058 2978 3062
rect 2982 3058 2986 3062
rect 3006 3068 3010 3072
rect 3022 3068 3026 3072
rect 2998 3058 3002 3062
rect 3030 3048 3034 3052
rect 2974 3038 2978 3042
rect 3126 3078 3130 3082
rect 3142 3078 3146 3082
rect 3022 3028 3026 3032
rect 3070 3028 3074 3032
rect 2982 3018 2986 3022
rect 3054 3008 3058 3012
rect 2958 2988 2962 2992
rect 2694 2968 2698 2972
rect 2726 2968 2730 2972
rect 2894 2968 2898 2972
rect 2686 2958 2690 2962
rect 2686 2948 2690 2952
rect 2702 2948 2706 2952
rect 2718 2948 2722 2952
rect 2734 2958 2738 2962
rect 2742 2948 2746 2952
rect 2806 2948 2810 2952
rect 2870 2948 2874 2952
rect 2782 2938 2786 2942
rect 2798 2938 2802 2942
rect 2654 2928 2658 2932
rect 2670 2928 2674 2932
rect 2766 2928 2770 2932
rect 2798 2928 2802 2932
rect 2886 2938 2890 2942
rect 2878 2928 2882 2932
rect 2886 2928 2890 2932
rect 2646 2918 2650 2922
rect 2702 2918 2706 2922
rect 2822 2918 2826 2922
rect 2838 2918 2842 2922
rect 2846 2918 2850 2922
rect 2638 2878 2642 2882
rect 2558 2868 2562 2872
rect 2630 2868 2634 2872
rect 2646 2868 2650 2872
rect 2598 2858 2602 2862
rect 2478 2778 2482 2782
rect 2430 2768 2434 2772
rect 2462 2747 2466 2751
rect 2254 2678 2258 2682
rect 2278 2678 2282 2682
rect 2334 2678 2338 2682
rect 2278 2668 2282 2672
rect 2286 2668 2290 2672
rect 2262 2658 2266 2662
rect 2326 2668 2330 2672
rect 2310 2658 2314 2662
rect 2406 2678 2410 2682
rect 2422 2678 2426 2682
rect 2374 2668 2378 2672
rect 2382 2658 2386 2662
rect 2294 2648 2298 2652
rect 2302 2648 2306 2652
rect 2350 2648 2354 2652
rect 2366 2648 2370 2652
rect 2414 2648 2418 2652
rect 2054 2628 2058 2632
rect 2110 2628 2114 2632
rect 2246 2628 2250 2632
rect 2334 2628 2338 2632
rect 1974 2618 1978 2622
rect 1998 2618 2002 2622
rect 2014 2618 2018 2622
rect 1950 2598 1954 2602
rect 1798 2578 1802 2582
rect 1950 2578 1954 2582
rect 1966 2578 1970 2582
rect 1814 2568 1818 2572
rect 1830 2548 1834 2552
rect 1822 2498 1826 2502
rect 1806 2468 1810 2472
rect 1798 2458 1802 2462
rect 1790 2448 1794 2452
rect 1798 2438 1802 2442
rect 1822 2438 1826 2442
rect 1814 2388 1818 2392
rect 1806 2368 1810 2372
rect 1774 2338 1778 2342
rect 1806 2338 1810 2342
rect 1798 2318 1802 2322
rect 1790 2258 1794 2262
rect 1702 2248 1706 2252
rect 1766 2248 1770 2252
rect 1718 2238 1722 2242
rect 1766 2238 1770 2242
rect 1654 2178 1658 2182
rect 1806 2178 1810 2182
rect 1654 2168 1658 2172
rect 1702 2168 1706 2172
rect 1654 2158 1658 2162
rect 1646 2148 1650 2152
rect 1638 2138 1642 2142
rect 1654 2138 1658 2142
rect 1742 2158 1746 2162
rect 1678 2148 1682 2152
rect 1662 2118 1666 2122
rect 1646 2108 1650 2112
rect 1598 1958 1602 1962
rect 1630 1958 1634 1962
rect 1446 1948 1450 1952
rect 1494 1948 1498 1952
rect 1510 1948 1514 1952
rect 1550 1948 1554 1952
rect 1590 1948 1594 1952
rect 1350 1938 1354 1942
rect 1502 1938 1506 1942
rect 1390 1928 1394 1932
rect 1326 1918 1330 1922
rect 1294 1898 1298 1902
rect 1270 1888 1274 1892
rect 1318 1878 1322 1882
rect 990 1868 994 1872
rect 1054 1868 1058 1872
rect 1254 1868 1258 1872
rect 942 1858 946 1862
rect 958 1858 962 1862
rect 1022 1858 1026 1862
rect 1038 1858 1042 1862
rect 1086 1858 1090 1862
rect 1142 1858 1146 1862
rect 950 1848 954 1852
rect 974 1848 978 1852
rect 1022 1848 1026 1852
rect 1038 1848 1042 1852
rect 998 1838 1002 1842
rect 1006 1818 1010 1822
rect 918 1788 922 1792
rect 1350 1868 1354 1872
rect 1310 1858 1314 1862
rect 1302 1848 1306 1852
rect 1270 1838 1274 1842
rect 1318 1798 1322 1802
rect 918 1778 922 1782
rect 998 1778 1002 1782
rect 1078 1778 1082 1782
rect 1150 1778 1154 1782
rect 902 1758 906 1762
rect 742 1748 746 1752
rect 766 1748 770 1752
rect 774 1748 778 1752
rect 798 1748 802 1752
rect 494 1738 498 1742
rect 686 1738 690 1742
rect 782 1738 786 1742
rect 830 1738 834 1742
rect 454 1728 458 1732
rect 486 1728 490 1732
rect 366 1708 370 1712
rect 318 1678 322 1682
rect 326 1666 330 1670
rect 342 1668 346 1672
rect 366 1668 370 1672
rect 286 1658 290 1662
rect 310 1658 314 1662
rect 366 1658 370 1662
rect 398 1658 402 1662
rect 262 1648 266 1652
rect 246 1608 250 1612
rect 278 1638 282 1642
rect 294 1638 298 1642
rect 398 1638 402 1642
rect 542 1708 546 1712
rect 614 1728 618 1732
rect 670 1728 674 1732
rect 694 1728 698 1732
rect 558 1698 562 1702
rect 694 1698 698 1702
rect 694 1688 698 1692
rect 718 1688 722 1692
rect 766 1728 770 1732
rect 858 1703 862 1707
rect 865 1703 869 1707
rect 758 1698 762 1702
rect 822 1698 826 1702
rect 486 1678 490 1682
rect 622 1678 626 1682
rect 686 1678 690 1682
rect 710 1678 714 1682
rect 750 1678 754 1682
rect 542 1668 546 1672
rect 902 1748 906 1752
rect 926 1768 930 1772
rect 1038 1768 1042 1772
rect 1142 1768 1146 1772
rect 1230 1768 1234 1772
rect 1006 1758 1010 1762
rect 950 1748 954 1752
rect 942 1738 946 1742
rect 814 1688 818 1692
rect 822 1688 826 1692
rect 886 1688 890 1692
rect 942 1688 946 1692
rect 974 1738 978 1742
rect 990 1728 994 1732
rect 1086 1758 1090 1762
rect 1182 1758 1186 1762
rect 1214 1758 1218 1762
rect 1022 1738 1026 1742
rect 1102 1738 1106 1742
rect 1014 1718 1018 1722
rect 1070 1728 1074 1732
rect 1142 1728 1146 1732
rect 1134 1718 1138 1722
rect 1046 1708 1050 1712
rect 790 1678 794 1682
rect 846 1678 850 1682
rect 862 1678 866 1682
rect 886 1678 890 1682
rect 934 1678 938 1682
rect 966 1678 970 1682
rect 670 1668 674 1672
rect 694 1668 698 1672
rect 718 1668 722 1672
rect 758 1668 762 1672
rect 422 1658 426 1662
rect 446 1658 450 1662
rect 478 1658 482 1662
rect 278 1618 282 1622
rect 254 1568 258 1572
rect 174 1558 178 1562
rect 190 1548 194 1552
rect 214 1548 218 1552
rect 230 1548 234 1552
rect 182 1538 186 1542
rect 206 1538 210 1542
rect 222 1538 226 1542
rect 254 1528 258 1532
rect 190 1498 194 1502
rect 182 1478 186 1482
rect 134 1358 138 1362
rect 142 1328 146 1332
rect 62 1268 66 1272
rect 94 1268 98 1272
rect 126 1268 130 1272
rect 30 1258 34 1262
rect 78 1258 82 1262
rect 38 1248 42 1252
rect 54 1248 58 1252
rect 14 1208 18 1212
rect 198 1488 202 1492
rect 222 1488 226 1492
rect 206 1478 210 1482
rect 206 1468 210 1472
rect 214 1458 218 1462
rect 230 1448 234 1452
rect 326 1608 330 1612
rect 346 1603 350 1607
rect 353 1603 357 1607
rect 294 1558 298 1562
rect 318 1558 322 1562
rect 286 1548 290 1552
rect 382 1568 386 1572
rect 390 1568 394 1572
rect 358 1558 362 1562
rect 334 1548 338 1552
rect 302 1538 306 1542
rect 342 1538 346 1542
rect 318 1528 322 1532
rect 278 1488 282 1492
rect 374 1548 378 1552
rect 510 1628 514 1632
rect 542 1628 546 1632
rect 414 1568 418 1572
rect 614 1658 618 1662
rect 638 1658 642 1662
rect 686 1658 690 1662
rect 782 1658 786 1662
rect 566 1648 570 1652
rect 574 1638 578 1642
rect 630 1638 634 1642
rect 630 1628 634 1632
rect 782 1648 786 1652
rect 742 1638 746 1642
rect 646 1608 650 1612
rect 638 1578 642 1582
rect 710 1578 714 1582
rect 558 1558 562 1562
rect 590 1558 594 1562
rect 430 1548 434 1552
rect 398 1528 402 1532
rect 478 1528 482 1532
rect 534 1528 538 1532
rect 510 1518 514 1522
rect 654 1568 658 1572
rect 678 1568 682 1572
rect 662 1548 666 1552
rect 614 1538 618 1542
rect 654 1538 658 1542
rect 894 1668 898 1672
rect 846 1658 850 1662
rect 798 1628 802 1632
rect 902 1658 906 1662
rect 918 1658 922 1662
rect 846 1648 850 1652
rect 886 1648 890 1652
rect 902 1648 906 1652
rect 806 1618 810 1622
rect 886 1628 890 1632
rect 830 1608 834 1612
rect 814 1598 818 1602
rect 822 1578 826 1582
rect 790 1568 794 1572
rect 814 1568 818 1572
rect 718 1548 722 1552
rect 742 1548 746 1552
rect 766 1548 770 1552
rect 726 1538 730 1542
rect 734 1538 738 1542
rect 598 1528 602 1532
rect 670 1528 674 1532
rect 678 1528 682 1532
rect 718 1528 722 1532
rect 462 1508 466 1512
rect 606 1518 610 1522
rect 470 1488 474 1492
rect 550 1488 554 1492
rect 254 1478 258 1482
rect 422 1478 426 1482
rect 486 1478 490 1482
rect 702 1518 706 1522
rect 686 1508 690 1512
rect 622 1498 626 1502
rect 310 1468 314 1472
rect 326 1458 330 1462
rect 422 1448 426 1452
rect 374 1438 378 1442
rect 222 1418 226 1422
rect 214 1348 218 1352
rect 346 1403 350 1407
rect 353 1403 357 1407
rect 454 1448 458 1452
rect 278 1378 282 1382
rect 430 1378 434 1382
rect 446 1378 450 1382
rect 254 1348 258 1352
rect 302 1368 306 1372
rect 310 1368 314 1372
rect 286 1358 290 1362
rect 366 1358 370 1362
rect 382 1358 386 1362
rect 358 1348 362 1352
rect 430 1358 434 1362
rect 438 1358 442 1362
rect 470 1358 474 1362
rect 494 1358 498 1362
rect 406 1348 410 1352
rect 310 1338 314 1342
rect 366 1338 370 1342
rect 390 1338 394 1342
rect 198 1328 202 1332
rect 214 1318 218 1322
rect 230 1328 234 1332
rect 270 1328 274 1332
rect 318 1328 322 1332
rect 382 1328 386 1332
rect 390 1328 394 1332
rect 222 1308 226 1312
rect 238 1288 242 1292
rect 286 1278 290 1282
rect 246 1268 250 1272
rect 222 1258 226 1262
rect 238 1248 242 1252
rect 262 1248 266 1252
rect 270 1248 274 1252
rect 286 1248 290 1252
rect 158 1238 162 1242
rect 158 1228 162 1232
rect 238 1228 242 1232
rect 46 1208 50 1212
rect 110 1208 114 1212
rect 22 1198 26 1202
rect 38 1198 42 1202
rect 214 1198 218 1202
rect 126 1188 130 1192
rect 158 1168 162 1172
rect 174 1168 178 1172
rect 214 1168 218 1172
rect 94 1148 98 1152
rect 110 1148 114 1152
rect 166 1158 170 1162
rect 134 1148 138 1152
rect 150 1148 154 1152
rect 174 1148 178 1152
rect 126 1138 130 1142
rect 54 1098 58 1102
rect 38 1068 42 1072
rect 190 1138 194 1142
rect 94 1128 98 1132
rect 126 1118 130 1122
rect 78 1078 82 1082
rect 86 1078 90 1082
rect 182 1108 186 1112
rect 262 1238 266 1242
rect 254 1218 258 1222
rect 286 1178 290 1182
rect 230 1148 234 1152
rect 310 1308 314 1312
rect 350 1278 354 1282
rect 310 1208 314 1212
rect 326 1258 330 1262
rect 462 1338 466 1342
rect 486 1338 490 1342
rect 486 1328 490 1332
rect 454 1318 458 1322
rect 446 1298 450 1302
rect 494 1298 498 1302
rect 814 1558 818 1562
rect 878 1598 882 1602
rect 838 1558 842 1562
rect 894 1618 898 1622
rect 958 1658 962 1662
rect 1166 1708 1170 1712
rect 1214 1708 1218 1712
rect 1142 1698 1146 1702
rect 1158 1688 1162 1692
rect 974 1668 978 1672
rect 974 1658 978 1662
rect 942 1648 946 1652
rect 974 1648 978 1652
rect 1054 1658 1058 1662
rect 1070 1658 1074 1662
rect 1094 1658 1098 1662
rect 1110 1658 1114 1662
rect 1142 1668 1146 1672
rect 1182 1688 1186 1692
rect 1206 1688 1210 1692
rect 1222 1698 1226 1702
rect 1174 1658 1178 1662
rect 1078 1648 1082 1652
rect 1134 1648 1138 1652
rect 1182 1648 1186 1652
rect 1038 1638 1042 1642
rect 1062 1638 1066 1642
rect 1078 1638 1082 1642
rect 1126 1638 1130 1642
rect 918 1608 922 1612
rect 966 1608 970 1612
rect 902 1598 906 1602
rect 950 1598 954 1602
rect 998 1598 1002 1602
rect 1102 1628 1106 1632
rect 1110 1628 1114 1632
rect 1038 1578 1042 1582
rect 966 1568 970 1572
rect 974 1568 978 1572
rect 1014 1568 1018 1572
rect 1054 1568 1058 1572
rect 1070 1568 1074 1572
rect 1142 1568 1146 1572
rect 902 1558 906 1562
rect 910 1558 914 1562
rect 998 1558 1002 1562
rect 806 1548 810 1552
rect 830 1548 834 1552
rect 870 1548 874 1552
rect 894 1548 898 1552
rect 918 1548 922 1552
rect 926 1548 930 1552
rect 942 1548 946 1552
rect 1006 1548 1010 1552
rect 846 1538 850 1542
rect 934 1538 938 1542
rect 950 1538 954 1542
rect 1022 1538 1026 1542
rect 1046 1538 1050 1542
rect 1206 1558 1210 1562
rect 1302 1738 1306 1742
rect 1430 1908 1434 1912
rect 1382 1898 1386 1902
rect 1526 1938 1530 1942
rect 1542 1938 1546 1942
rect 1534 1928 1538 1932
rect 1446 1918 1450 1922
rect 1574 1918 1578 1922
rect 1446 1908 1450 1912
rect 1438 1878 1442 1882
rect 1370 1803 1374 1807
rect 1377 1803 1381 1807
rect 1430 1758 1434 1762
rect 1422 1748 1426 1752
rect 1382 1738 1386 1742
rect 1398 1718 1402 1722
rect 1326 1658 1330 1662
rect 1270 1648 1274 1652
rect 1286 1648 1290 1652
rect 1318 1648 1322 1652
rect 1334 1638 1338 1642
rect 1398 1618 1402 1622
rect 1370 1603 1374 1607
rect 1377 1603 1381 1607
rect 1334 1588 1338 1592
rect 1078 1548 1082 1552
rect 1126 1548 1130 1552
rect 1166 1548 1170 1552
rect 1318 1548 1322 1552
rect 1086 1538 1090 1542
rect 1118 1538 1122 1542
rect 1134 1538 1138 1542
rect 1150 1538 1154 1542
rect 1174 1538 1178 1542
rect 1310 1538 1314 1542
rect 758 1528 762 1532
rect 782 1528 786 1532
rect 790 1528 794 1532
rect 1030 1528 1034 1532
rect 1054 1528 1058 1532
rect 1126 1528 1130 1532
rect 1142 1528 1146 1532
rect 742 1498 746 1502
rect 726 1488 730 1492
rect 766 1488 770 1492
rect 686 1478 690 1482
rect 646 1468 650 1472
rect 638 1458 642 1462
rect 646 1448 650 1452
rect 858 1503 862 1507
rect 865 1503 869 1507
rect 902 1488 906 1492
rect 1118 1488 1122 1492
rect 742 1478 746 1482
rect 774 1478 778 1482
rect 694 1468 698 1472
rect 734 1468 738 1472
rect 758 1468 762 1472
rect 862 1468 866 1472
rect 878 1458 882 1462
rect 662 1438 666 1442
rect 558 1428 562 1432
rect 558 1418 562 1422
rect 694 1448 698 1452
rect 990 1458 994 1462
rect 1030 1458 1034 1462
rect 1110 1458 1114 1462
rect 1094 1448 1098 1452
rect 974 1438 978 1442
rect 790 1418 794 1422
rect 1022 1418 1026 1422
rect 742 1408 746 1412
rect 686 1398 690 1402
rect 606 1358 610 1362
rect 630 1358 634 1362
rect 670 1358 674 1362
rect 518 1348 522 1352
rect 550 1348 554 1352
rect 582 1348 586 1352
rect 614 1348 618 1352
rect 662 1348 666 1352
rect 1158 1468 1162 1472
rect 1134 1398 1138 1402
rect 1254 1528 1258 1532
rect 1222 1478 1226 1482
rect 1294 1478 1298 1482
rect 1190 1468 1194 1472
rect 1246 1468 1250 1472
rect 1182 1438 1186 1442
rect 1230 1448 1234 1452
rect 1238 1448 1242 1452
rect 1254 1448 1258 1452
rect 1302 1468 1306 1472
rect 1310 1468 1314 1472
rect 1294 1458 1298 1462
rect 1310 1448 1314 1452
rect 1278 1438 1282 1442
rect 1310 1428 1314 1432
rect 1174 1388 1178 1392
rect 1110 1378 1114 1382
rect 958 1368 962 1372
rect 966 1368 970 1372
rect 814 1358 818 1362
rect 822 1358 826 1362
rect 750 1348 754 1352
rect 518 1338 522 1342
rect 558 1338 562 1342
rect 510 1318 514 1322
rect 430 1288 434 1292
rect 502 1288 506 1292
rect 422 1278 426 1282
rect 414 1268 418 1272
rect 454 1278 458 1282
rect 502 1278 506 1282
rect 558 1328 562 1332
rect 622 1328 626 1332
rect 526 1298 530 1302
rect 550 1298 554 1302
rect 582 1298 586 1302
rect 566 1288 570 1292
rect 590 1278 594 1282
rect 486 1268 490 1272
rect 678 1318 682 1322
rect 694 1318 698 1322
rect 702 1318 706 1322
rect 814 1318 818 1322
rect 614 1268 618 1272
rect 414 1258 418 1262
rect 454 1258 458 1262
rect 358 1248 362 1252
rect 398 1238 402 1242
rect 334 1228 338 1232
rect 406 1228 410 1232
rect 326 1198 330 1202
rect 346 1203 350 1207
rect 353 1203 357 1207
rect 318 1188 322 1192
rect 486 1238 490 1242
rect 486 1228 490 1232
rect 462 1188 466 1192
rect 318 1178 322 1182
rect 438 1178 442 1182
rect 406 1158 410 1162
rect 414 1158 418 1162
rect 438 1158 442 1162
rect 254 1138 258 1142
rect 286 1138 290 1142
rect 302 1138 306 1142
rect 230 1128 234 1132
rect 270 1128 274 1132
rect 462 1148 466 1152
rect 534 1168 538 1172
rect 510 1158 514 1162
rect 494 1148 498 1152
rect 414 1138 418 1142
rect 606 1238 610 1242
rect 614 1228 618 1232
rect 766 1308 770 1312
rect 1134 1368 1138 1372
rect 838 1318 842 1322
rect 858 1303 862 1307
rect 865 1303 869 1307
rect 758 1288 762 1292
rect 822 1288 826 1292
rect 854 1288 858 1292
rect 862 1288 866 1292
rect 838 1278 842 1282
rect 846 1278 850 1282
rect 726 1268 730 1272
rect 766 1268 770 1272
rect 734 1258 738 1262
rect 710 1248 714 1252
rect 742 1248 746 1252
rect 830 1268 834 1272
rect 782 1258 786 1262
rect 774 1248 778 1252
rect 806 1258 810 1262
rect 830 1258 834 1262
rect 710 1238 714 1242
rect 750 1238 754 1242
rect 670 1208 674 1212
rect 710 1208 714 1212
rect 622 1188 626 1192
rect 726 1188 730 1192
rect 622 1178 626 1182
rect 742 1168 746 1172
rect 766 1168 770 1172
rect 558 1158 562 1162
rect 558 1148 562 1152
rect 598 1148 602 1152
rect 678 1148 682 1152
rect 718 1148 722 1152
rect 742 1148 746 1152
rect 774 1148 778 1152
rect 574 1138 578 1142
rect 582 1138 586 1142
rect 646 1138 650 1142
rect 694 1138 698 1142
rect 358 1128 362 1132
rect 422 1128 426 1132
rect 542 1128 546 1132
rect 566 1128 570 1132
rect 526 1118 530 1122
rect 558 1118 562 1122
rect 574 1118 578 1122
rect 262 1108 266 1112
rect 310 1108 314 1112
rect 326 1108 330 1112
rect 518 1098 522 1102
rect 230 1088 234 1092
rect 278 1088 282 1092
rect 374 1088 378 1092
rect 470 1088 474 1092
rect 150 1078 154 1082
rect 174 1078 178 1082
rect 214 1078 218 1082
rect 270 1078 274 1082
rect 62 1068 66 1072
rect 70 1068 74 1072
rect 550 1108 554 1112
rect 374 1078 378 1082
rect 406 1078 410 1082
rect 478 1078 482 1082
rect 174 1068 178 1072
rect 278 1068 282 1072
rect 78 1058 82 1062
rect 126 1058 130 1062
rect 142 1058 146 1062
rect 62 1048 66 1052
rect 150 1048 154 1052
rect 190 1048 194 1052
rect 30 1038 34 1042
rect 102 1038 106 1042
rect 126 988 130 992
rect 78 968 82 972
rect 110 888 114 892
rect 62 868 66 872
rect 166 978 170 982
rect 198 978 202 982
rect 142 958 146 962
rect 182 958 186 962
rect 198 958 202 962
rect 158 948 162 952
rect 198 938 202 942
rect 286 1058 290 1062
rect 294 1058 298 1062
rect 246 1038 250 1042
rect 346 1003 350 1007
rect 353 1003 357 1007
rect 302 978 306 982
rect 246 968 250 972
rect 222 948 226 952
rect 278 938 282 942
rect 222 928 226 932
rect 390 1058 394 1062
rect 430 1058 434 1062
rect 470 1058 474 1062
rect 382 998 386 1002
rect 502 1048 506 1052
rect 446 1038 450 1042
rect 454 1038 458 1042
rect 438 1008 442 1012
rect 414 968 418 972
rect 398 958 402 962
rect 438 958 442 962
rect 414 948 418 952
rect 286 928 290 932
rect 270 918 274 922
rect 206 888 210 892
rect 214 888 218 892
rect 262 878 266 882
rect 334 878 338 882
rect 158 868 162 872
rect 126 859 130 862
rect 126 858 130 859
rect 390 938 394 942
rect 398 928 402 932
rect 390 918 394 922
rect 390 868 394 872
rect 278 858 282 862
rect 294 858 298 862
rect 478 978 482 982
rect 470 968 474 972
rect 454 938 458 942
rect 422 928 426 932
rect 446 918 450 922
rect 406 878 410 882
rect 446 898 450 902
rect 510 1028 514 1032
rect 534 1048 538 1052
rect 542 1048 546 1052
rect 566 1068 570 1072
rect 558 1048 562 1052
rect 542 1038 546 1042
rect 534 1018 538 1022
rect 518 998 522 1002
rect 510 968 514 972
rect 518 968 522 972
rect 510 948 514 952
rect 486 908 490 912
rect 502 908 506 912
rect 470 898 474 902
rect 446 878 450 882
rect 590 1068 594 1072
rect 582 1058 586 1062
rect 702 1128 706 1132
rect 742 1128 746 1132
rect 662 1108 666 1112
rect 678 1108 682 1112
rect 630 1078 634 1082
rect 606 1068 610 1072
rect 646 1068 650 1072
rect 630 1058 634 1062
rect 758 1118 762 1122
rect 702 1078 706 1082
rect 734 1078 738 1082
rect 814 1188 818 1192
rect 806 1168 810 1172
rect 822 1168 826 1172
rect 918 1358 922 1362
rect 1006 1358 1010 1362
rect 894 1338 898 1342
rect 934 1338 938 1342
rect 974 1338 978 1342
rect 902 1328 906 1332
rect 958 1328 962 1332
rect 886 1308 890 1312
rect 886 1288 890 1292
rect 894 1278 898 1282
rect 902 1268 906 1272
rect 926 1208 930 1212
rect 902 1188 906 1192
rect 790 1158 794 1162
rect 822 1158 826 1162
rect 806 1148 810 1152
rect 830 1148 834 1152
rect 942 1298 946 1302
rect 1014 1348 1018 1352
rect 1038 1358 1042 1362
rect 1062 1358 1066 1362
rect 1086 1358 1090 1362
rect 1142 1358 1146 1362
rect 1046 1348 1050 1352
rect 1070 1348 1074 1352
rect 1134 1348 1138 1352
rect 1174 1348 1178 1352
rect 1022 1338 1026 1342
rect 1054 1338 1058 1342
rect 1078 1338 1082 1342
rect 1086 1338 1090 1342
rect 1126 1338 1130 1342
rect 1142 1338 1146 1342
rect 1182 1338 1186 1342
rect 998 1328 1002 1332
rect 1150 1328 1154 1332
rect 1262 1328 1266 1332
rect 990 1318 994 1322
rect 942 1278 946 1282
rect 958 1278 962 1282
rect 966 1278 970 1282
rect 990 1278 994 1282
rect 1014 1318 1018 1322
rect 1182 1318 1186 1322
rect 1030 1298 1034 1302
rect 1086 1288 1090 1292
rect 1022 1278 1026 1282
rect 1126 1278 1130 1282
rect 1182 1278 1186 1282
rect 1054 1268 1058 1272
rect 1062 1268 1066 1272
rect 1094 1268 1098 1272
rect 1118 1268 1122 1272
rect 998 1258 1002 1262
rect 966 1208 970 1212
rect 1006 1248 1010 1252
rect 990 1198 994 1202
rect 1030 1198 1034 1202
rect 1134 1268 1138 1272
rect 1142 1248 1146 1252
rect 1262 1318 1266 1322
rect 1206 1288 1210 1292
rect 1254 1288 1258 1292
rect 1214 1278 1218 1282
rect 1230 1278 1234 1282
rect 1198 1268 1202 1272
rect 1206 1248 1210 1252
rect 1222 1268 1226 1272
rect 1550 1888 1554 1892
rect 1598 1908 1602 1912
rect 1606 1898 1610 1902
rect 1654 2098 1658 2102
rect 1710 2148 1714 2152
rect 1726 2148 1730 2152
rect 1702 2138 1706 2142
rect 1718 2138 1722 2142
rect 1694 2118 1698 2122
rect 1886 2538 1890 2542
rect 1874 2503 1878 2507
rect 1881 2503 1885 2507
rect 2206 2608 2210 2612
rect 2142 2598 2146 2602
rect 2270 2588 2274 2592
rect 2206 2558 2210 2562
rect 2038 2548 2042 2552
rect 2022 2538 2026 2542
rect 2078 2538 2082 2542
rect 2310 2547 2314 2551
rect 2214 2538 2218 2542
rect 2238 2538 2242 2542
rect 2254 2528 2258 2532
rect 2382 2638 2386 2642
rect 2246 2518 2250 2522
rect 2262 2518 2266 2522
rect 2358 2518 2362 2522
rect 2246 2508 2250 2512
rect 2134 2498 2138 2502
rect 2158 2498 2162 2502
rect 1998 2478 2002 2482
rect 2102 2478 2106 2482
rect 2158 2478 2162 2482
rect 1854 2468 1858 2472
rect 1878 2459 1882 2463
rect 1926 2418 1930 2422
rect 1918 2398 1922 2402
rect 1926 2398 1930 2402
rect 1830 2378 1834 2382
rect 1846 2368 1850 2372
rect 1886 2368 1890 2372
rect 1918 2368 1922 2372
rect 1822 2348 1826 2352
rect 1838 2348 1842 2352
rect 1854 2348 1858 2352
rect 1894 2348 1898 2352
rect 1910 2348 1914 2352
rect 2014 2468 2018 2472
rect 2038 2468 2042 2472
rect 1966 2398 1970 2402
rect 1942 2378 1946 2382
rect 1982 2398 1986 2402
rect 2022 2458 2026 2462
rect 2150 2468 2154 2472
rect 2006 2448 2010 2452
rect 2070 2448 2074 2452
rect 2006 2418 2010 2422
rect 1990 2378 1994 2382
rect 2006 2378 2010 2382
rect 2078 2368 2082 2372
rect 1942 2358 1946 2362
rect 1950 2358 1954 2362
rect 1974 2358 1978 2362
rect 1998 2358 2002 2362
rect 2022 2358 2026 2362
rect 1934 2348 1938 2352
rect 1862 2328 1866 2332
rect 1878 2328 1882 2332
rect 1894 2328 1898 2332
rect 1902 2328 1906 2332
rect 1874 2303 1878 2307
rect 1881 2303 1885 2307
rect 1854 2288 1858 2292
rect 1878 2288 1882 2292
rect 1830 2278 1834 2282
rect 1870 2268 1874 2272
rect 1878 2268 1882 2272
rect 1838 2218 1842 2222
rect 1830 2188 1834 2192
rect 1878 2258 1882 2262
rect 1846 2188 1850 2192
rect 1902 2318 1906 2322
rect 1926 2318 1930 2322
rect 1942 2318 1946 2322
rect 1902 2308 1906 2312
rect 1934 2308 1938 2312
rect 1918 2238 1922 2242
rect 2006 2328 2010 2332
rect 1966 2308 1970 2312
rect 1950 2298 1954 2302
rect 1966 2298 1970 2302
rect 1958 2288 1962 2292
rect 1942 2258 1946 2262
rect 1950 2228 1954 2232
rect 2014 2308 2018 2312
rect 2030 2338 2034 2342
rect 2030 2318 2034 2322
rect 2062 2318 2066 2322
rect 2118 2448 2122 2452
rect 2094 2278 2098 2282
rect 2110 2278 2114 2282
rect 2062 2268 2066 2272
rect 2102 2268 2106 2272
rect 1990 2258 1994 2262
rect 2070 2258 2074 2262
rect 2102 2258 2106 2262
rect 2198 2448 2202 2452
rect 2222 2448 2226 2452
rect 2190 2438 2194 2442
rect 2166 2418 2170 2422
rect 2158 2408 2162 2412
rect 2126 2398 2130 2402
rect 2254 2498 2258 2502
rect 2286 2478 2290 2482
rect 2126 2378 2130 2382
rect 2222 2348 2226 2352
rect 2190 2338 2194 2342
rect 2214 2338 2218 2342
rect 2182 2328 2186 2332
rect 2214 2328 2218 2332
rect 2254 2318 2258 2322
rect 2238 2308 2242 2312
rect 2198 2288 2202 2292
rect 2022 2248 2026 2252
rect 2054 2248 2058 2252
rect 1974 2228 1978 2232
rect 2078 2208 2082 2212
rect 1990 2198 1994 2202
rect 2070 2198 2074 2202
rect 1934 2168 1938 2172
rect 1958 2168 1962 2172
rect 1654 2048 1658 2052
rect 1758 2118 1762 2122
rect 1894 2138 1898 2142
rect 1942 2138 1946 2142
rect 1878 2128 1882 2132
rect 1874 2103 1878 2107
rect 1881 2103 1885 2107
rect 1814 2098 1818 2102
rect 1774 2078 1778 2082
rect 1782 2078 1786 2082
rect 1758 2068 1762 2072
rect 1846 2068 1850 2072
rect 1910 2088 1914 2092
rect 1926 2088 1930 2092
rect 2102 2178 2106 2182
rect 2014 2147 2018 2151
rect 2006 2138 2010 2142
rect 2086 2138 2090 2142
rect 2062 2118 2066 2122
rect 1998 2108 2002 2112
rect 2094 2108 2098 2112
rect 2246 2278 2250 2282
rect 2134 2248 2138 2252
rect 2150 2248 2154 2252
rect 2126 2208 2130 2212
rect 2190 2258 2194 2262
rect 2222 2258 2226 2262
rect 2246 2258 2250 2262
rect 2174 2248 2178 2252
rect 2222 2248 2226 2252
rect 2182 2238 2186 2242
rect 2222 2218 2226 2222
rect 2174 2208 2178 2212
rect 2190 2208 2194 2212
rect 2150 2198 2154 2202
rect 2158 2198 2162 2202
rect 2118 2168 2122 2172
rect 2142 2168 2146 2172
rect 2182 2158 2186 2162
rect 2150 2148 2154 2152
rect 2118 2138 2122 2142
rect 2142 2138 2146 2142
rect 2158 2128 2162 2132
rect 2206 2138 2210 2142
rect 2302 2448 2306 2452
rect 2318 2448 2322 2452
rect 2350 2448 2354 2452
rect 2342 2398 2346 2402
rect 2394 2603 2398 2607
rect 2401 2603 2405 2607
rect 2454 2648 2458 2652
rect 2422 2628 2426 2632
rect 2438 2628 2442 2632
rect 2518 2808 2522 2812
rect 2518 2768 2522 2772
rect 2510 2748 2514 2752
rect 2550 2738 2554 2742
rect 2526 2678 2530 2682
rect 2630 2848 2634 2852
rect 2686 2868 2690 2872
rect 2742 2868 2746 2872
rect 2774 2868 2778 2872
rect 2790 2868 2794 2872
rect 2662 2858 2666 2862
rect 2678 2848 2682 2852
rect 2686 2848 2690 2852
rect 2734 2858 2738 2862
rect 2686 2828 2690 2832
rect 2622 2818 2626 2822
rect 2654 2818 2658 2822
rect 3038 2958 3042 2962
rect 2942 2948 2946 2952
rect 2958 2948 2962 2952
rect 3046 2948 3050 2952
rect 2894 2908 2898 2912
rect 2906 2903 2910 2907
rect 2913 2903 2917 2907
rect 2942 2888 2946 2892
rect 2998 2888 3002 2892
rect 3006 2878 3010 2882
rect 2862 2868 2866 2872
rect 2918 2868 2922 2872
rect 2814 2858 2818 2862
rect 2774 2848 2778 2852
rect 2758 2838 2762 2842
rect 2798 2838 2802 2842
rect 2806 2838 2810 2842
rect 2830 2838 2834 2842
rect 2846 2838 2850 2842
rect 2862 2838 2866 2842
rect 2894 2858 2898 2862
rect 2926 2858 2930 2862
rect 2982 2858 2986 2862
rect 2878 2848 2882 2852
rect 2918 2848 2922 2852
rect 2942 2848 2946 2852
rect 2966 2848 2970 2852
rect 2990 2848 2994 2852
rect 2886 2838 2890 2842
rect 2870 2828 2874 2832
rect 2750 2818 2754 2822
rect 2702 2808 2706 2812
rect 2726 2808 2730 2812
rect 2614 2798 2618 2802
rect 2782 2798 2786 2802
rect 2630 2778 2634 2782
rect 2734 2758 2738 2762
rect 2630 2738 2634 2742
rect 2694 2738 2698 2742
rect 2702 2728 2706 2732
rect 2830 2768 2834 2772
rect 2854 2768 2858 2772
rect 2894 2828 2898 2832
rect 2950 2828 2954 2832
rect 2974 2828 2978 2832
rect 3038 2908 3042 2912
rect 3102 3058 3106 3062
rect 3134 3058 3138 3062
rect 3134 2998 3138 3002
rect 3126 2988 3130 2992
rect 3078 2978 3082 2982
rect 3070 2958 3074 2962
rect 3118 2958 3122 2962
rect 3134 2958 3138 2962
rect 3086 2948 3090 2952
rect 3070 2938 3074 2942
rect 3086 2928 3090 2932
rect 3262 3098 3266 3102
rect 3342 3208 3346 3212
rect 3294 3158 3298 3162
rect 3334 3148 3338 3152
rect 3358 3148 3362 3152
rect 3326 3138 3330 3142
rect 3430 3328 3434 3332
rect 3454 3328 3458 3332
rect 3422 3298 3426 3302
rect 3398 3268 3402 3272
rect 3406 3268 3410 3272
rect 3446 3318 3450 3322
rect 3510 3318 3514 3322
rect 3550 3288 3554 3292
rect 3462 3268 3466 3272
rect 3494 3268 3498 3272
rect 3510 3268 3514 3272
rect 3438 3258 3442 3262
rect 3430 3228 3434 3232
rect 3382 3218 3386 3222
rect 3382 3208 3386 3212
rect 3418 3203 3422 3207
rect 3425 3203 3429 3207
rect 3406 3168 3410 3172
rect 3462 3168 3466 3172
rect 3374 3128 3378 3132
rect 3238 3088 3242 3092
rect 3206 3058 3210 3062
rect 3222 3058 3226 3062
rect 3318 3108 3322 3112
rect 3310 3078 3314 3082
rect 3318 3078 3322 3082
rect 3262 3058 3266 3062
rect 3182 3048 3186 3052
rect 3222 3048 3226 3052
rect 3270 3048 3274 3052
rect 3238 3038 3242 3042
rect 3262 3038 3266 3042
rect 3206 2998 3210 3002
rect 3174 2958 3178 2962
rect 3142 2948 3146 2952
rect 3222 2948 3226 2952
rect 3150 2938 3154 2942
rect 3190 2938 3194 2942
rect 3142 2918 3146 2922
rect 3102 2898 3106 2902
rect 3134 2888 3138 2892
rect 3126 2878 3130 2882
rect 3022 2868 3026 2872
rect 3262 3028 3266 3032
rect 3254 2968 3258 2972
rect 3278 2978 3282 2982
rect 3326 3068 3330 3072
rect 3478 3238 3482 3242
rect 3502 3258 3506 3262
rect 3494 3238 3498 3242
rect 3486 3228 3490 3232
rect 3542 3248 3546 3252
rect 3654 3328 3658 3332
rect 3606 3298 3610 3302
rect 3566 3268 3570 3272
rect 3574 3268 3578 3272
rect 3654 3258 3658 3262
rect 3718 3308 3722 3312
rect 3742 3308 3746 3312
rect 3766 3308 3770 3312
rect 3902 3508 3906 3512
rect 3982 3558 3986 3562
rect 4070 3618 4074 3622
rect 4046 3588 4050 3592
rect 3926 3538 3930 3542
rect 3930 3503 3934 3507
rect 3937 3503 3941 3507
rect 3918 3478 3922 3482
rect 4062 3538 4066 3542
rect 4102 3578 4106 3582
rect 4094 3558 4098 3562
rect 4086 3538 4090 3542
rect 4182 3688 4186 3692
rect 4190 3678 4194 3682
rect 4174 3658 4178 3662
rect 4182 3648 4186 3652
rect 4134 3588 4138 3592
rect 4182 3578 4186 3582
rect 4174 3558 4178 3562
rect 4166 3548 4170 3552
rect 4126 3538 4130 3542
rect 4150 3538 4154 3542
rect 4190 3538 4194 3542
rect 4214 3698 4218 3702
rect 4238 3698 4242 3702
rect 4294 3698 4298 3702
rect 4342 3688 4346 3692
rect 4302 3668 4306 3672
rect 4238 3648 4242 3652
rect 4246 3638 4250 3642
rect 4374 3698 4378 3702
rect 4374 3688 4378 3692
rect 4326 3658 4330 3662
rect 4446 3678 4450 3682
rect 4662 3678 4666 3682
rect 4710 3678 4714 3682
rect 4726 3678 4730 3682
rect 4734 3678 4738 3682
rect 4846 3678 4850 3682
rect 4366 3658 4370 3662
rect 4358 3648 4362 3652
rect 4350 3638 4354 3642
rect 4398 3648 4402 3652
rect 4390 3638 4394 3642
rect 4422 3668 4426 3672
rect 4534 3668 4538 3672
rect 4558 3668 4562 3672
rect 4702 3668 4706 3672
rect 4430 3658 4434 3662
rect 4446 3658 4450 3662
rect 4510 3658 4514 3662
rect 4462 3638 4466 3642
rect 4414 3628 4418 3632
rect 4390 3588 4394 3592
rect 4374 3578 4378 3582
rect 4310 3568 4314 3572
rect 4334 3568 4338 3572
rect 4350 3568 4354 3572
rect 4374 3568 4378 3572
rect 4222 3558 4226 3562
rect 4310 3558 4314 3562
rect 4214 3548 4218 3552
rect 4326 3538 4330 3542
rect 4118 3508 4122 3512
rect 4062 3478 4066 3482
rect 3950 3468 3954 3472
rect 4038 3468 4042 3472
rect 4110 3468 4114 3472
rect 3862 3458 3866 3462
rect 3798 3428 3802 3432
rect 3846 3428 3850 3432
rect 3814 3358 3818 3362
rect 3950 3448 3954 3452
rect 3950 3388 3954 3392
rect 3886 3368 3890 3372
rect 3854 3358 3858 3362
rect 3854 3348 3858 3352
rect 3926 3348 3930 3352
rect 3798 3328 3802 3332
rect 3782 3318 3786 3322
rect 3838 3338 3842 3342
rect 3902 3338 3906 3342
rect 3894 3328 3898 3332
rect 3918 3328 3922 3332
rect 3822 3298 3826 3302
rect 3846 3298 3850 3302
rect 3702 3248 3706 3252
rect 3758 3248 3762 3252
rect 3614 3238 3618 3242
rect 3638 3238 3642 3242
rect 3710 3238 3714 3242
rect 3718 3238 3722 3242
rect 3558 3228 3562 3232
rect 3510 3168 3514 3172
rect 3534 3168 3538 3172
rect 3574 3168 3578 3172
rect 3430 3158 3434 3162
rect 3494 3158 3498 3162
rect 3566 3158 3570 3162
rect 3598 3158 3602 3162
rect 3694 3158 3698 3162
rect 3438 3148 3442 3152
rect 3454 3148 3458 3152
rect 3430 3138 3434 3142
rect 3438 3128 3442 3132
rect 3558 3148 3562 3152
rect 3486 3138 3490 3142
rect 3510 3138 3514 3142
rect 3382 3118 3386 3122
rect 3446 3118 3450 3122
rect 3366 3088 3370 3092
rect 3358 3078 3362 3082
rect 3350 3068 3354 3072
rect 3374 3068 3378 3072
rect 3342 3048 3346 3052
rect 3350 3048 3354 3052
rect 3366 3038 3370 3042
rect 3310 3028 3314 3032
rect 3294 2968 3298 2972
rect 3430 3078 3434 3082
rect 3446 3078 3450 3082
rect 3398 3068 3402 3072
rect 3406 3068 3410 3072
rect 3462 3068 3466 3072
rect 3398 3048 3402 3052
rect 3398 3038 3402 3042
rect 3438 3038 3442 3042
rect 3454 3038 3458 3042
rect 3462 3038 3466 3042
rect 3390 3028 3394 3032
rect 3382 2988 3386 2992
rect 3326 2978 3330 2982
rect 3374 2978 3378 2982
rect 3310 2968 3314 2972
rect 3342 2968 3346 2972
rect 3350 2968 3354 2972
rect 3382 2958 3386 2962
rect 3302 2948 3306 2952
rect 3326 2948 3330 2952
rect 3358 2948 3362 2952
rect 3262 2938 3266 2942
rect 3318 2938 3322 2942
rect 3334 2938 3338 2942
rect 3230 2928 3234 2932
rect 3182 2908 3186 2912
rect 3214 2908 3218 2912
rect 3150 2888 3154 2892
rect 3078 2858 3082 2862
rect 3110 2858 3114 2862
rect 3142 2858 3146 2862
rect 3014 2848 3018 2852
rect 3046 2848 3050 2852
rect 3126 2848 3130 2852
rect 3086 2838 3090 2842
rect 2958 2778 2962 2782
rect 2910 2768 2914 2772
rect 2926 2768 2930 2772
rect 2990 2768 2994 2772
rect 2798 2758 2802 2762
rect 2822 2758 2826 2762
rect 2846 2758 2850 2762
rect 2870 2758 2874 2762
rect 2790 2748 2794 2752
rect 2806 2748 2810 2752
rect 2838 2748 2842 2752
rect 2862 2748 2866 2752
rect 2878 2748 2882 2752
rect 2830 2738 2834 2742
rect 2662 2718 2666 2722
rect 2638 2698 2642 2702
rect 2582 2678 2586 2682
rect 2630 2678 2634 2682
rect 2550 2658 2554 2662
rect 2518 2598 2522 2602
rect 2502 2578 2506 2582
rect 2486 2558 2490 2562
rect 2406 2538 2410 2542
rect 2414 2448 2418 2452
rect 2394 2403 2398 2407
rect 2401 2403 2405 2407
rect 2374 2368 2378 2372
rect 2366 2348 2370 2352
rect 2398 2348 2402 2352
rect 2278 2338 2282 2342
rect 2366 2328 2370 2332
rect 2494 2528 2498 2532
rect 2494 2498 2498 2502
rect 2558 2518 2562 2522
rect 2750 2688 2754 2692
rect 2694 2658 2698 2662
rect 2854 2728 2858 2732
rect 2806 2708 2810 2712
rect 2854 2708 2858 2712
rect 2790 2658 2794 2662
rect 2598 2628 2602 2632
rect 2742 2628 2746 2632
rect 2742 2618 2746 2622
rect 2790 2618 2794 2622
rect 2654 2608 2658 2612
rect 2662 2598 2666 2602
rect 2614 2568 2618 2572
rect 2726 2538 2730 2542
rect 2630 2508 2634 2512
rect 2582 2498 2586 2502
rect 2622 2498 2626 2502
rect 2518 2478 2522 2482
rect 2518 2448 2522 2452
rect 2622 2448 2626 2452
rect 2518 2438 2522 2442
rect 2526 2418 2530 2422
rect 2550 2418 2554 2422
rect 2478 2408 2482 2412
rect 2590 2388 2594 2392
rect 2614 2388 2618 2392
rect 2502 2348 2506 2352
rect 2430 2338 2434 2342
rect 2398 2328 2402 2332
rect 2374 2298 2378 2302
rect 2454 2288 2458 2292
rect 2374 2278 2378 2282
rect 2286 2268 2290 2272
rect 2350 2268 2354 2272
rect 2366 2268 2370 2272
rect 2462 2278 2466 2282
rect 2534 2308 2538 2312
rect 2494 2268 2498 2272
rect 2510 2268 2514 2272
rect 2302 2258 2306 2262
rect 2262 2248 2266 2252
rect 2406 2248 2410 2252
rect 2254 2238 2258 2242
rect 2518 2238 2522 2242
rect 2358 2228 2362 2232
rect 2270 2188 2274 2192
rect 2254 2178 2258 2182
rect 2502 2218 2506 2222
rect 2394 2203 2398 2207
rect 2401 2203 2405 2207
rect 2382 2198 2386 2202
rect 2478 2168 2482 2172
rect 2326 2158 2330 2162
rect 2358 2158 2362 2162
rect 2438 2158 2442 2162
rect 2454 2158 2458 2162
rect 2470 2158 2474 2162
rect 2270 2148 2274 2152
rect 2286 2148 2290 2152
rect 2302 2148 2306 2152
rect 2214 2128 2218 2132
rect 2262 2128 2266 2132
rect 2270 2128 2274 2132
rect 2174 2118 2178 2122
rect 2190 2098 2194 2102
rect 2006 2078 2010 2082
rect 2078 2078 2082 2082
rect 1926 2068 1930 2072
rect 1726 2048 1730 2052
rect 1750 2048 1754 2052
rect 1774 2048 1778 2052
rect 1798 2048 1802 2052
rect 1822 2048 1826 2052
rect 1686 2038 1690 2042
rect 1718 2028 1722 2032
rect 1734 2008 1738 2012
rect 1686 1978 1690 1982
rect 1718 1978 1722 1982
rect 1662 1958 1666 1962
rect 1702 1968 1706 1972
rect 1814 2038 1818 2042
rect 1862 2048 1866 2052
rect 1782 2028 1786 2032
rect 1790 2028 1794 2032
rect 1838 2028 1842 2032
rect 1742 1968 1746 1972
rect 1774 1968 1778 1972
rect 1806 2018 1810 2022
rect 1814 2008 1818 2012
rect 1846 2008 1850 2012
rect 1838 1978 1842 1982
rect 1734 1948 1738 1952
rect 1742 1948 1746 1952
rect 1774 1948 1778 1952
rect 1790 1948 1794 1952
rect 1742 1938 1746 1942
rect 1654 1928 1658 1932
rect 1702 1918 1706 1922
rect 1718 1898 1722 1902
rect 1822 1928 1826 1932
rect 1846 1958 1850 1962
rect 1862 1958 1866 1962
rect 1894 2008 1898 2012
rect 1918 2008 1922 2012
rect 1926 2008 1930 2012
rect 1926 1998 1930 2002
rect 1950 1978 1954 1982
rect 1838 1938 1842 1942
rect 1582 1888 1586 1892
rect 1614 1888 1618 1892
rect 1766 1888 1770 1892
rect 1838 1888 1842 1892
rect 1874 1903 1878 1907
rect 1881 1903 1885 1907
rect 1598 1868 1602 1872
rect 1614 1868 1618 1872
rect 1494 1848 1498 1852
rect 1710 1878 1714 1882
rect 1590 1858 1594 1862
rect 1678 1858 1682 1862
rect 1606 1848 1610 1852
rect 1526 1838 1530 1842
rect 1582 1838 1586 1842
rect 1470 1828 1474 1832
rect 1462 1738 1466 1742
rect 1598 1818 1602 1822
rect 1542 1778 1546 1782
rect 1494 1758 1498 1762
rect 1542 1758 1546 1762
rect 1670 1848 1674 1852
rect 1686 1848 1690 1852
rect 1630 1778 1634 1782
rect 1686 1798 1690 1802
rect 1734 1868 1738 1872
rect 1750 1868 1754 1872
rect 1830 1868 1834 1872
rect 1742 1858 1746 1862
rect 1766 1858 1770 1862
rect 1750 1848 1754 1852
rect 1758 1808 1762 1812
rect 1718 1788 1722 1792
rect 1694 1768 1698 1772
rect 1718 1758 1722 1762
rect 1678 1748 1682 1752
rect 1702 1748 1706 1752
rect 1718 1748 1722 1752
rect 1734 1748 1738 1752
rect 1598 1738 1602 1742
rect 1566 1728 1570 1732
rect 1502 1698 1506 1702
rect 1614 1698 1618 1702
rect 1702 1728 1706 1732
rect 1622 1688 1626 1692
rect 1638 1688 1642 1692
rect 1486 1678 1490 1682
rect 1662 1678 1666 1682
rect 1670 1678 1674 1682
rect 1534 1668 1538 1672
rect 1654 1668 1658 1672
rect 1486 1648 1490 1652
rect 1494 1618 1498 1622
rect 1598 1658 1602 1662
rect 1678 1658 1682 1662
rect 1694 1658 1698 1662
rect 1678 1648 1682 1652
rect 1566 1598 1570 1602
rect 1870 1818 1874 1822
rect 1774 1758 1778 1762
rect 1766 1718 1770 1722
rect 1942 1948 1946 1952
rect 1910 1938 1914 1942
rect 1934 1938 1938 1942
rect 1902 1918 1906 1922
rect 1926 1918 1930 1922
rect 1918 1908 1922 1912
rect 1934 1888 1938 1892
rect 2046 2068 2050 2072
rect 2094 2068 2098 2072
rect 2022 2058 2026 2062
rect 2086 2058 2090 2062
rect 2118 2058 2122 2062
rect 2174 2058 2178 2062
rect 2198 2058 2202 2062
rect 2094 2048 2098 2052
rect 2190 2048 2194 2052
rect 1990 2038 1994 2042
rect 2150 2028 2154 2032
rect 2270 2118 2274 2122
rect 2286 2118 2290 2122
rect 2414 2148 2418 2152
rect 2462 2148 2466 2152
rect 2414 2138 2418 2142
rect 2430 2138 2434 2142
rect 2446 2138 2450 2142
rect 2502 2128 2506 2132
rect 2558 2158 2562 2162
rect 2622 2368 2626 2372
rect 2798 2588 2802 2592
rect 2758 2538 2762 2542
rect 2782 2538 2786 2542
rect 2790 2538 2794 2542
rect 2782 2518 2786 2522
rect 2750 2508 2754 2512
rect 2774 2508 2778 2512
rect 2790 2478 2794 2482
rect 2678 2448 2682 2452
rect 2670 2378 2674 2382
rect 2710 2378 2714 2382
rect 2734 2358 2738 2362
rect 2646 2328 2650 2332
rect 2686 2278 2690 2282
rect 2694 2268 2698 2272
rect 2574 2208 2578 2212
rect 2638 2258 2642 2262
rect 2678 2248 2682 2252
rect 2590 2198 2594 2202
rect 2582 2158 2586 2162
rect 2614 2158 2618 2162
rect 2398 2118 2402 2122
rect 2534 2098 2538 2102
rect 2262 2088 2266 2092
rect 2302 2088 2306 2092
rect 2366 2088 2370 2092
rect 2542 2088 2546 2092
rect 2294 2078 2298 2082
rect 2318 2078 2322 2082
rect 2326 2078 2330 2082
rect 2374 2078 2378 2082
rect 2422 2078 2426 2082
rect 2454 2078 2458 2082
rect 2502 2078 2506 2082
rect 2302 2068 2306 2072
rect 2246 2038 2250 2042
rect 2230 2018 2234 2022
rect 2030 1998 2034 2002
rect 2046 1998 2050 2002
rect 2038 1978 2042 1982
rect 2014 1968 2018 1972
rect 1982 1948 1986 1952
rect 2014 1938 2018 1942
rect 2030 1938 2034 1942
rect 1958 1908 1962 1912
rect 1998 1898 2002 1902
rect 2014 1898 2018 1902
rect 1974 1888 1978 1892
rect 1942 1868 1946 1872
rect 2054 1978 2058 1982
rect 2270 1978 2274 1982
rect 2134 1968 2138 1972
rect 2166 1968 2170 1972
rect 2230 1968 2234 1972
rect 2254 1968 2258 1972
rect 2062 1958 2066 1962
rect 2110 1958 2114 1962
rect 2142 1958 2146 1962
rect 2070 1938 2074 1942
rect 2094 1938 2098 1942
rect 2118 1938 2122 1942
rect 2150 1938 2154 1942
rect 2198 1938 2202 1942
rect 2062 1928 2066 1932
rect 2078 1928 2082 1932
rect 2134 1928 2138 1932
rect 2126 1918 2130 1922
rect 2086 1898 2090 1902
rect 2086 1888 2090 1892
rect 2102 1888 2106 1892
rect 2046 1868 2050 1872
rect 2062 1868 2066 1872
rect 1950 1858 1954 1862
rect 2046 1858 2050 1862
rect 2110 1878 2114 1882
rect 2094 1868 2098 1872
rect 2110 1858 2114 1862
rect 2174 1928 2178 1932
rect 2206 1928 2210 1932
rect 2158 1918 2162 1922
rect 2390 2068 2394 2072
rect 2334 2058 2338 2062
rect 2542 2068 2546 2072
rect 2574 2078 2578 2082
rect 2646 2148 2650 2152
rect 2694 2148 2698 2152
rect 2622 2108 2626 2112
rect 2566 2068 2570 2072
rect 2574 2068 2578 2072
rect 2446 2058 2450 2062
rect 2478 2058 2482 2062
rect 2494 2058 2498 2062
rect 2318 2048 2322 2052
rect 2326 2048 2330 2052
rect 2430 2048 2434 2052
rect 2462 2048 2466 2052
rect 2486 2038 2490 2042
rect 2510 2038 2514 2042
rect 2542 2048 2546 2052
rect 2574 2048 2578 2052
rect 2422 2028 2426 2032
rect 2526 2028 2530 2032
rect 2614 2048 2618 2052
rect 2334 2018 2338 2022
rect 2454 2018 2458 2022
rect 2598 2018 2602 2022
rect 2614 2018 2618 2022
rect 2278 1968 2282 1972
rect 2302 1968 2306 1972
rect 2310 1968 2314 1972
rect 2270 1958 2274 1962
rect 2222 1938 2226 1942
rect 2238 1938 2242 1942
rect 2254 1928 2258 1932
rect 2214 1918 2218 1922
rect 2166 1908 2170 1912
rect 2190 1908 2194 1912
rect 2190 1888 2194 1892
rect 2394 2003 2398 2007
rect 2401 2003 2405 2007
rect 2422 1998 2426 2002
rect 2358 1968 2362 1972
rect 2374 1968 2378 1972
rect 2294 1938 2298 1942
rect 2278 1928 2282 1932
rect 2302 1928 2306 1932
rect 2318 1918 2322 1922
rect 2238 1898 2242 1902
rect 2270 1898 2274 1902
rect 2278 1898 2282 1902
rect 2294 1888 2298 1892
rect 2150 1878 2154 1882
rect 2166 1858 2170 1862
rect 1926 1848 1930 1852
rect 1998 1848 2002 1852
rect 2102 1848 2106 1852
rect 1926 1838 1930 1842
rect 1998 1838 2002 1842
rect 1814 1788 1818 1792
rect 1838 1788 1842 1792
rect 1854 1748 1858 1752
rect 1878 1748 1882 1752
rect 1934 1818 1938 1822
rect 1950 1798 1954 1802
rect 1966 1798 1970 1802
rect 2014 1808 2018 1812
rect 2022 1808 2026 1812
rect 2014 1778 2018 1782
rect 1990 1758 1994 1762
rect 1974 1748 1978 1752
rect 1990 1748 1994 1752
rect 1806 1728 1810 1732
rect 1838 1728 1842 1732
rect 1854 1728 1858 1732
rect 1894 1718 1898 1722
rect 1790 1708 1794 1712
rect 1806 1708 1810 1712
rect 1782 1698 1786 1702
rect 1874 1703 1878 1707
rect 1881 1703 1885 1707
rect 1814 1688 1818 1692
rect 1846 1688 1850 1692
rect 1894 1688 1898 1692
rect 1902 1678 1906 1682
rect 1942 1678 1946 1682
rect 1798 1668 1802 1672
rect 1814 1668 1818 1672
rect 1934 1668 1938 1672
rect 1726 1658 1730 1662
rect 1718 1648 1722 1652
rect 1726 1648 1730 1652
rect 1790 1658 1794 1662
rect 1726 1638 1730 1642
rect 1742 1638 1746 1642
rect 1718 1608 1722 1612
rect 1694 1578 1698 1582
rect 1510 1568 1514 1572
rect 1646 1558 1650 1562
rect 1502 1548 1506 1552
rect 1614 1548 1618 1552
rect 1686 1548 1690 1552
rect 1494 1538 1498 1542
rect 1582 1538 1586 1542
rect 1686 1538 1690 1542
rect 1446 1528 1450 1532
rect 1374 1518 1378 1522
rect 1478 1518 1482 1522
rect 1510 1518 1514 1522
rect 1462 1498 1466 1502
rect 1334 1478 1338 1482
rect 1342 1478 1346 1482
rect 1494 1488 1498 1492
rect 1526 1488 1530 1492
rect 1486 1478 1490 1482
rect 1478 1468 1482 1472
rect 1334 1458 1338 1462
rect 1358 1458 1362 1462
rect 1326 1388 1330 1392
rect 1390 1448 1394 1452
rect 1370 1403 1374 1407
rect 1377 1403 1381 1407
rect 1334 1378 1338 1382
rect 1382 1358 1386 1362
rect 1390 1338 1394 1342
rect 1374 1298 1378 1302
rect 1350 1278 1354 1282
rect 1294 1268 1298 1272
rect 1310 1268 1314 1272
rect 1334 1268 1338 1272
rect 1350 1268 1354 1272
rect 1222 1258 1226 1262
rect 1254 1258 1258 1262
rect 1070 1228 1074 1232
rect 1078 1228 1082 1232
rect 1110 1228 1114 1232
rect 1150 1228 1154 1232
rect 1174 1228 1178 1232
rect 1190 1228 1194 1232
rect 1062 1198 1066 1202
rect 934 1178 938 1182
rect 1030 1158 1034 1162
rect 958 1148 962 1152
rect 1014 1138 1018 1142
rect 830 1118 834 1122
rect 878 1118 882 1122
rect 1510 1478 1514 1482
rect 1518 1478 1522 1482
rect 1622 1488 1626 1492
rect 1502 1468 1506 1472
rect 1518 1468 1522 1472
rect 1510 1458 1514 1462
rect 1478 1388 1482 1392
rect 1470 1368 1474 1372
rect 1462 1348 1466 1352
rect 1478 1328 1482 1332
rect 1398 1318 1402 1322
rect 1438 1318 1442 1322
rect 1422 1308 1426 1312
rect 1406 1278 1410 1282
rect 1470 1268 1474 1272
rect 1566 1388 1570 1392
rect 1702 1528 1706 1532
rect 1718 1508 1722 1512
rect 1710 1488 1714 1492
rect 1718 1478 1722 1482
rect 1782 1628 1786 1632
rect 1822 1658 1826 1662
rect 1910 1658 1914 1662
rect 1926 1658 1930 1662
rect 1878 1648 1882 1652
rect 1894 1648 1898 1652
rect 1878 1638 1882 1642
rect 1854 1608 1858 1612
rect 1854 1568 1858 1572
rect 1766 1558 1770 1562
rect 1758 1548 1762 1552
rect 1750 1538 1754 1542
rect 1766 1538 1770 1542
rect 1758 1528 1762 1532
rect 1822 1548 1826 1552
rect 1806 1528 1810 1532
rect 1798 1508 1802 1512
rect 1758 1478 1762 1482
rect 1790 1478 1794 1482
rect 1734 1468 1738 1472
rect 1750 1468 1754 1472
rect 1646 1458 1650 1462
rect 1710 1458 1714 1462
rect 1742 1458 1746 1462
rect 1646 1438 1650 1442
rect 1766 1438 1770 1442
rect 1630 1428 1634 1432
rect 1790 1438 1794 1442
rect 1654 1428 1658 1432
rect 1774 1428 1778 1432
rect 1630 1348 1634 1352
rect 1542 1338 1546 1342
rect 1614 1338 1618 1342
rect 1638 1318 1642 1322
rect 1686 1418 1690 1422
rect 1678 1338 1682 1342
rect 1654 1288 1658 1292
rect 1710 1408 1714 1412
rect 1814 1488 1818 1492
rect 1822 1478 1826 1482
rect 1878 1528 1882 1532
rect 1886 1528 1890 1532
rect 1822 1458 1826 1462
rect 1838 1418 1842 1422
rect 1758 1398 1762 1402
rect 1798 1398 1802 1402
rect 1874 1503 1878 1507
rect 1881 1503 1885 1507
rect 1918 1628 1922 1632
rect 1934 1568 1938 1572
rect 1926 1558 1930 1562
rect 1982 1728 1986 1732
rect 2038 1788 2042 1792
rect 2030 1768 2034 1772
rect 2014 1748 2018 1752
rect 1974 1688 1978 1692
rect 1958 1678 1962 1682
rect 1966 1668 1970 1672
rect 2006 1658 2010 1662
rect 1966 1648 1970 1652
rect 1990 1648 1994 1652
rect 2006 1648 2010 1652
rect 1974 1628 1978 1632
rect 2094 1808 2098 1812
rect 2126 1818 2130 1822
rect 2182 1818 2186 1822
rect 2134 1798 2138 1802
rect 2142 1798 2146 1802
rect 2142 1778 2146 1782
rect 2046 1708 2050 1712
rect 2038 1688 2042 1692
rect 2062 1678 2066 1682
rect 2022 1658 2026 1662
rect 2030 1608 2034 1612
rect 2006 1588 2010 1592
rect 2134 1748 2138 1752
rect 2118 1738 2122 1742
rect 2110 1698 2114 1702
rect 2110 1688 2114 1692
rect 2086 1678 2090 1682
rect 2158 1768 2162 1772
rect 2150 1758 2154 1762
rect 2342 1908 2346 1912
rect 2374 1938 2378 1942
rect 2374 1918 2378 1922
rect 2350 1898 2354 1902
rect 2462 1978 2466 1982
rect 2454 1968 2458 1972
rect 2430 1958 2434 1962
rect 2446 1958 2450 1962
rect 2510 1998 2514 2002
rect 2606 1998 2610 2002
rect 2678 2108 2682 2112
rect 2630 2048 2634 2052
rect 2662 2058 2666 2062
rect 2678 2058 2682 2062
rect 2686 2058 2690 2062
rect 2670 2048 2674 2052
rect 2782 2408 2786 2412
rect 2782 2398 2786 2402
rect 2766 2378 2770 2382
rect 2758 2298 2762 2302
rect 2750 2218 2754 2222
rect 2758 2158 2762 2162
rect 2718 2148 2722 2152
rect 2918 2758 2922 2762
rect 2906 2703 2910 2707
rect 2913 2703 2917 2707
rect 2902 2668 2906 2672
rect 2950 2748 2954 2752
rect 2966 2748 2970 2752
rect 2966 2728 2970 2732
rect 3150 2808 3154 2812
rect 3022 2798 3026 2802
rect 3246 2898 3250 2902
rect 3278 2928 3282 2932
rect 3302 2928 3306 2932
rect 3398 3018 3402 3022
rect 3418 3003 3422 3007
rect 3425 3003 3429 3007
rect 3422 2968 3426 2972
rect 3414 2958 3418 2962
rect 3406 2938 3410 2942
rect 3590 3128 3594 3132
rect 3662 3148 3666 3152
rect 3926 3318 3930 3322
rect 3918 3308 3922 3312
rect 3930 3303 3934 3307
rect 3937 3303 3941 3307
rect 3958 3368 3962 3372
rect 3974 3328 3978 3332
rect 4014 3378 4018 3382
rect 4142 3488 4146 3492
rect 4126 3468 4130 3472
rect 4094 3458 4098 3462
rect 4094 3418 4098 3422
rect 4078 3368 4082 3372
rect 4086 3368 4090 3372
rect 4054 3358 4058 3362
rect 4022 3348 4026 3352
rect 4086 3348 4090 3352
rect 3998 3308 4002 3312
rect 4078 3328 4082 3332
rect 4038 3318 4042 3322
rect 4030 3308 4034 3312
rect 4038 3308 4042 3312
rect 4054 3288 4058 3292
rect 4118 3388 4122 3392
rect 4110 3368 4114 3372
rect 4110 3358 4114 3362
rect 4102 3328 4106 3332
rect 4094 3308 4098 3312
rect 4342 3558 4346 3562
rect 4406 3558 4410 3562
rect 4350 3548 4354 3552
rect 4302 3528 4306 3532
rect 4150 3438 4154 3442
rect 4190 3488 4194 3492
rect 4174 3478 4178 3482
rect 4278 3488 4282 3492
rect 4182 3468 4186 3472
rect 4206 3468 4210 3472
rect 4230 3468 4234 3472
rect 4270 3468 4274 3472
rect 4182 3458 4186 3462
rect 4198 3458 4202 3462
rect 4206 3458 4210 3462
rect 4222 3458 4226 3462
rect 4190 3448 4194 3452
rect 4214 3438 4218 3442
rect 4174 3378 4178 3382
rect 4382 3548 4386 3552
rect 4398 3548 4402 3552
rect 4442 3603 4446 3607
rect 4449 3603 4453 3607
rect 4438 3588 4442 3592
rect 4358 3538 4362 3542
rect 4374 3538 4378 3542
rect 4430 3538 4434 3542
rect 4358 3488 4362 3492
rect 4302 3468 4306 3472
rect 4342 3468 4346 3472
rect 4294 3458 4298 3462
rect 4326 3458 4330 3462
rect 4254 3448 4258 3452
rect 4294 3448 4298 3452
rect 4334 3448 4338 3452
rect 4342 3448 4346 3452
rect 4246 3438 4250 3442
rect 4270 3438 4274 3442
rect 4406 3488 4410 3492
rect 4422 3488 4426 3492
rect 4390 3468 4394 3472
rect 4406 3468 4410 3472
rect 4374 3448 4378 3452
rect 4238 3398 4242 3402
rect 4238 3368 4242 3372
rect 4350 3348 4354 3352
rect 4398 3438 4402 3442
rect 4390 3428 4394 3432
rect 4390 3348 4394 3352
rect 4278 3338 4282 3342
rect 4126 3288 4130 3292
rect 4150 3258 4154 3262
rect 4246 3318 4250 3322
rect 4230 3298 4234 3302
rect 4326 3328 4330 3332
rect 4358 3328 4362 3332
rect 4390 3308 4394 3312
rect 4446 3578 4450 3582
rect 4462 3568 4466 3572
rect 4470 3558 4474 3562
rect 4446 3528 4450 3532
rect 4502 3638 4506 3642
rect 4574 3648 4578 3652
rect 4598 3648 4602 3652
rect 4526 3638 4530 3642
rect 4718 3648 4722 3652
rect 4678 3628 4682 3632
rect 4518 3578 4522 3582
rect 4558 3578 4562 3582
rect 4518 3568 4522 3572
rect 4486 3548 4490 3552
rect 4494 3548 4498 3552
rect 4526 3558 4530 3562
rect 4590 3568 4594 3572
rect 4582 3558 4586 3562
rect 4614 3558 4618 3562
rect 4670 3558 4674 3562
rect 4630 3548 4634 3552
rect 4638 3548 4642 3552
rect 4662 3548 4666 3552
rect 4510 3538 4514 3542
rect 4542 3538 4546 3542
rect 4566 3538 4570 3542
rect 4606 3538 4610 3542
rect 4646 3538 4650 3542
rect 4670 3538 4674 3542
rect 4494 3498 4498 3502
rect 4470 3488 4474 3492
rect 4486 3488 4490 3492
rect 4494 3488 4498 3492
rect 4470 3478 4474 3482
rect 4486 3468 4490 3472
rect 4494 3468 4498 3472
rect 4462 3458 4466 3462
rect 4550 3498 4554 3502
rect 4526 3488 4530 3492
rect 4542 3488 4546 3492
rect 4518 3478 4522 3482
rect 4462 3438 4466 3442
rect 4478 3438 4482 3442
rect 4442 3403 4446 3407
rect 4449 3403 4453 3407
rect 4574 3468 4578 3472
rect 4606 3468 4610 3472
rect 4694 3578 4698 3582
rect 4830 3668 4834 3672
rect 4766 3658 4770 3662
rect 4782 3658 4786 3662
rect 4766 3638 4770 3642
rect 4734 3618 4738 3622
rect 4814 3628 4818 3632
rect 4766 3568 4770 3572
rect 4702 3558 4706 3562
rect 4718 3558 4722 3562
rect 4734 3558 4738 3562
rect 4702 3538 4706 3542
rect 4662 3528 4666 3532
rect 4678 3528 4682 3532
rect 4710 3528 4714 3532
rect 4646 3478 4650 3482
rect 4630 3458 4634 3462
rect 4438 3358 4442 3362
rect 4542 3348 4546 3352
rect 4462 3338 4466 3342
rect 4438 3328 4442 3332
rect 4486 3338 4490 3342
rect 4542 3338 4546 3342
rect 4414 3298 4418 3302
rect 4470 3298 4474 3302
rect 4358 3288 4362 3292
rect 4214 3278 4218 3282
rect 4502 3308 4506 3312
rect 4534 3308 4538 3312
rect 4494 3298 4498 3302
rect 4382 3278 4386 3282
rect 4406 3278 4410 3282
rect 4486 3278 4490 3282
rect 4558 3318 4562 3322
rect 4550 3288 4554 3292
rect 4622 3448 4626 3452
rect 4590 3408 4594 3412
rect 4654 3398 4658 3402
rect 4598 3348 4602 3352
rect 4718 3508 4722 3512
rect 4846 3558 4850 3562
rect 4954 3703 4958 3707
rect 4961 3703 4965 3707
rect 5062 3688 5066 3692
rect 5150 3688 5154 3692
rect 4894 3678 4898 3682
rect 4998 3678 5002 3682
rect 4894 3658 4898 3662
rect 4982 3658 4986 3662
rect 4902 3648 4906 3652
rect 4990 3648 4994 3652
rect 4886 3618 4890 3622
rect 5038 3668 5042 3672
rect 5014 3648 5018 3652
rect 5006 3618 5010 3622
rect 4782 3548 4786 3552
rect 4806 3548 4810 3552
rect 4886 3548 4890 3552
rect 4918 3548 4922 3552
rect 4990 3548 4994 3552
rect 4822 3538 4826 3542
rect 4750 3518 4754 3522
rect 4766 3498 4770 3502
rect 4774 3488 4778 3492
rect 4798 3488 4802 3492
rect 4758 3468 4762 3472
rect 4862 3538 4866 3542
rect 4942 3538 4946 3542
rect 4838 3528 4842 3532
rect 4894 3528 4898 3532
rect 4918 3528 4922 3532
rect 4926 3528 4930 3532
rect 4854 3518 4858 3522
rect 4830 3498 4834 3502
rect 4854 3498 4858 3502
rect 4902 3488 4906 3492
rect 4846 3478 4850 3482
rect 4878 3478 4882 3482
rect 4718 3438 4722 3442
rect 4782 3448 4786 3452
rect 4726 3418 4730 3422
rect 4750 3418 4754 3422
rect 4694 3378 4698 3382
rect 4678 3358 4682 3362
rect 4614 3338 4618 3342
rect 4646 3338 4650 3342
rect 4614 3328 4618 3332
rect 4630 3328 4634 3332
rect 4606 3318 4610 3322
rect 4582 3308 4586 3312
rect 4606 3308 4610 3312
rect 4566 3278 4570 3282
rect 4326 3268 4330 3272
rect 4390 3268 4394 3272
rect 4510 3268 4514 3272
rect 3982 3248 3986 3252
rect 4038 3248 4042 3252
rect 4110 3248 4114 3252
rect 4166 3248 4170 3252
rect 4470 3258 4474 3262
rect 4550 3258 4554 3262
rect 4574 3258 4578 3262
rect 4270 3248 4274 3252
rect 4414 3238 4418 3242
rect 4462 3238 4466 3242
rect 4470 3238 4474 3242
rect 4398 3228 4402 3232
rect 4198 3208 4202 3212
rect 4214 3208 4218 3212
rect 4246 3208 4250 3212
rect 4334 3208 4338 3212
rect 3934 3188 3938 3192
rect 4158 3168 4162 3172
rect 4286 3158 4290 3162
rect 3774 3148 3778 3152
rect 3950 3148 3954 3152
rect 4014 3148 4018 3152
rect 4158 3148 4162 3152
rect 4182 3148 4186 3152
rect 3726 3138 3730 3142
rect 3870 3138 3874 3142
rect 3894 3138 3898 3142
rect 3990 3138 3994 3142
rect 4006 3138 4010 3142
rect 4070 3138 4074 3142
rect 3646 3128 3650 3132
rect 3830 3128 3834 3132
rect 3990 3128 3994 3132
rect 3582 3118 3586 3122
rect 3630 3118 3634 3122
rect 3502 3108 3506 3112
rect 3930 3103 3934 3107
rect 3937 3103 3941 3107
rect 3878 3098 3882 3102
rect 3814 3088 3818 3092
rect 4014 3088 4018 3092
rect 4086 3108 4090 3112
rect 3518 3078 3522 3082
rect 3542 3078 3546 3082
rect 3550 3078 3554 3082
rect 3590 3078 3594 3082
rect 3614 3078 3618 3082
rect 3638 3078 3642 3082
rect 3782 3078 3786 3082
rect 3950 3078 3954 3082
rect 3518 3068 3522 3072
rect 3486 3058 3490 3062
rect 3534 3058 3538 3062
rect 3494 3038 3498 3042
rect 3558 3068 3562 3072
rect 3598 3068 3602 3072
rect 3494 2978 3498 2982
rect 3510 2978 3514 2982
rect 3518 2978 3522 2982
rect 3526 2978 3530 2982
rect 3470 2958 3474 2962
rect 3366 2918 3370 2922
rect 3278 2908 3282 2912
rect 3302 2898 3306 2902
rect 3278 2878 3282 2882
rect 3294 2878 3298 2882
rect 3206 2868 3210 2872
rect 3198 2858 3202 2862
rect 3190 2848 3194 2852
rect 3206 2848 3210 2852
rect 3166 2798 3170 2802
rect 3118 2788 3122 2792
rect 3030 2768 3034 2772
rect 2990 2738 2994 2742
rect 2982 2718 2986 2722
rect 2878 2658 2882 2662
rect 2934 2658 2938 2662
rect 2838 2628 2842 2632
rect 2910 2628 2914 2632
rect 2974 2648 2978 2652
rect 2958 2628 2962 2632
rect 3150 2778 3154 2782
rect 3174 2778 3178 2782
rect 3198 2778 3202 2782
rect 3134 2748 3138 2752
rect 3038 2738 3042 2742
rect 3054 2738 3058 2742
rect 3038 2728 3042 2732
rect 3062 2718 3066 2722
rect 3126 2718 3130 2722
rect 3038 2698 3042 2702
rect 3102 2698 3106 2702
rect 3222 2828 3226 2832
rect 3238 2858 3242 2862
rect 3230 2808 3234 2812
rect 3222 2798 3226 2802
rect 3254 2868 3258 2872
rect 3486 2948 3490 2952
rect 3446 2928 3450 2932
rect 3534 2968 3538 2972
rect 3518 2948 3522 2952
rect 3494 2938 3498 2942
rect 3550 2948 3554 2952
rect 3558 2948 3562 2952
rect 3622 3068 3626 3072
rect 3694 3068 3698 3072
rect 3662 3058 3666 3062
rect 3686 3058 3690 3062
rect 3606 3048 3610 3052
rect 3622 3048 3626 3052
rect 3670 3048 3674 3052
rect 3702 3048 3706 3052
rect 3598 3028 3602 3032
rect 3582 2968 3586 2972
rect 3574 2958 3578 2962
rect 3718 3038 3722 3042
rect 3630 2988 3634 2992
rect 3678 2988 3682 2992
rect 3614 2958 3618 2962
rect 3670 2958 3674 2962
rect 3702 2958 3706 2962
rect 3630 2948 3634 2952
rect 3646 2948 3650 2952
rect 3558 2938 3562 2942
rect 3470 2928 3474 2932
rect 3430 2918 3434 2922
rect 3454 2918 3458 2922
rect 3494 2918 3498 2922
rect 3558 2918 3562 2922
rect 3422 2908 3426 2912
rect 3310 2878 3314 2882
rect 3254 2838 3258 2842
rect 3270 2828 3274 2832
rect 3462 2908 3466 2912
rect 3438 2898 3442 2902
rect 3470 2888 3474 2892
rect 3566 2888 3570 2892
rect 3438 2878 3442 2882
rect 3366 2868 3370 2872
rect 3686 2948 3690 2952
rect 3758 3058 3762 3062
rect 3838 3058 3842 3062
rect 3846 3048 3850 3052
rect 3870 3048 3874 3052
rect 3838 3038 3842 3042
rect 3790 3028 3794 3032
rect 4030 3068 4034 3072
rect 4134 3128 4138 3132
rect 4142 3128 4146 3132
rect 4166 3088 4170 3092
rect 4222 3138 4226 3142
rect 4230 3138 4234 3142
rect 4254 3128 4258 3132
rect 4270 3148 4274 3152
rect 4350 3158 4354 3162
rect 4318 3128 4322 3132
rect 4270 3118 4274 3122
rect 4262 3108 4266 3112
rect 4230 3088 4234 3092
rect 4094 3068 4098 3072
rect 3902 3058 3906 3062
rect 3926 3058 3930 3062
rect 4006 3058 4010 3062
rect 4038 3058 4042 3062
rect 4054 3058 4058 3062
rect 4070 3058 4074 3062
rect 4086 3058 4090 3062
rect 4158 3058 4162 3062
rect 4166 3058 4170 3062
rect 3974 3048 3978 3052
rect 4046 3048 4050 3052
rect 4110 3048 4114 3052
rect 3894 3038 3898 3042
rect 4078 3038 4082 3042
rect 4110 3038 4114 3042
rect 4158 3038 4162 3042
rect 4158 3028 4162 3032
rect 4110 3018 4114 3022
rect 3734 2978 3738 2982
rect 3750 2978 3754 2982
rect 3766 2978 3770 2982
rect 3734 2948 3738 2952
rect 3614 2938 3618 2942
rect 3662 2938 3666 2942
rect 3630 2928 3634 2932
rect 3710 2938 3714 2942
rect 3638 2918 3642 2922
rect 3654 2918 3658 2922
rect 3694 2918 3698 2922
rect 3598 2908 3602 2912
rect 3622 2908 3626 2912
rect 3638 2898 3642 2902
rect 3798 2968 3802 2972
rect 4442 3203 4446 3207
rect 4449 3203 4453 3207
rect 4422 3178 4426 3182
rect 4550 3168 4554 3172
rect 4462 3108 4466 3112
rect 4510 3118 4514 3122
rect 4438 3088 4442 3092
rect 4462 3088 4466 3092
rect 4534 3088 4538 3092
rect 4342 3078 4346 3082
rect 4358 3078 4362 3082
rect 4438 3078 4442 3082
rect 4302 3068 4306 3072
rect 4366 3068 4370 3072
rect 4406 3068 4410 3072
rect 4494 3068 4498 3072
rect 4510 3068 4514 3072
rect 4670 3328 4674 3332
rect 4710 3318 4714 3322
rect 4662 3288 4666 3292
rect 4654 3278 4658 3282
rect 4686 3278 4690 3282
rect 4694 3278 4698 3282
rect 4798 3448 4802 3452
rect 4814 3448 4818 3452
rect 4830 3448 4834 3452
rect 4798 3408 4802 3412
rect 4734 3338 4738 3342
rect 4790 3338 4794 3342
rect 4814 3368 4818 3372
rect 4798 3308 4802 3312
rect 4838 3358 4842 3362
rect 5030 3648 5034 3652
rect 5094 3648 5098 3652
rect 5078 3628 5082 3632
rect 5070 3618 5074 3622
rect 5062 3568 5066 3572
rect 5022 3558 5026 3562
rect 4982 3528 4986 3532
rect 4950 3518 4954 3522
rect 4954 3503 4958 3507
rect 4961 3503 4965 3507
rect 4998 3488 5002 3492
rect 5006 3478 5010 3482
rect 4854 3468 4858 3472
rect 4886 3468 4890 3472
rect 4926 3468 4930 3472
rect 5006 3468 5010 3472
rect 5022 3468 5026 3472
rect 4854 3368 4858 3372
rect 4894 3458 4898 3462
rect 4934 3458 4938 3462
rect 4998 3458 5002 3462
rect 4886 3448 4890 3452
rect 4878 3438 4882 3442
rect 4910 3368 4914 3372
rect 4902 3358 4906 3362
rect 4886 3348 4890 3352
rect 4926 3348 4930 3352
rect 4838 3328 4842 3332
rect 4822 3318 4826 3322
rect 4854 3318 4858 3322
rect 4726 3298 4730 3302
rect 4774 3298 4778 3302
rect 4814 3298 4818 3302
rect 4838 3298 4842 3302
rect 4758 3288 4762 3292
rect 4742 3278 4746 3282
rect 4734 3268 4738 3272
rect 4742 3268 4746 3272
rect 4630 3258 4634 3262
rect 4670 3258 4674 3262
rect 4614 3248 4618 3252
rect 4726 3248 4730 3252
rect 4662 3158 4666 3162
rect 4630 3148 4634 3152
rect 5014 3448 5018 3452
rect 5078 3548 5082 3552
rect 5086 3548 5090 3552
rect 5126 3548 5130 3552
rect 5062 3478 5066 3482
rect 5222 3618 5226 3622
rect 5214 3568 5218 3572
rect 5158 3558 5162 3562
rect 5094 3488 5098 3492
rect 5030 3428 5034 3432
rect 4982 3368 4986 3372
rect 5078 3368 5082 3372
rect 4982 3358 4986 3362
rect 4990 3358 4994 3362
rect 5006 3358 5010 3362
rect 5022 3358 5026 3362
rect 5006 3348 5010 3352
rect 4878 3338 4882 3342
rect 4902 3338 4906 3342
rect 4934 3338 4938 3342
rect 5046 3338 5050 3342
rect 4870 3328 4874 3332
rect 4966 3328 4970 3332
rect 4894 3308 4898 3312
rect 4870 3298 4874 3302
rect 4862 3288 4866 3292
rect 4854 3278 4858 3282
rect 4954 3303 4958 3307
rect 4961 3303 4965 3307
rect 4902 3288 4906 3292
rect 4934 3288 4938 3292
rect 4894 3278 4898 3282
rect 5238 3698 5242 3702
rect 5254 3658 5258 3662
rect 5246 3648 5250 3652
rect 5278 3648 5282 3652
rect 5302 3568 5306 3572
rect 5294 3558 5298 3562
rect 5246 3548 5250 3552
rect 5278 3548 5282 3552
rect 5262 3528 5266 3532
rect 5206 3478 5210 3482
rect 5110 3458 5114 3462
rect 5262 3468 5266 3472
rect 5142 3448 5146 3452
rect 5270 3448 5274 3452
rect 5262 3438 5266 3442
rect 5110 3378 5114 3382
rect 5102 3368 5106 3372
rect 5126 3368 5130 3372
rect 5142 3368 5146 3372
rect 5182 3358 5186 3362
rect 5094 3348 5098 3352
rect 5102 3348 5106 3352
rect 5278 3428 5282 3432
rect 5238 3388 5242 3392
rect 5270 3368 5274 3372
rect 5278 3358 5282 3362
rect 5286 3358 5290 3362
rect 5086 3338 5090 3342
rect 5102 3338 5106 3342
rect 5134 3338 5138 3342
rect 5246 3338 5250 3342
rect 5190 3328 5194 3332
rect 5150 3318 5154 3322
rect 4918 3278 4922 3282
rect 4942 3278 4946 3282
rect 4950 3278 4954 3282
rect 4998 3278 5002 3282
rect 5022 3278 5026 3282
rect 5062 3278 5066 3282
rect 5110 3278 5114 3282
rect 5142 3278 5146 3282
rect 5206 3278 5210 3282
rect 4894 3268 4898 3272
rect 4910 3268 4914 3272
rect 4934 3268 4938 3272
rect 4958 3268 4962 3272
rect 5046 3268 5050 3272
rect 4830 3258 4834 3262
rect 4998 3258 5002 3262
rect 4806 3248 4810 3252
rect 4982 3248 4986 3252
rect 4910 3218 4914 3222
rect 4758 3158 4762 3162
rect 4862 3188 4866 3192
rect 4846 3168 4850 3172
rect 4862 3158 4866 3162
rect 4870 3158 4874 3162
rect 4774 3148 4778 3152
rect 4790 3148 4794 3152
rect 4694 3138 4698 3142
rect 4622 3118 4626 3122
rect 4550 3088 4554 3092
rect 4590 3078 4594 3082
rect 4638 3088 4642 3092
rect 4622 3068 4626 3072
rect 4334 3058 4338 3062
rect 4398 3058 4402 3062
rect 4526 3058 4530 3062
rect 4278 3038 4282 3042
rect 4190 3028 4194 3032
rect 4246 3028 4250 3032
rect 4326 3048 4330 3052
rect 4318 3028 4322 3032
rect 3806 2958 3810 2962
rect 4006 2958 4010 2962
rect 4086 2958 4090 2962
rect 4134 2958 4138 2962
rect 3838 2948 3842 2952
rect 3910 2948 3914 2952
rect 3758 2928 3762 2932
rect 3846 2938 3850 2942
rect 3902 2928 3906 2932
rect 3798 2918 3802 2922
rect 3822 2918 3826 2922
rect 3846 2918 3850 2922
rect 3950 2918 3954 2922
rect 3742 2898 3746 2902
rect 3726 2888 3730 2892
rect 3830 2908 3834 2912
rect 3654 2878 3658 2882
rect 3710 2878 3714 2882
rect 3782 2878 3786 2882
rect 3694 2868 3698 2872
rect 3326 2858 3330 2862
rect 3454 2858 3458 2862
rect 3470 2858 3474 2862
rect 3510 2858 3514 2862
rect 3670 2858 3674 2862
rect 3678 2858 3682 2862
rect 3542 2848 3546 2852
rect 3638 2848 3642 2852
rect 3646 2848 3650 2852
rect 3670 2848 3674 2852
rect 3614 2838 3618 2842
rect 3686 2838 3690 2842
rect 3694 2828 3698 2832
rect 3534 2818 3538 2822
rect 3334 2808 3338 2812
rect 3470 2808 3474 2812
rect 3494 2808 3498 2812
rect 3418 2803 3422 2807
rect 3425 2803 3429 2807
rect 3806 2868 3810 2872
rect 3814 2868 3818 2872
rect 3930 2903 3934 2907
rect 3937 2903 3941 2907
rect 3846 2888 3850 2892
rect 3870 2868 3874 2872
rect 3894 2868 3898 2872
rect 3734 2858 3738 2862
rect 3862 2848 3866 2852
rect 3766 2838 3770 2842
rect 3878 2828 3882 2832
rect 3782 2818 3786 2822
rect 3454 2788 3458 2792
rect 3710 2788 3714 2792
rect 3310 2778 3314 2782
rect 3254 2768 3258 2772
rect 3278 2748 3282 2752
rect 3166 2738 3170 2742
rect 3174 2738 3178 2742
rect 3206 2738 3210 2742
rect 3174 2728 3178 2732
rect 3190 2728 3194 2732
rect 3158 2718 3162 2722
rect 3158 2708 3162 2712
rect 3006 2678 3010 2682
rect 3094 2678 3098 2682
rect 3118 2678 3122 2682
rect 3062 2628 3066 2632
rect 2942 2618 2946 2622
rect 2982 2618 2986 2622
rect 3054 2618 3058 2622
rect 3030 2598 3034 2602
rect 2846 2548 2850 2552
rect 2886 2548 2890 2552
rect 2838 2538 2842 2542
rect 2862 2538 2866 2542
rect 2814 2528 2818 2532
rect 2806 2508 2810 2512
rect 2830 2498 2834 2502
rect 2822 2448 2826 2452
rect 2798 2398 2802 2402
rect 3110 2598 3114 2602
rect 3126 2598 3130 2602
rect 3126 2568 3130 2572
rect 3078 2558 3082 2562
rect 3102 2558 3106 2562
rect 3150 2628 3154 2632
rect 3190 2698 3194 2702
rect 3174 2668 3178 2672
rect 3150 2578 3154 2582
rect 3230 2698 3234 2702
rect 3774 2778 3778 2782
rect 3734 2768 3738 2772
rect 3766 2768 3770 2772
rect 3486 2758 3490 2762
rect 3606 2758 3610 2762
rect 3638 2758 3642 2762
rect 3662 2758 3666 2762
rect 3678 2758 3682 2762
rect 3294 2748 3298 2752
rect 3342 2748 3346 2752
rect 3406 2748 3410 2752
rect 3286 2728 3290 2732
rect 3246 2708 3250 2712
rect 3326 2708 3330 2712
rect 3542 2748 3546 2752
rect 3606 2748 3610 2752
rect 3510 2718 3514 2722
rect 3566 2718 3570 2722
rect 3630 2728 3634 2732
rect 3462 2708 3466 2712
rect 3582 2708 3586 2712
rect 3310 2698 3314 2702
rect 3374 2698 3378 2702
rect 3214 2668 3218 2672
rect 3230 2668 3234 2672
rect 3238 2668 3242 2672
rect 3254 2668 3258 2672
rect 3190 2658 3194 2662
rect 3454 2688 3458 2692
rect 3462 2688 3466 2692
rect 3614 2678 3618 2682
rect 3638 2718 3642 2722
rect 3294 2668 3298 2672
rect 3630 2668 3634 2672
rect 3310 2658 3314 2662
rect 3214 2648 3218 2652
rect 3262 2648 3266 2652
rect 3278 2648 3282 2652
rect 3326 2648 3330 2652
rect 3174 2638 3178 2642
rect 3302 2638 3306 2642
rect 3222 2628 3226 2632
rect 3294 2628 3298 2632
rect 3262 2618 3266 2622
rect 3198 2558 3202 2562
rect 3062 2548 3066 2552
rect 3086 2548 3090 2552
rect 3118 2548 3122 2552
rect 3150 2548 3154 2552
rect 3342 2638 3346 2642
rect 3502 2658 3506 2662
rect 3518 2658 3522 2662
rect 3414 2648 3418 2652
rect 3382 2608 3386 2612
rect 3418 2603 3422 2607
rect 3425 2603 3429 2607
rect 3542 2558 3546 2562
rect 2894 2538 2898 2542
rect 2966 2538 2970 2542
rect 3038 2538 3042 2542
rect 3070 2538 3074 2542
rect 3110 2538 3114 2542
rect 2846 2478 2850 2482
rect 2906 2503 2910 2507
rect 2913 2503 2917 2507
rect 2974 2478 2978 2482
rect 3022 2468 3026 2472
rect 2830 2438 2834 2442
rect 2854 2438 2858 2442
rect 2806 2368 2810 2372
rect 3150 2518 3154 2522
rect 3054 2498 3058 2502
rect 3086 2478 3090 2482
rect 3246 2498 3250 2502
rect 3374 2538 3378 2542
rect 3294 2488 3298 2492
rect 3038 2458 3042 2462
rect 3070 2458 3074 2462
rect 3166 2458 3170 2462
rect 3350 2478 3354 2482
rect 3278 2458 3282 2462
rect 3342 2458 3346 2462
rect 3366 2468 3370 2472
rect 3182 2448 3186 2452
rect 3310 2448 3314 2452
rect 3342 2448 3346 2452
rect 3390 2448 3394 2452
rect 2990 2438 2994 2442
rect 3382 2438 3386 2442
rect 2894 2408 2898 2412
rect 2870 2398 2874 2402
rect 2990 2388 2994 2392
rect 3174 2388 3178 2392
rect 3214 2388 3218 2392
rect 2950 2378 2954 2382
rect 3014 2378 3018 2382
rect 3054 2378 3058 2382
rect 2910 2368 2914 2372
rect 2798 2358 2802 2362
rect 2878 2358 2882 2362
rect 2950 2358 2954 2362
rect 2966 2358 2970 2362
rect 2822 2338 2826 2342
rect 2790 2268 2794 2272
rect 2798 2258 2802 2262
rect 2822 2198 2826 2202
rect 2814 2148 2818 2152
rect 2750 2128 2754 2132
rect 2886 2348 2890 2352
rect 2926 2348 2930 2352
rect 2942 2348 2946 2352
rect 2854 2338 2858 2342
rect 2862 2338 2866 2342
rect 2846 2298 2850 2302
rect 2982 2340 2986 2344
rect 3038 2358 3042 2362
rect 3062 2358 3066 2362
rect 3142 2358 3146 2362
rect 3150 2358 3154 2362
rect 2998 2338 3002 2342
rect 3030 2338 3034 2342
rect 2870 2328 2874 2332
rect 2918 2328 2922 2332
rect 2906 2303 2910 2307
rect 2913 2303 2917 2307
rect 2886 2288 2890 2292
rect 2918 2278 2922 2282
rect 2974 2278 2978 2282
rect 2902 2268 2906 2272
rect 2958 2258 2962 2262
rect 2966 2258 2970 2262
rect 2982 2258 2986 2262
rect 2966 2238 2970 2242
rect 2902 2218 2906 2222
rect 2862 2198 2866 2202
rect 2870 2198 2874 2202
rect 2854 2178 2858 2182
rect 2886 2178 2890 2182
rect 2846 2158 2850 2162
rect 2870 2158 2874 2162
rect 2718 2118 2722 2122
rect 2726 2118 2730 2122
rect 2814 2118 2818 2122
rect 2702 2098 2706 2102
rect 2702 2058 2706 2062
rect 2646 2038 2650 2042
rect 2686 2038 2690 2042
rect 2694 2038 2698 2042
rect 2670 2028 2674 2032
rect 2694 2028 2698 2032
rect 2630 2008 2634 2012
rect 2614 1978 2618 1982
rect 2622 1978 2626 1982
rect 2470 1958 2474 1962
rect 2454 1938 2458 1942
rect 2462 1928 2466 1932
rect 2534 1928 2538 1932
rect 2438 1908 2442 1912
rect 2510 1918 2514 1922
rect 2470 1898 2474 1902
rect 2438 1888 2442 1892
rect 2566 1878 2570 1882
rect 2214 1868 2218 1872
rect 2230 1868 2234 1872
rect 2270 1866 2274 1870
rect 2294 1868 2298 1872
rect 2422 1868 2426 1872
rect 2374 1858 2378 1862
rect 2302 1838 2306 1842
rect 2270 1818 2274 1822
rect 2198 1798 2202 1802
rect 2190 1768 2194 1772
rect 2326 1808 2330 1812
rect 2166 1758 2170 1762
rect 2198 1758 2202 1762
rect 2294 1758 2298 1762
rect 2310 1758 2314 1762
rect 2318 1758 2322 1762
rect 2414 1858 2418 1862
rect 2366 1848 2370 1852
rect 2382 1848 2386 1852
rect 2398 1818 2402 1822
rect 2394 1803 2398 1807
rect 2401 1803 2405 1807
rect 2446 1848 2450 1852
rect 2430 1818 2434 1822
rect 2390 1768 2394 1772
rect 2414 1768 2418 1772
rect 2350 1758 2354 1762
rect 2366 1758 2370 1762
rect 2342 1748 2346 1752
rect 2262 1738 2266 1742
rect 2318 1738 2322 1742
rect 2206 1728 2210 1732
rect 2278 1728 2282 1732
rect 2294 1728 2298 1732
rect 2158 1708 2162 1712
rect 2142 1678 2146 1682
rect 2166 1688 2170 1692
rect 2166 1678 2170 1682
rect 2086 1658 2090 1662
rect 2078 1578 2082 1582
rect 1950 1558 1954 1562
rect 1942 1548 1946 1552
rect 1958 1548 1962 1552
rect 2054 1548 2058 1552
rect 1990 1538 1994 1542
rect 2038 1538 2042 1542
rect 2230 1718 2234 1722
rect 2238 1718 2242 1722
rect 2182 1698 2186 1702
rect 2206 1688 2210 1692
rect 2182 1668 2186 1672
rect 2222 1678 2226 1682
rect 2222 1668 2226 1672
rect 2254 1688 2258 1692
rect 2262 1688 2266 1692
rect 2270 1678 2274 1682
rect 2198 1648 2202 1652
rect 2126 1628 2130 1632
rect 2214 1628 2218 1632
rect 2166 1618 2170 1622
rect 2142 1598 2146 1602
rect 2102 1558 2106 1562
rect 2094 1548 2098 1552
rect 2062 1538 2066 1542
rect 2086 1538 2090 1542
rect 1918 1528 1922 1532
rect 1966 1528 1970 1532
rect 1990 1528 1994 1532
rect 2046 1528 2050 1532
rect 2078 1528 2082 1532
rect 1990 1518 1994 1522
rect 2022 1508 2026 1512
rect 2070 1498 2074 1502
rect 1894 1488 1898 1492
rect 1926 1488 1930 1492
rect 1902 1478 1906 1482
rect 1974 1478 1978 1482
rect 1982 1478 1986 1482
rect 1862 1458 1866 1462
rect 1806 1388 1810 1392
rect 1854 1388 1858 1392
rect 1838 1378 1842 1382
rect 1910 1468 1914 1472
rect 1934 1468 1938 1472
rect 1910 1458 1914 1462
rect 1958 1458 1962 1462
rect 1894 1438 1898 1442
rect 1870 1418 1874 1422
rect 1862 1368 1866 1372
rect 1878 1348 1882 1352
rect 1926 1448 1930 1452
rect 1910 1428 1914 1432
rect 1950 1408 1954 1412
rect 2006 1468 2010 1472
rect 2022 1468 2026 1472
rect 2038 1468 2042 1472
rect 2102 1528 2106 1532
rect 2134 1548 2138 1552
rect 2206 1548 2210 1552
rect 2158 1538 2162 1542
rect 2182 1528 2186 1532
rect 2110 1508 2114 1512
rect 2094 1498 2098 1502
rect 2110 1498 2114 1502
rect 2102 1488 2106 1492
rect 2118 1488 2122 1492
rect 2142 1488 2146 1492
rect 2182 1488 2186 1492
rect 2102 1468 2106 1472
rect 2030 1458 2034 1462
rect 2006 1448 2010 1452
rect 2022 1448 2026 1452
rect 1982 1438 1986 1442
rect 2062 1418 2066 1422
rect 2038 1398 2042 1402
rect 1934 1388 1938 1392
rect 1942 1388 1946 1392
rect 1974 1388 1978 1392
rect 1918 1378 1922 1382
rect 1926 1378 1930 1382
rect 1918 1348 1922 1352
rect 1798 1338 1802 1342
rect 1878 1338 1882 1342
rect 1902 1338 1906 1342
rect 1934 1338 1938 1342
rect 1734 1318 1738 1322
rect 1718 1298 1722 1302
rect 1518 1278 1522 1282
rect 1534 1278 1538 1282
rect 1678 1278 1682 1282
rect 1734 1278 1738 1282
rect 1302 1258 1306 1262
rect 1326 1258 1330 1262
rect 1390 1258 1394 1262
rect 1558 1268 1562 1272
rect 1606 1268 1610 1272
rect 1622 1268 1626 1272
rect 1638 1268 1642 1272
rect 1662 1268 1666 1272
rect 1678 1268 1682 1272
rect 1582 1258 1586 1262
rect 1318 1248 1322 1252
rect 1334 1248 1338 1252
rect 1486 1248 1490 1252
rect 1518 1248 1522 1252
rect 1542 1248 1546 1252
rect 1606 1248 1610 1252
rect 1590 1238 1594 1242
rect 1286 1218 1290 1222
rect 1478 1218 1482 1222
rect 1566 1218 1570 1222
rect 1086 1198 1090 1202
rect 1198 1198 1202 1202
rect 1370 1203 1374 1207
rect 1377 1203 1381 1207
rect 1142 1168 1146 1172
rect 1262 1168 1266 1172
rect 1238 1158 1242 1162
rect 974 1118 978 1122
rect 782 1098 786 1102
rect 858 1103 862 1107
rect 865 1103 869 1107
rect 910 1098 914 1102
rect 830 1088 834 1092
rect 710 1068 714 1072
rect 830 1068 834 1072
rect 942 1098 946 1102
rect 1070 1118 1074 1122
rect 1494 1158 1498 1162
rect 1094 1098 1098 1102
rect 1062 1088 1066 1092
rect 1126 1108 1130 1112
rect 1286 1148 1290 1152
rect 1134 1098 1138 1102
rect 1126 1088 1130 1092
rect 1134 1088 1138 1092
rect 966 1078 970 1082
rect 1014 1078 1018 1082
rect 1046 1078 1050 1082
rect 1102 1078 1106 1082
rect 726 1058 730 1062
rect 742 1058 746 1062
rect 766 1058 770 1062
rect 926 1058 930 1062
rect 934 1058 938 1062
rect 630 1048 634 1052
rect 750 1048 754 1052
rect 622 1038 626 1042
rect 830 1038 834 1042
rect 598 1008 602 1012
rect 550 958 554 962
rect 574 958 578 962
rect 614 958 618 962
rect 542 948 546 952
rect 566 948 570 952
rect 582 948 586 952
rect 1054 1068 1058 1072
rect 958 1048 962 1052
rect 990 1048 994 1052
rect 1030 1048 1034 1052
rect 998 1038 1002 1042
rect 1030 1038 1034 1042
rect 1046 1038 1050 1042
rect 1014 1028 1018 1032
rect 686 1018 690 1022
rect 710 1018 714 1022
rect 846 1018 850 1022
rect 630 978 634 982
rect 646 968 650 972
rect 678 968 682 972
rect 638 948 642 952
rect 526 938 530 942
rect 550 938 554 942
rect 662 938 666 942
rect 534 928 538 932
rect 558 928 562 932
rect 614 898 618 902
rect 550 888 554 892
rect 558 888 562 892
rect 502 878 506 882
rect 542 878 546 882
rect 606 878 610 882
rect 494 868 498 872
rect 718 948 722 952
rect 678 938 682 942
rect 670 908 674 912
rect 670 888 674 892
rect 654 878 658 882
rect 734 898 738 902
rect 718 888 722 892
rect 710 878 714 882
rect 638 868 642 872
rect 534 858 538 862
rect 590 858 594 862
rect 646 858 650 862
rect 694 858 698 862
rect 774 888 778 892
rect 734 858 738 862
rect 598 848 602 852
rect 622 848 626 852
rect 686 848 690 852
rect 358 838 362 842
rect 38 747 42 751
rect 110 748 114 752
rect 126 748 130 752
rect 182 748 186 752
rect 94 708 98 712
rect 150 738 154 742
rect 174 738 178 742
rect 142 688 146 692
rect 134 668 138 672
rect 174 708 178 712
rect 190 708 194 712
rect 166 678 170 682
rect 638 818 642 822
rect 346 803 350 807
rect 353 803 357 807
rect 294 778 298 782
rect 206 758 210 762
rect 238 758 242 762
rect 270 758 274 762
rect 222 748 226 752
rect 214 738 218 742
rect 206 718 210 722
rect 238 718 242 722
rect 318 728 322 732
rect 278 708 282 712
rect 230 698 234 702
rect 262 698 266 702
rect 206 678 210 682
rect 262 678 266 682
rect 182 668 186 672
rect 198 668 202 672
rect 238 668 242 672
rect 150 658 154 662
rect 198 658 202 662
rect 222 658 226 662
rect 110 648 114 652
rect 222 648 226 652
rect 62 588 66 592
rect 62 568 66 572
rect 38 508 42 512
rect 222 628 226 632
rect 182 568 186 572
rect 206 568 210 572
rect 158 558 162 562
rect 190 558 194 562
rect 118 508 122 512
rect 302 678 306 682
rect 294 668 298 672
rect 262 658 266 662
rect 278 658 282 662
rect 342 748 346 752
rect 414 768 418 772
rect 454 768 458 772
rect 478 768 482 772
rect 486 768 490 772
rect 686 768 690 772
rect 374 748 378 752
rect 334 738 338 742
rect 350 738 354 742
rect 374 728 378 732
rect 334 708 338 712
rect 358 698 362 702
rect 438 748 442 752
rect 446 728 450 732
rect 438 718 442 722
rect 446 698 450 702
rect 478 728 482 732
rect 446 688 450 692
rect 390 678 394 682
rect 502 758 506 762
rect 518 758 522 762
rect 510 748 514 752
rect 550 748 554 752
rect 590 748 594 752
rect 502 728 506 732
rect 526 728 530 732
rect 534 728 538 732
rect 558 728 562 732
rect 590 728 594 732
rect 1030 978 1034 982
rect 846 968 850 972
rect 950 968 954 972
rect 958 968 962 972
rect 974 968 978 972
rect 998 968 1002 972
rect 1014 968 1018 972
rect 1046 968 1050 972
rect 798 958 802 962
rect 838 958 842 962
rect 918 958 922 962
rect 838 938 842 942
rect 846 938 850 942
rect 858 903 862 907
rect 865 903 869 907
rect 902 938 906 942
rect 926 948 930 952
rect 942 948 946 952
rect 862 878 866 882
rect 918 878 922 882
rect 974 958 978 962
rect 966 948 970 952
rect 966 878 970 882
rect 1150 1108 1154 1112
rect 1286 1138 1290 1142
rect 1182 1128 1186 1132
rect 1230 1128 1234 1132
rect 1166 1118 1170 1122
rect 1158 1098 1162 1102
rect 1094 1068 1098 1072
rect 1150 1068 1154 1072
rect 1070 1058 1074 1062
rect 1070 1048 1074 1052
rect 1110 1048 1114 1052
rect 1166 1058 1170 1062
rect 1262 1098 1266 1102
rect 1230 1078 1234 1082
rect 1398 1148 1402 1152
rect 1446 1148 1450 1152
rect 1334 1138 1338 1142
rect 1302 1128 1306 1132
rect 1398 1128 1402 1132
rect 1390 1118 1394 1122
rect 1366 1098 1370 1102
rect 1270 1078 1274 1082
rect 1198 1068 1202 1072
rect 1310 1068 1314 1072
rect 1142 1048 1146 1052
rect 1342 1068 1346 1072
rect 1198 1058 1202 1062
rect 1214 1058 1218 1062
rect 1350 1058 1354 1062
rect 1270 1048 1274 1052
rect 1286 1048 1290 1052
rect 1302 1048 1306 1052
rect 1182 1038 1186 1042
rect 1214 1038 1218 1042
rect 1118 1028 1122 1032
rect 1230 978 1234 982
rect 1094 968 1098 972
rect 1086 958 1090 962
rect 1206 958 1210 962
rect 1030 948 1034 952
rect 1062 948 1066 952
rect 1134 948 1138 952
rect 1174 948 1178 952
rect 1230 948 1234 952
rect 1358 1028 1362 1032
rect 1370 1003 1374 1007
rect 1377 1003 1381 1007
rect 1510 1148 1514 1152
rect 1630 1258 1634 1262
rect 1654 1258 1658 1262
rect 1646 1248 1650 1252
rect 1662 1248 1666 1252
rect 1614 1188 1618 1192
rect 1598 1178 1602 1182
rect 1606 1168 1610 1172
rect 1646 1168 1650 1172
rect 1590 1138 1594 1142
rect 1614 1138 1618 1142
rect 1622 1138 1626 1142
rect 1454 1128 1458 1132
rect 1422 1118 1426 1122
rect 1438 1118 1442 1122
rect 1454 1108 1458 1112
rect 1430 1088 1434 1092
rect 1446 1068 1450 1072
rect 1446 1058 1450 1062
rect 1462 1088 1466 1092
rect 1470 1058 1474 1062
rect 1414 1048 1418 1052
rect 1422 1048 1426 1052
rect 1430 1038 1434 1042
rect 1414 998 1418 1002
rect 1302 988 1306 992
rect 1406 988 1410 992
rect 1430 978 1434 982
rect 1318 968 1322 972
rect 1462 998 1466 1002
rect 1374 958 1378 962
rect 1454 948 1458 952
rect 990 938 994 942
rect 942 868 946 872
rect 958 868 962 872
rect 790 858 794 862
rect 854 848 858 852
rect 886 848 890 852
rect 918 848 922 852
rect 950 848 954 852
rect 830 778 834 782
rect 798 758 802 762
rect 718 748 722 752
rect 814 748 818 752
rect 710 738 714 742
rect 950 738 954 742
rect 654 728 658 732
rect 566 718 570 722
rect 598 718 602 722
rect 630 718 634 722
rect 662 718 666 722
rect 550 708 554 712
rect 542 688 546 692
rect 406 678 410 682
rect 470 678 474 682
rect 494 678 498 682
rect 310 668 314 672
rect 326 668 330 672
rect 358 668 362 672
rect 390 668 394 672
rect 398 668 402 672
rect 286 648 290 652
rect 318 648 322 652
rect 270 638 274 642
rect 422 658 426 662
rect 334 648 338 652
rect 366 648 370 652
rect 398 648 402 652
rect 438 648 442 652
rect 326 628 330 632
rect 346 603 350 607
rect 353 603 357 607
rect 326 548 330 552
rect 198 538 202 542
rect 222 538 226 542
rect 158 488 162 492
rect 198 488 202 492
rect 222 488 226 492
rect 182 468 186 472
rect 70 348 74 352
rect 38 328 42 332
rect 294 498 298 502
rect 414 628 418 632
rect 438 628 442 632
rect 414 618 418 622
rect 470 618 474 622
rect 518 668 522 672
rect 534 668 538 672
rect 654 678 658 682
rect 702 678 706 682
rect 790 728 794 732
rect 870 728 874 732
rect 782 698 786 702
rect 858 703 862 707
rect 865 703 869 707
rect 926 718 930 722
rect 918 708 922 712
rect 806 698 810 702
rect 902 698 906 702
rect 566 668 570 672
rect 582 668 586 672
rect 526 658 530 662
rect 590 658 594 662
rect 494 638 498 642
rect 518 648 522 652
rect 526 648 530 652
rect 518 638 522 642
rect 550 638 554 642
rect 502 628 506 632
rect 934 708 938 712
rect 950 708 954 712
rect 926 688 930 692
rect 942 688 946 692
rect 870 678 874 682
rect 838 668 842 672
rect 822 658 826 662
rect 790 648 794 652
rect 646 638 650 642
rect 798 628 802 632
rect 702 618 706 622
rect 566 578 570 582
rect 678 578 682 582
rect 486 568 490 572
rect 518 568 522 572
rect 550 568 554 572
rect 630 568 634 572
rect 406 558 410 562
rect 462 558 466 562
rect 302 488 306 492
rect 390 488 394 492
rect 502 558 506 562
rect 494 548 498 552
rect 534 548 538 552
rect 630 548 634 552
rect 638 548 642 552
rect 518 538 522 542
rect 510 528 514 532
rect 558 528 562 532
rect 526 498 530 502
rect 310 468 314 472
rect 454 468 458 472
rect 206 458 210 462
rect 262 458 266 462
rect 278 458 282 462
rect 398 458 402 462
rect 558 458 562 462
rect 374 448 378 452
rect 406 448 410 452
rect 446 448 450 452
rect 470 448 474 452
rect 486 448 490 452
rect 310 438 314 442
rect 518 408 522 412
rect 346 403 350 407
rect 353 403 357 407
rect 342 358 346 362
rect 134 348 138 352
rect 198 348 202 352
rect 238 348 242 352
rect 310 348 314 352
rect 358 348 362 352
rect 398 348 402 352
rect 214 338 218 342
rect 246 338 250 342
rect 22 318 26 322
rect 78 318 82 322
rect 174 328 178 332
rect 78 298 82 302
rect 142 298 146 302
rect 46 268 50 272
rect 70 268 74 272
rect 110 258 114 262
rect 134 258 138 262
rect 38 248 42 252
rect 62 248 66 252
rect 86 248 90 252
rect 102 248 106 252
rect 142 248 146 252
rect 166 248 170 252
rect 46 228 50 232
rect 94 218 98 222
rect 22 198 26 202
rect 14 138 18 142
rect 494 347 498 351
rect 606 478 610 482
rect 622 458 626 462
rect 606 448 610 452
rect 574 368 578 372
rect 534 358 538 362
rect 566 358 570 362
rect 542 348 546 352
rect 646 458 650 462
rect 598 358 602 362
rect 622 358 626 362
rect 630 358 634 362
rect 582 348 586 352
rect 598 348 602 352
rect 358 338 362 342
rect 438 338 442 342
rect 446 338 450 342
rect 534 338 538 342
rect 558 338 562 342
rect 574 338 578 342
rect 598 338 602 342
rect 214 328 218 332
rect 254 328 258 332
rect 294 328 298 332
rect 230 308 234 312
rect 214 278 218 282
rect 230 268 234 272
rect 222 258 226 262
rect 270 278 274 282
rect 262 268 266 272
rect 310 328 314 332
rect 286 288 290 292
rect 430 308 434 312
rect 350 298 354 302
rect 414 288 418 292
rect 326 278 330 282
rect 350 278 354 282
rect 310 268 314 272
rect 246 258 250 262
rect 278 258 282 262
rect 302 258 306 262
rect 334 258 338 262
rect 414 268 418 272
rect 318 248 322 252
rect 190 238 194 242
rect 78 178 82 182
rect 150 228 154 232
rect 134 208 138 212
rect 86 168 90 172
rect 118 168 122 172
rect 126 158 130 162
rect 366 258 370 262
rect 398 248 402 252
rect 390 238 394 242
rect 310 218 314 222
rect 166 178 170 182
rect 214 208 218 212
rect 270 198 274 202
rect 238 188 242 192
rect 230 178 234 182
rect 158 158 162 162
rect 182 158 186 162
rect 190 158 194 162
rect 142 148 146 152
rect 54 138 58 142
rect 30 128 34 132
rect 126 118 130 122
rect 246 148 250 152
rect 254 148 258 152
rect 334 208 338 212
rect 318 178 322 182
rect 346 203 350 207
rect 353 203 357 207
rect 366 178 370 182
rect 390 168 394 172
rect 438 298 442 302
rect 478 278 482 282
rect 582 328 586 332
rect 686 538 690 542
rect 694 528 698 532
rect 766 608 770 612
rect 950 668 954 672
rect 862 658 866 662
rect 886 658 890 662
rect 846 628 850 632
rect 974 858 978 862
rect 990 858 994 862
rect 1038 938 1042 942
rect 1110 938 1114 942
rect 1142 938 1146 942
rect 1254 938 1258 942
rect 1270 938 1274 942
rect 1414 938 1418 942
rect 1438 938 1442 942
rect 1446 938 1450 942
rect 1078 928 1082 932
rect 1102 918 1106 922
rect 1094 898 1098 902
rect 1134 908 1138 912
rect 1134 898 1138 902
rect 1150 908 1154 912
rect 1166 908 1170 912
rect 1198 908 1202 912
rect 1150 898 1154 902
rect 1078 878 1082 882
rect 1134 878 1138 882
rect 1166 868 1170 872
rect 1038 858 1042 862
rect 1054 858 1058 862
rect 1022 848 1026 852
rect 1078 858 1082 862
rect 1046 848 1050 852
rect 1006 828 1010 832
rect 1006 808 1010 812
rect 1014 798 1018 802
rect 1054 768 1058 772
rect 1246 918 1250 922
rect 1238 908 1242 912
rect 1222 898 1226 902
rect 1214 878 1218 882
rect 1238 878 1242 882
rect 1238 868 1242 872
rect 1246 868 1250 872
rect 1158 858 1162 862
rect 1174 858 1178 862
rect 1198 858 1202 862
rect 1230 858 1234 862
rect 1094 848 1098 852
rect 1270 928 1274 932
rect 1278 908 1282 912
rect 1278 878 1282 882
rect 1262 868 1266 872
rect 1254 858 1258 862
rect 1326 908 1330 912
rect 1302 898 1306 902
rect 1302 878 1306 882
rect 1318 878 1322 882
rect 1478 1028 1482 1032
rect 1486 1028 1490 1032
rect 1526 1098 1530 1102
rect 1502 1078 1506 1082
rect 1510 1048 1514 1052
rect 1558 1098 1562 1102
rect 1550 1088 1554 1092
rect 1574 1068 1578 1072
rect 1550 1058 1554 1062
rect 1582 1058 1586 1062
rect 1814 1328 1818 1332
rect 1918 1328 1922 1332
rect 1926 1328 1930 1332
rect 1806 1318 1810 1322
rect 1894 1318 1898 1322
rect 1918 1318 1922 1322
rect 1874 1303 1878 1307
rect 1881 1303 1885 1307
rect 1846 1298 1850 1302
rect 1766 1278 1770 1282
rect 1790 1278 1794 1282
rect 1838 1278 1842 1282
rect 1750 1268 1754 1272
rect 1774 1268 1778 1272
rect 1710 1258 1714 1262
rect 1758 1258 1762 1262
rect 1782 1258 1786 1262
rect 2030 1358 2034 1362
rect 2118 1468 2122 1472
rect 2134 1468 2138 1472
rect 2166 1468 2170 1472
rect 2134 1438 2138 1442
rect 2302 1708 2306 1712
rect 2342 1728 2346 1732
rect 2382 1728 2386 1732
rect 2358 1718 2362 1722
rect 2366 1718 2370 1722
rect 2310 1698 2314 1702
rect 2294 1688 2298 1692
rect 2422 1748 2426 1752
rect 2502 1858 2506 1862
rect 2534 1858 2538 1862
rect 2566 1858 2570 1862
rect 2574 1858 2578 1862
rect 2646 1948 2650 1952
rect 2726 2098 2730 2102
rect 2894 2158 2898 2162
rect 2942 2198 2946 2202
rect 3078 2338 3082 2342
rect 3102 2338 3106 2342
rect 3054 2328 3058 2332
rect 3262 2378 3266 2382
rect 3358 2378 3362 2382
rect 3198 2368 3202 2372
rect 3230 2368 3234 2372
rect 3254 2368 3258 2372
rect 3206 2358 3210 2362
rect 3278 2368 3282 2372
rect 3326 2368 3330 2372
rect 3318 2358 3322 2362
rect 3350 2358 3354 2362
rect 3366 2358 3370 2362
rect 3166 2348 3170 2352
rect 3270 2348 3274 2352
rect 3318 2348 3322 2352
rect 3366 2348 3370 2352
rect 3382 2358 3386 2362
rect 3406 2498 3410 2502
rect 3406 2478 3410 2482
rect 3454 2528 3458 2532
rect 3470 2508 3474 2512
rect 3654 2718 3658 2722
rect 3694 2758 3698 2762
rect 3710 2758 3714 2762
rect 3702 2748 3706 2752
rect 3662 2708 3666 2712
rect 3646 2678 3650 2682
rect 4214 2948 4218 2952
rect 4246 2948 4250 2952
rect 4046 2938 4050 2942
rect 4078 2938 4082 2942
rect 3974 2918 3978 2922
rect 4070 2928 4074 2932
rect 4038 2908 4042 2912
rect 4078 2918 4082 2922
rect 4054 2908 4058 2912
rect 4046 2888 4050 2892
rect 3966 2878 3970 2882
rect 4014 2878 4018 2882
rect 4142 2908 4146 2912
rect 4086 2888 4090 2892
rect 4094 2888 4098 2892
rect 4118 2888 4122 2892
rect 3990 2868 3994 2872
rect 3958 2858 3962 2862
rect 3974 2858 3978 2862
rect 3918 2838 3922 2842
rect 3942 2838 3946 2842
rect 3974 2838 3978 2842
rect 4038 2858 4042 2862
rect 3998 2838 4002 2842
rect 3990 2828 3994 2832
rect 4022 2838 4026 2842
rect 4046 2838 4050 2842
rect 4014 2828 4018 2832
rect 4030 2828 4034 2832
rect 3998 2818 4002 2822
rect 4014 2818 4018 2822
rect 3950 2808 3954 2812
rect 3798 2778 3802 2782
rect 3886 2768 3890 2772
rect 3782 2758 3786 2762
rect 3854 2758 3858 2762
rect 3742 2748 3746 2752
rect 3814 2748 3818 2752
rect 3846 2748 3850 2752
rect 3798 2738 3802 2742
rect 3822 2738 3826 2742
rect 3846 2738 3850 2742
rect 3854 2738 3858 2742
rect 3686 2728 3690 2732
rect 3718 2728 3722 2732
rect 3750 2728 3754 2732
rect 3678 2708 3682 2712
rect 3782 2718 3786 2722
rect 3814 2728 3818 2732
rect 3726 2708 3730 2712
rect 3806 2698 3810 2702
rect 3782 2678 3786 2682
rect 3702 2668 3706 2672
rect 3646 2648 3650 2652
rect 3654 2648 3658 2652
rect 3678 2648 3682 2652
rect 3630 2618 3634 2622
rect 3606 2598 3610 2602
rect 3718 2648 3722 2652
rect 3710 2588 3714 2592
rect 3574 2558 3578 2562
rect 3670 2558 3674 2562
rect 3894 2748 3898 2752
rect 3942 2738 3946 2742
rect 3870 2728 3874 2732
rect 3930 2703 3934 2707
rect 3937 2703 3941 2707
rect 3878 2698 3882 2702
rect 3822 2668 3826 2672
rect 3830 2668 3834 2672
rect 4110 2868 4114 2872
rect 4110 2848 4114 2852
rect 4142 2878 4146 2882
rect 4134 2858 4138 2862
rect 4302 2998 4306 3002
rect 4318 2998 4322 3002
rect 4342 3048 4346 3052
rect 4414 3048 4418 3052
rect 4430 3048 4434 3052
rect 4382 3038 4386 3042
rect 4350 2948 4354 2952
rect 4326 2938 4330 2942
rect 4206 2918 4210 2922
rect 4150 2868 4154 2872
rect 4174 2858 4178 2862
rect 4030 2808 4034 2812
rect 4038 2808 4042 2812
rect 4078 2808 4082 2812
rect 4094 2788 4098 2792
rect 4142 2848 4146 2852
rect 4166 2848 4170 2852
rect 4198 2848 4202 2852
rect 4190 2818 4194 2822
rect 4046 2778 4050 2782
rect 4134 2778 4138 2782
rect 3974 2768 3978 2772
rect 4022 2768 4026 2772
rect 4062 2768 4066 2772
rect 3966 2758 3970 2762
rect 3998 2758 4002 2762
rect 4094 2758 4098 2762
rect 3982 2748 3986 2752
rect 4046 2748 4050 2752
rect 4094 2748 4098 2752
rect 4414 2928 4418 2932
rect 4230 2888 4234 2892
rect 4214 2868 4218 2872
rect 4278 2868 4282 2872
rect 4286 2848 4290 2852
rect 4270 2818 4274 2822
rect 4310 2808 4314 2812
rect 4358 2859 4362 2862
rect 4358 2858 4362 2859
rect 4358 2798 4362 2802
rect 4590 3058 4594 3062
rect 4542 3048 4546 3052
rect 4478 3038 4482 3042
rect 4494 3038 4498 3042
rect 4442 3003 4446 3007
rect 4449 3003 4453 3007
rect 4510 2968 4514 2972
rect 4542 2968 4546 2972
rect 4446 2958 4450 2962
rect 4518 2958 4522 2962
rect 4470 2948 4474 2952
rect 4494 2948 4498 2952
rect 4462 2938 4466 2942
rect 4526 2938 4530 2942
rect 4470 2928 4474 2932
rect 4438 2918 4442 2922
rect 4574 2958 4578 2962
rect 4558 2938 4562 2942
rect 4558 2928 4562 2932
rect 4502 2918 4506 2922
rect 4542 2888 4546 2892
rect 4494 2878 4498 2882
rect 4606 2918 4610 2922
rect 4598 2878 4602 2882
rect 4590 2868 4594 2872
rect 4494 2828 4498 2832
rect 4442 2803 4446 2807
rect 4449 2803 4453 2807
rect 4750 3128 4754 3132
rect 4686 3098 4690 3102
rect 4718 3068 4722 3072
rect 4846 3068 4850 3072
rect 4734 3058 4738 3062
rect 4862 3058 4866 3062
rect 5014 3238 5018 3242
rect 5086 3258 5090 3262
rect 5134 3268 5138 3272
rect 5214 3268 5218 3272
rect 5110 3258 5114 3262
rect 5166 3258 5170 3262
rect 5070 3238 5074 3242
rect 5094 3238 5098 3242
rect 4998 3228 5002 3232
rect 5062 3228 5066 3232
rect 4982 3178 4986 3182
rect 4918 3158 4922 3162
rect 4934 3148 4938 3152
rect 4918 3138 4922 3142
rect 4942 3138 4946 3142
rect 4950 3128 4954 3132
rect 4942 3118 4946 3122
rect 4974 3118 4978 3122
rect 4954 3103 4958 3107
rect 4961 3103 4965 3107
rect 4958 3088 4962 3092
rect 4950 3078 4954 3082
rect 4942 3058 4946 3062
rect 4750 3048 4754 3052
rect 4822 3048 4826 3052
rect 4830 3048 4834 3052
rect 4934 3048 4938 3052
rect 4854 2988 4858 2992
rect 4782 2958 4786 2962
rect 4702 2948 4706 2952
rect 4742 2948 4746 2952
rect 4766 2928 4770 2932
rect 4638 2918 4642 2922
rect 4670 2888 4674 2892
rect 4750 2888 4754 2892
rect 4614 2878 4618 2882
rect 4638 2858 4642 2862
rect 4574 2848 4578 2852
rect 4622 2848 4626 2852
rect 4694 2868 4698 2872
rect 4726 2868 4730 2872
rect 4854 2878 4858 2882
rect 4790 2868 4794 2872
rect 4830 2868 4834 2872
rect 4686 2858 4690 2862
rect 4718 2858 4722 2862
rect 4774 2858 4778 2862
rect 4886 2878 4890 2882
rect 4958 2938 4962 2942
rect 4982 3068 4986 3072
rect 5094 3178 5098 3182
rect 5030 3168 5034 3172
rect 5070 3168 5074 3172
rect 5022 3128 5026 3132
rect 5038 3118 5042 3122
rect 5006 3088 5010 3092
rect 5078 3158 5082 3162
rect 5086 3078 5090 3082
rect 5030 3068 5034 3072
rect 5022 3058 5026 3062
rect 5030 3048 5034 3052
rect 5086 3048 5090 3052
rect 4998 2988 5002 2992
rect 5030 2988 5034 2992
rect 5054 2978 5058 2982
rect 5262 3288 5266 3292
rect 5214 3258 5218 3262
rect 5198 3248 5202 3252
rect 5270 3248 5274 3252
rect 5118 3228 5122 3232
rect 5294 3258 5298 3262
rect 5286 3228 5290 3232
rect 5270 3188 5274 3192
rect 5246 3178 5250 3182
rect 5198 3158 5202 3162
rect 5214 3148 5218 3152
rect 5278 3178 5282 3182
rect 5286 3158 5290 3162
rect 5126 3138 5130 3142
rect 5118 3118 5122 3122
rect 4982 2948 4986 2952
rect 5054 2948 5058 2952
rect 5078 2948 5082 2952
rect 5102 2948 5106 2952
rect 5006 2938 5010 2942
rect 4958 2918 4962 2922
rect 4954 2903 4958 2907
rect 4961 2903 4965 2907
rect 5142 3118 5146 3122
rect 5142 3088 5146 3092
rect 5246 3138 5250 3142
rect 5262 3138 5266 3142
rect 5254 3088 5258 3092
rect 5246 3078 5250 3082
rect 5134 2988 5138 2992
rect 5198 2958 5202 2962
rect 5142 2948 5146 2952
rect 5166 2948 5170 2952
rect 5110 2928 5114 2932
rect 5078 2898 5082 2902
rect 5038 2888 5042 2892
rect 4910 2878 4914 2882
rect 4942 2878 4946 2882
rect 4990 2878 4994 2882
rect 5014 2878 5018 2882
rect 4918 2868 4922 2872
rect 4982 2868 4986 2872
rect 4870 2858 4874 2862
rect 4902 2858 4906 2862
rect 4934 2858 4938 2862
rect 4814 2848 4818 2852
rect 4582 2838 4586 2842
rect 4598 2838 4602 2842
rect 4646 2838 4650 2842
rect 4566 2828 4570 2832
rect 4430 2788 4434 2792
rect 4518 2788 4522 2792
rect 4390 2778 4394 2782
rect 4398 2768 4402 2772
rect 4414 2768 4418 2772
rect 4598 2768 4602 2772
rect 4630 2768 4634 2772
rect 4358 2758 4362 2762
rect 4430 2758 4434 2762
rect 4454 2758 4458 2762
rect 4502 2758 4506 2762
rect 4526 2758 4530 2762
rect 4278 2748 4282 2752
rect 4054 2738 4058 2742
rect 3862 2658 3866 2662
rect 3918 2658 3922 2662
rect 4102 2738 4106 2742
rect 4134 2738 4138 2742
rect 4086 2678 4090 2682
rect 3838 2648 3842 2652
rect 3926 2648 3930 2652
rect 3854 2638 3858 2642
rect 3902 2638 3906 2642
rect 4094 2658 4098 2662
rect 4070 2648 4074 2652
rect 4014 2638 4018 2642
rect 3982 2628 3986 2632
rect 3958 2588 3962 2592
rect 3838 2578 3842 2582
rect 3646 2547 3650 2551
rect 3726 2548 3730 2552
rect 3662 2538 3666 2542
rect 3462 2498 3466 2502
rect 3478 2498 3482 2502
rect 3446 2478 3450 2482
rect 3486 2468 3490 2472
rect 3526 2458 3530 2462
rect 3534 2458 3538 2462
rect 3494 2448 3498 2452
rect 3542 2448 3546 2452
rect 3598 2478 3602 2482
rect 3630 2478 3634 2482
rect 3566 2468 3570 2472
rect 3606 2458 3610 2462
rect 3630 2458 3634 2462
rect 3646 2458 3650 2462
rect 3582 2448 3586 2452
rect 3638 2448 3642 2452
rect 3742 2528 3746 2532
rect 3870 2568 3874 2572
rect 3862 2558 3866 2562
rect 3782 2518 3786 2522
rect 3822 2518 3826 2522
rect 3686 2478 3690 2482
rect 3734 2478 3738 2482
rect 3670 2468 3674 2472
rect 3822 2478 3826 2482
rect 3798 2468 3802 2472
rect 3758 2458 3762 2462
rect 3718 2448 3722 2452
rect 3502 2438 3506 2442
rect 3526 2438 3530 2442
rect 3558 2438 3562 2442
rect 3406 2428 3410 2432
rect 3398 2348 3402 2352
rect 3190 2338 3194 2342
rect 3278 2338 3282 2342
rect 3310 2338 3314 2342
rect 3358 2338 3362 2342
rect 3374 2338 3378 2342
rect 3150 2328 3154 2332
rect 3158 2328 3162 2332
rect 3182 2328 3186 2332
rect 3246 2328 3250 2332
rect 3294 2328 3298 2332
rect 3310 2328 3314 2332
rect 3070 2318 3074 2322
rect 3118 2318 3122 2322
rect 3006 2308 3010 2312
rect 3006 2288 3010 2292
rect 3086 2288 3090 2292
rect 3070 2278 3074 2282
rect 3062 2268 3066 2272
rect 3014 2248 3018 2252
rect 3206 2318 3210 2322
rect 3214 2318 3218 2322
rect 3142 2308 3146 2312
rect 3142 2288 3146 2292
rect 3102 2268 3106 2272
rect 3134 2268 3138 2272
rect 3102 2258 3106 2262
rect 3134 2258 3138 2262
rect 3166 2278 3170 2282
rect 3222 2288 3226 2292
rect 3278 2268 3282 2272
rect 3294 2268 3298 2272
rect 3382 2328 3386 2332
rect 3382 2318 3386 2322
rect 3638 2428 3642 2432
rect 3526 2418 3530 2422
rect 3418 2403 3422 2407
rect 3425 2403 3429 2407
rect 3454 2398 3458 2402
rect 3582 2388 3586 2392
rect 3478 2368 3482 2372
rect 3518 2368 3522 2372
rect 3494 2358 3498 2362
rect 3494 2348 3498 2352
rect 3414 2338 3418 2342
rect 3470 2328 3474 2332
rect 3526 2348 3530 2352
rect 3622 2358 3626 2362
rect 3590 2348 3594 2352
rect 3614 2348 3618 2352
rect 3646 2348 3650 2352
rect 3518 2338 3522 2342
rect 3526 2338 3530 2342
rect 3510 2318 3514 2322
rect 3614 2318 3618 2322
rect 3366 2288 3370 2292
rect 3526 2308 3530 2312
rect 3550 2298 3554 2302
rect 3638 2298 3642 2302
rect 3558 2288 3562 2292
rect 3422 2278 3426 2282
rect 3478 2278 3482 2282
rect 3582 2278 3586 2282
rect 3590 2278 3594 2282
rect 3374 2268 3378 2272
rect 3390 2268 3394 2272
rect 3286 2248 3290 2252
rect 3326 2248 3330 2252
rect 3366 2248 3370 2252
rect 3382 2238 3386 2242
rect 3334 2228 3338 2232
rect 3190 2218 3194 2222
rect 3246 2208 3250 2212
rect 3142 2198 3146 2202
rect 3046 2178 3050 2182
rect 3070 2158 3074 2162
rect 2894 2148 2898 2152
rect 2926 2148 2930 2152
rect 3046 2148 3050 2152
rect 3190 2158 3194 2162
rect 3198 2158 3202 2162
rect 3214 2158 3218 2162
rect 3230 2158 3234 2162
rect 3062 2148 3066 2152
rect 3078 2148 3082 2152
rect 3134 2148 3138 2152
rect 3054 2138 3058 2142
rect 2926 2128 2930 2132
rect 2974 2128 2978 2132
rect 2982 2128 2986 2132
rect 2906 2103 2910 2107
rect 2913 2103 2917 2107
rect 3094 2138 3098 2142
rect 3118 2138 3122 2142
rect 3158 2138 3162 2142
rect 3214 2148 3218 2152
rect 3230 2148 3234 2152
rect 3254 2158 3258 2162
rect 3262 2148 3266 2152
rect 3278 2148 3282 2152
rect 3366 2198 3370 2202
rect 3478 2258 3482 2262
rect 3398 2218 3402 2222
rect 3478 2218 3482 2222
rect 3418 2203 3422 2207
rect 3425 2203 3429 2207
rect 3406 2198 3410 2202
rect 3302 2148 3306 2152
rect 3318 2148 3322 2152
rect 3334 2148 3338 2152
rect 3390 2148 3394 2152
rect 3406 2148 3410 2152
rect 3238 2138 3242 2142
rect 3270 2138 3274 2142
rect 3286 2138 3290 2142
rect 3294 2138 3298 2142
rect 3070 2128 3074 2132
rect 3142 2128 3146 2132
rect 3078 2108 3082 2112
rect 3054 2088 3058 2092
rect 2854 2078 2858 2082
rect 2870 2078 2874 2082
rect 2926 2078 2930 2082
rect 3006 2078 3010 2082
rect 3046 2078 3050 2082
rect 2742 2068 2746 2072
rect 2774 2068 2778 2072
rect 2790 2068 2794 2072
rect 2822 2068 2826 2072
rect 2766 2058 2770 2062
rect 2798 2058 2802 2062
rect 2830 2058 2834 2062
rect 2726 2048 2730 2052
rect 2766 2048 2770 2052
rect 2982 2068 2986 2072
rect 2798 2048 2802 2052
rect 2838 2048 2842 2052
rect 2782 2038 2786 2042
rect 2726 1998 2730 2002
rect 2838 1998 2842 2002
rect 2782 1948 2786 1952
rect 2806 1948 2810 1952
rect 2830 1948 2834 1952
rect 2838 1948 2842 1952
rect 2614 1918 2618 1922
rect 2606 1878 2610 1882
rect 2590 1858 2594 1862
rect 2510 1848 2514 1852
rect 2526 1838 2530 1842
rect 2558 1838 2562 1842
rect 2566 1838 2570 1842
rect 2534 1818 2538 1822
rect 2470 1808 2474 1812
rect 2438 1768 2442 1772
rect 2446 1768 2450 1772
rect 2462 1768 2466 1772
rect 2550 1768 2554 1772
rect 2518 1758 2522 1762
rect 2462 1748 2466 1752
rect 2478 1748 2482 1752
rect 2502 1748 2506 1752
rect 2430 1738 2434 1742
rect 2438 1738 2442 1742
rect 2486 1738 2490 1742
rect 2510 1738 2514 1742
rect 2582 1768 2586 1772
rect 2566 1758 2570 1762
rect 2606 1818 2610 1822
rect 2630 1898 2634 1902
rect 2734 1908 2738 1912
rect 2662 1898 2666 1902
rect 2694 1898 2698 1902
rect 2718 1898 2722 1902
rect 2726 1898 2730 1902
rect 2638 1888 2642 1892
rect 2694 1878 2698 1882
rect 2718 1878 2722 1882
rect 2622 1868 2626 1872
rect 2654 1868 2658 1872
rect 2670 1868 2674 1872
rect 2702 1866 2706 1870
rect 2670 1858 2674 1862
rect 2630 1848 2634 1852
rect 2646 1848 2650 1852
rect 2814 1938 2818 1942
rect 2798 1928 2802 1932
rect 2822 1928 2826 1932
rect 2830 1918 2834 1922
rect 2798 1908 2802 1912
rect 2806 1908 2810 1912
rect 2766 1898 2770 1902
rect 2758 1888 2762 1892
rect 2814 1898 2818 1902
rect 2734 1858 2738 1862
rect 2750 1848 2754 1852
rect 2686 1838 2690 1842
rect 2774 1858 2778 1862
rect 2774 1848 2778 1852
rect 2782 1848 2786 1852
rect 2638 1818 2642 1822
rect 2638 1758 2642 1762
rect 2646 1758 2650 1762
rect 2542 1748 2546 1752
rect 2550 1748 2554 1752
rect 2574 1748 2578 1752
rect 2598 1748 2602 1752
rect 2606 1748 2610 1752
rect 2670 1748 2674 1752
rect 2542 1738 2546 1742
rect 2534 1728 2538 1732
rect 2558 1728 2562 1732
rect 2462 1708 2466 1712
rect 2446 1698 2450 1702
rect 2582 1738 2586 1742
rect 2646 1738 2650 1742
rect 2718 1828 2722 1832
rect 2726 1738 2730 1742
rect 2662 1728 2666 1732
rect 2566 1718 2570 1722
rect 2574 1698 2578 1702
rect 2598 1688 2602 1692
rect 2414 1678 2418 1682
rect 2510 1678 2514 1682
rect 2534 1678 2538 1682
rect 2558 1678 2562 1682
rect 2646 1678 2650 1682
rect 2694 1728 2698 1732
rect 2702 1728 2706 1732
rect 2734 1728 2738 1732
rect 2742 1718 2746 1722
rect 2350 1668 2354 1672
rect 2366 1668 2370 1672
rect 2374 1668 2378 1672
rect 2454 1668 2458 1672
rect 2478 1668 2482 1672
rect 2518 1668 2522 1672
rect 2326 1658 2330 1662
rect 2270 1648 2274 1652
rect 2310 1648 2314 1652
rect 2342 1648 2346 1652
rect 2366 1648 2370 1652
rect 2390 1648 2394 1652
rect 2246 1608 2250 1612
rect 2262 1588 2266 1592
rect 2350 1608 2354 1612
rect 2318 1588 2322 1592
rect 2246 1578 2250 1582
rect 2294 1578 2298 1582
rect 2222 1548 2226 1552
rect 2294 1568 2298 1572
rect 2406 1648 2410 1652
rect 2462 1648 2466 1652
rect 2470 1648 2474 1652
rect 2398 1618 2402 1622
rect 2394 1603 2398 1607
rect 2401 1603 2405 1607
rect 2382 1598 2386 1602
rect 2278 1558 2282 1562
rect 2326 1558 2330 1562
rect 2294 1548 2298 1552
rect 2366 1548 2370 1552
rect 2238 1528 2242 1532
rect 2278 1498 2282 1502
rect 2342 1528 2346 1532
rect 2318 1508 2322 1512
rect 2406 1578 2410 1582
rect 2414 1568 2418 1572
rect 2446 1548 2450 1552
rect 2574 1658 2578 1662
rect 2614 1658 2618 1662
rect 2702 1658 2706 1662
rect 2518 1648 2522 1652
rect 2590 1648 2594 1652
rect 2622 1648 2626 1652
rect 2646 1648 2650 1652
rect 2542 1628 2546 1632
rect 2502 1568 2506 1572
rect 2478 1508 2482 1512
rect 2382 1498 2386 1502
rect 2742 1638 2746 1642
rect 2694 1608 2698 1612
rect 2630 1588 2634 1592
rect 2742 1568 2746 1572
rect 2590 1558 2594 1562
rect 2582 1538 2586 1542
rect 2574 1518 2578 1522
rect 2518 1498 2522 1502
rect 2534 1498 2538 1502
rect 2270 1478 2274 1482
rect 2278 1478 2282 1482
rect 2302 1478 2306 1482
rect 2366 1478 2370 1482
rect 2494 1478 2498 1482
rect 2510 1478 2514 1482
rect 2478 1468 2482 1472
rect 2494 1468 2498 1472
rect 2198 1458 2202 1462
rect 2222 1459 2226 1463
rect 2278 1458 2282 1462
rect 2182 1448 2186 1452
rect 2150 1428 2154 1432
rect 2174 1428 2178 1432
rect 2174 1408 2178 1412
rect 2142 1398 2146 1402
rect 2078 1378 2082 1382
rect 2110 1378 2114 1382
rect 2118 1358 2122 1362
rect 2014 1348 2018 1352
rect 1966 1318 1970 1322
rect 1958 1308 1962 1312
rect 2222 1398 2226 1402
rect 2310 1448 2314 1452
rect 2334 1448 2338 1452
rect 2286 1438 2290 1442
rect 2302 1438 2306 1442
rect 2486 1458 2490 1462
rect 2494 1458 2498 1462
rect 3174 2098 3178 2102
rect 3102 2078 3106 2082
rect 3134 2078 3138 2082
rect 3198 2078 3202 2082
rect 3078 2068 3082 2072
rect 3094 2068 3098 2072
rect 3158 2068 3162 2072
rect 2894 2038 2898 2042
rect 2942 2018 2946 2022
rect 2926 2008 2930 2012
rect 2886 1948 2890 1952
rect 2878 1938 2882 1942
rect 2854 1928 2858 1932
rect 2862 1918 2866 1922
rect 2846 1898 2850 1902
rect 2830 1868 2834 1872
rect 2846 1868 2850 1872
rect 2870 1868 2874 1872
rect 2822 1858 2826 1862
rect 2798 1748 2802 1752
rect 2822 1748 2826 1752
rect 2854 1858 2858 1862
rect 2870 1848 2874 1852
rect 2906 1903 2910 1907
rect 2913 1903 2917 1907
rect 2990 1948 2994 1952
rect 3070 2058 3074 2062
rect 3078 2058 3082 2062
rect 3054 2018 3058 2022
rect 3022 1938 3026 1942
rect 2942 1928 2946 1932
rect 2934 1918 2938 1922
rect 2998 1918 3002 1922
rect 2958 1908 2962 1912
rect 2958 1898 2962 1902
rect 2910 1868 2914 1872
rect 2918 1868 2922 1872
rect 2894 1858 2898 1862
rect 2902 1858 2906 1862
rect 2918 1858 2922 1862
rect 2878 1838 2882 1842
rect 2854 1818 2858 1822
rect 2870 1818 2874 1822
rect 2894 1758 2898 1762
rect 2862 1748 2866 1752
rect 2854 1738 2858 1742
rect 2870 1738 2874 1742
rect 2766 1718 2770 1722
rect 2958 1868 2962 1872
rect 2990 1868 2994 1872
rect 2934 1858 2938 1862
rect 2966 1858 2970 1862
rect 3022 1818 3026 1822
rect 3078 1998 3082 2002
rect 3102 2058 3106 2062
rect 3134 2058 3138 2062
rect 3230 2068 3234 2072
rect 3190 2058 3194 2062
rect 3214 2058 3218 2062
rect 3134 2048 3138 2052
rect 3174 2048 3178 2052
rect 3182 2048 3186 2052
rect 3110 2028 3114 2032
rect 3150 2028 3154 2032
rect 3102 1998 3106 2002
rect 3158 1998 3162 2002
rect 3118 1948 3122 1952
rect 3086 1928 3090 1932
rect 3062 1858 3066 1862
rect 2990 1768 2994 1772
rect 2934 1758 2938 1762
rect 2958 1758 2962 1762
rect 2982 1758 2986 1762
rect 2990 1758 2994 1762
rect 2934 1748 2938 1752
rect 2926 1728 2930 1732
rect 2942 1728 2946 1732
rect 2798 1718 2802 1722
rect 2774 1708 2778 1712
rect 2846 1708 2850 1712
rect 2814 1688 2818 1692
rect 2906 1703 2910 1707
rect 2913 1703 2917 1707
rect 2966 1748 2970 1752
rect 3014 1748 3018 1752
rect 3006 1738 3010 1742
rect 2982 1718 2986 1722
rect 2974 1698 2978 1702
rect 2958 1688 2962 1692
rect 2774 1668 2778 1672
rect 2942 1668 2946 1672
rect 2758 1658 2762 1662
rect 2814 1658 2818 1662
rect 3030 1768 3034 1772
rect 3046 1748 3050 1752
rect 3038 1738 3042 1742
rect 3118 1888 3122 1892
rect 3142 1948 3146 1952
rect 3142 1928 3146 1932
rect 3110 1868 3114 1872
rect 3126 1868 3130 1872
rect 3174 1938 3178 1942
rect 3326 2098 3330 2102
rect 3254 2078 3258 2082
rect 3318 2068 3322 2072
rect 3286 2058 3290 2062
rect 3206 2048 3210 2052
rect 3294 2048 3298 2052
rect 3350 2098 3354 2102
rect 3358 2078 3362 2082
rect 3566 2248 3570 2252
rect 3494 2208 3498 2212
rect 3622 2228 3626 2232
rect 3614 2198 3618 2202
rect 3566 2168 3570 2172
rect 3606 2148 3610 2152
rect 3726 2438 3730 2442
rect 3726 2408 3730 2412
rect 3694 2378 3698 2382
rect 3742 2428 3746 2432
rect 3734 2388 3738 2392
rect 3806 2448 3810 2452
rect 3806 2428 3810 2432
rect 3942 2558 3946 2562
rect 3886 2548 3890 2552
rect 3910 2548 3914 2552
rect 3878 2528 3882 2532
rect 3910 2528 3914 2532
rect 3982 2578 3986 2582
rect 4070 2598 4074 2602
rect 4142 2668 4146 2672
rect 4158 2668 4162 2672
rect 4126 2658 4130 2662
rect 4166 2658 4170 2662
rect 4118 2648 4122 2652
rect 4302 2747 4306 2751
rect 4510 2748 4514 2752
rect 4230 2738 4234 2742
rect 4382 2738 4386 2742
rect 4270 2718 4274 2722
rect 4374 2718 4378 2722
rect 4206 2688 4210 2692
rect 4190 2678 4194 2682
rect 4230 2678 4234 2682
rect 4238 2678 4242 2682
rect 4286 2678 4290 2682
rect 4174 2638 4178 2642
rect 4182 2588 4186 2592
rect 4102 2568 4106 2572
rect 3982 2558 3986 2562
rect 3990 2558 3994 2562
rect 4014 2558 4018 2562
rect 4022 2558 4026 2562
rect 4046 2558 4050 2562
rect 3974 2528 3978 2532
rect 3958 2518 3962 2522
rect 3930 2503 3934 2507
rect 3937 2503 3941 2507
rect 3902 2488 3906 2492
rect 3878 2478 3882 2482
rect 3854 2458 3858 2462
rect 3870 2458 3874 2462
rect 3894 2458 3898 2462
rect 3918 2458 3922 2462
rect 3934 2458 3938 2462
rect 3886 2448 3890 2452
rect 3910 2448 3914 2452
rect 4014 2548 4018 2552
rect 3982 2518 3986 2522
rect 3982 2508 3986 2512
rect 4054 2548 4058 2552
rect 4134 2547 4138 2551
rect 4030 2518 4034 2522
rect 4038 2518 4042 2522
rect 4062 2518 4066 2522
rect 3990 2498 3994 2502
rect 3998 2488 4002 2492
rect 3974 2468 3978 2472
rect 4014 2488 4018 2492
rect 4014 2478 4018 2482
rect 4062 2498 4066 2502
rect 4046 2468 4050 2472
rect 3950 2458 3954 2462
rect 4030 2458 4034 2462
rect 4046 2458 4050 2462
rect 3998 2448 4002 2452
rect 3942 2438 3946 2442
rect 4006 2438 4010 2442
rect 4086 2518 4090 2522
rect 4462 2738 4466 2742
rect 4494 2738 4498 2742
rect 4382 2678 4386 2682
rect 4262 2668 4266 2672
rect 4350 2668 4354 2672
rect 4302 2658 4306 2662
rect 4334 2658 4338 2662
rect 4534 2748 4538 2752
rect 4574 2738 4578 2742
rect 4742 2838 4746 2842
rect 4710 2828 4714 2832
rect 4694 2778 4698 2782
rect 4718 2778 4722 2782
rect 4678 2768 4682 2772
rect 4710 2768 4714 2772
rect 4758 2828 4762 2832
rect 4726 2758 4730 2762
rect 4742 2758 4746 2762
rect 4662 2748 4666 2752
rect 4694 2748 4698 2752
rect 4734 2748 4738 2752
rect 4622 2738 4626 2742
rect 4878 2768 4882 2772
rect 4862 2758 4866 2762
rect 4798 2748 4802 2752
rect 4846 2748 4850 2752
rect 4798 2738 4802 2742
rect 4806 2738 4810 2742
rect 4822 2738 4826 2742
rect 4486 2728 4490 2732
rect 4542 2728 4546 2732
rect 4614 2728 4618 2732
rect 4638 2728 4642 2732
rect 4894 2758 4898 2762
rect 4926 2748 4930 2752
rect 4894 2738 4898 2742
rect 4926 2738 4930 2742
rect 4750 2728 4754 2732
rect 4822 2728 4826 2732
rect 4894 2728 4898 2732
rect 4646 2718 4650 2722
rect 4686 2718 4690 2722
rect 4758 2718 4762 2722
rect 4790 2718 4794 2722
rect 4622 2688 4626 2692
rect 4670 2698 4674 2702
rect 4598 2678 4602 2682
rect 4638 2678 4642 2682
rect 4590 2668 4594 2672
rect 4622 2668 4626 2672
rect 4646 2668 4650 2672
rect 4510 2658 4514 2662
rect 4222 2648 4226 2652
rect 4238 2648 4242 2652
rect 4262 2648 4266 2652
rect 4278 2648 4282 2652
rect 4326 2648 4330 2652
rect 4358 2648 4362 2652
rect 4214 2638 4218 2642
rect 4254 2638 4258 2642
rect 4198 2628 4202 2632
rect 4198 2538 4202 2542
rect 4190 2528 4194 2532
rect 4158 2518 4162 2522
rect 4190 2508 4194 2512
rect 4342 2638 4346 2642
rect 4542 2658 4546 2662
rect 4686 2658 4690 2662
rect 4574 2648 4578 2652
rect 4606 2648 4610 2652
rect 4750 2698 4754 2702
rect 4782 2698 4786 2702
rect 4790 2688 4794 2692
rect 4726 2678 4730 2682
rect 4718 2668 4722 2672
rect 4734 2668 4738 2672
rect 4814 2718 4818 2722
rect 4870 2718 4874 2722
rect 4822 2708 4826 2712
rect 4846 2698 4850 2702
rect 4814 2688 4818 2692
rect 4822 2678 4826 2682
rect 4702 2648 4706 2652
rect 4926 2718 4930 2722
rect 4854 2678 4858 2682
rect 4878 2678 4882 2682
rect 4862 2648 4866 2652
rect 4710 2638 4714 2642
rect 4734 2638 4738 2642
rect 4534 2628 4538 2632
rect 4646 2628 4650 2632
rect 4678 2628 4682 2632
rect 4334 2618 4338 2622
rect 4414 2618 4418 2622
rect 4462 2618 4466 2622
rect 4638 2618 4642 2622
rect 4534 2608 4538 2612
rect 4442 2603 4446 2607
rect 4449 2603 4453 2607
rect 4478 2578 4482 2582
rect 4390 2568 4394 2572
rect 4422 2568 4426 2572
rect 4462 2568 4466 2572
rect 4502 2568 4506 2572
rect 4622 2568 4626 2572
rect 4422 2558 4426 2562
rect 4494 2558 4498 2562
rect 4558 2558 4562 2562
rect 4590 2558 4594 2562
rect 4366 2548 4370 2552
rect 4406 2548 4410 2552
rect 4350 2538 4354 2542
rect 4382 2538 4386 2542
rect 4398 2538 4402 2542
rect 4422 2538 4426 2542
rect 4478 2538 4482 2542
rect 4246 2528 4250 2532
rect 4246 2518 4250 2522
rect 4238 2488 4242 2492
rect 4230 2478 4234 2482
rect 4270 2478 4274 2482
rect 4190 2468 4194 2472
rect 4222 2468 4226 2472
rect 4238 2468 4242 2472
rect 4246 2468 4250 2472
rect 4094 2458 4098 2462
rect 4086 2448 4090 2452
rect 4070 2438 4074 2442
rect 3798 2388 3802 2392
rect 3830 2388 3834 2392
rect 3766 2378 3770 2382
rect 3758 2368 3762 2372
rect 3750 2358 3754 2362
rect 3774 2358 3778 2362
rect 3782 2358 3786 2362
rect 3678 2348 3682 2352
rect 3830 2378 3834 2382
rect 3822 2358 3826 2362
rect 3662 2338 3666 2342
rect 3710 2338 3714 2342
rect 3758 2338 3762 2342
rect 3790 2338 3794 2342
rect 3678 2328 3682 2332
rect 3670 2278 3674 2282
rect 3726 2308 3730 2312
rect 3662 2258 3666 2262
rect 3870 2348 3874 2352
rect 3854 2338 3858 2342
rect 3934 2408 3938 2412
rect 3974 2408 3978 2412
rect 3942 2378 3946 2382
rect 3950 2378 3954 2382
rect 3918 2358 3922 2362
rect 3926 2358 3930 2362
rect 3902 2340 3906 2344
rect 3878 2328 3882 2332
rect 3886 2328 3890 2332
rect 3758 2318 3762 2322
rect 3774 2318 3778 2322
rect 3750 2308 3754 2312
rect 3878 2298 3882 2302
rect 3742 2288 3746 2292
rect 3766 2288 3770 2292
rect 3854 2288 3858 2292
rect 3878 2288 3882 2292
rect 3734 2278 3738 2282
rect 3942 2338 3946 2342
rect 3966 2368 3970 2372
rect 4054 2378 4058 2382
rect 4070 2378 4074 2382
rect 4006 2368 4010 2372
rect 4030 2368 4034 2372
rect 4062 2368 4066 2372
rect 3974 2348 3978 2352
rect 3982 2338 3986 2342
rect 3998 2338 4002 2342
rect 4118 2448 4122 2452
rect 4142 2428 4146 2432
rect 4134 2378 4138 2382
rect 4110 2368 4114 2372
rect 4126 2368 4130 2372
rect 4094 2358 4098 2362
rect 4118 2358 4122 2362
rect 4046 2348 4050 2352
rect 4070 2348 4074 2352
rect 4078 2348 4082 2352
rect 4014 2338 4018 2342
rect 4214 2458 4218 2462
rect 4174 2448 4178 2452
rect 4206 2448 4210 2452
rect 4222 2448 4226 2452
rect 4150 2418 4154 2422
rect 4190 2428 4194 2432
rect 4206 2428 4210 2432
rect 4166 2418 4170 2422
rect 4158 2388 4162 2392
rect 4174 2408 4178 2412
rect 4262 2458 4266 2462
rect 4254 2358 4258 2362
rect 4182 2348 4186 2352
rect 4142 2338 4146 2342
rect 4166 2338 4170 2342
rect 4078 2328 4082 2332
rect 4126 2328 4130 2332
rect 3958 2318 3962 2322
rect 3910 2308 3914 2312
rect 3930 2303 3934 2307
rect 3937 2303 3941 2307
rect 3926 2288 3930 2292
rect 3758 2278 3762 2282
rect 3886 2278 3890 2282
rect 3894 2278 3898 2282
rect 3918 2278 3922 2282
rect 3718 2248 3722 2252
rect 3694 2228 3698 2232
rect 3694 2218 3698 2222
rect 3670 2168 3674 2172
rect 3742 2208 3746 2212
rect 3718 2198 3722 2202
rect 3678 2148 3682 2152
rect 3790 2268 3794 2272
rect 3766 2258 3770 2262
rect 3782 2248 3786 2252
rect 3806 2248 3810 2252
rect 3846 2258 3850 2262
rect 3854 2258 3858 2262
rect 3790 2238 3794 2242
rect 3814 2238 3818 2242
rect 3846 2228 3850 2232
rect 3902 2268 3906 2272
rect 3902 2238 3906 2242
rect 3870 2218 3874 2222
rect 3910 2218 3914 2222
rect 3846 2168 3850 2172
rect 3910 2158 3914 2162
rect 3942 2278 3946 2282
rect 3934 2268 3938 2272
rect 3942 2248 3946 2252
rect 3926 2238 3930 2242
rect 3926 2158 3930 2162
rect 3798 2148 3802 2152
rect 3830 2148 3834 2152
rect 3902 2148 3906 2152
rect 4206 2338 4210 2342
rect 4198 2308 4202 2312
rect 4310 2458 4314 2462
rect 4278 2448 4282 2452
rect 4566 2548 4570 2552
rect 4574 2548 4578 2552
rect 4526 2538 4530 2542
rect 4622 2538 4626 2542
rect 4510 2528 4514 2532
rect 4430 2518 4434 2522
rect 4390 2508 4394 2512
rect 4406 2468 4410 2472
rect 4590 2528 4594 2532
rect 4534 2508 4538 2512
rect 4558 2508 4562 2512
rect 4630 2508 4634 2512
rect 4654 2588 4658 2592
rect 4542 2488 4546 2492
rect 4486 2478 4490 2482
rect 4462 2468 4466 2472
rect 4358 2448 4362 2452
rect 4390 2448 4394 2452
rect 4422 2448 4426 2452
rect 4462 2448 4466 2452
rect 4478 2448 4482 2452
rect 4510 2468 4514 2472
rect 4534 2468 4538 2472
rect 4510 2458 4514 2462
rect 4518 2448 4522 2452
rect 4350 2398 4354 2402
rect 4326 2388 4330 2392
rect 4270 2368 4274 2372
rect 4334 2368 4338 2372
rect 4278 2358 4282 2362
rect 4302 2358 4306 2362
rect 4262 2348 4266 2352
rect 4278 2338 4282 2342
rect 4302 2338 4306 2342
rect 4270 2328 4274 2332
rect 3966 2288 3970 2292
rect 4022 2288 4026 2292
rect 3990 2278 3994 2282
rect 4078 2278 4082 2282
rect 4134 2278 4138 2282
rect 4166 2278 4170 2282
rect 3982 2268 3986 2272
rect 4014 2268 4018 2272
rect 4030 2268 4034 2272
rect 4102 2268 4106 2272
rect 4110 2268 4114 2272
rect 4158 2268 4162 2272
rect 4014 2258 4018 2262
rect 4054 2258 4058 2262
rect 4094 2258 4098 2262
rect 4102 2258 4106 2262
rect 4134 2258 4138 2262
rect 4150 2258 4154 2262
rect 4054 2248 4058 2252
rect 4022 2228 4026 2232
rect 4062 2228 4066 2232
rect 4030 2218 4034 2222
rect 3998 2198 4002 2202
rect 3990 2178 3994 2182
rect 3990 2168 3994 2172
rect 3982 2148 3986 2152
rect 4062 2188 4066 2192
rect 4062 2168 4066 2172
rect 4094 2168 4098 2172
rect 4022 2158 4026 2162
rect 3750 2138 3754 2142
rect 3846 2138 3850 2142
rect 3910 2138 3914 2142
rect 3206 2038 3210 2042
rect 3214 2038 3218 2042
rect 3254 2038 3258 2042
rect 3294 2038 3298 2042
rect 3286 2018 3290 2022
rect 3310 2018 3314 2022
rect 3190 1998 3194 2002
rect 3318 1968 3322 1972
rect 3238 1958 3242 1962
rect 3254 1958 3258 1962
rect 3310 1958 3314 1962
rect 3198 1948 3202 1952
rect 3214 1948 3218 1952
rect 3214 1938 3218 1942
rect 3190 1918 3194 1922
rect 3230 1918 3234 1922
rect 3214 1908 3218 1912
rect 3158 1888 3162 1892
rect 3262 1938 3266 1942
rect 3350 2068 3354 2072
rect 3366 2068 3370 2072
rect 3358 2058 3362 2062
rect 3374 2058 3378 2062
rect 3342 2048 3346 2052
rect 3366 2038 3370 2042
rect 3358 2028 3362 2032
rect 3366 2028 3370 2032
rect 3358 1958 3362 1962
rect 3366 1948 3370 1952
rect 3390 2068 3394 2072
rect 3454 2118 3458 2122
rect 3414 2098 3418 2102
rect 3486 2108 3490 2112
rect 3502 2098 3506 2102
rect 3654 2088 3658 2092
rect 3710 2088 3714 2092
rect 3726 2088 3730 2092
rect 3422 2078 3426 2082
rect 3430 2068 3434 2072
rect 3494 2068 3498 2072
rect 3502 2068 3506 2072
rect 3566 2078 3570 2082
rect 3622 2078 3626 2082
rect 3630 2078 3634 2082
rect 3758 2078 3762 2082
rect 3830 2128 3834 2132
rect 3838 2128 3842 2132
rect 3854 2128 3858 2132
rect 3870 2108 3874 2112
rect 4006 2128 4010 2132
rect 4022 2128 4026 2132
rect 4030 2128 4034 2132
rect 4150 2188 4154 2192
rect 4102 2158 4106 2162
rect 4078 2128 4082 2132
rect 4094 2128 4098 2132
rect 4038 2118 4042 2122
rect 4054 2118 4058 2122
rect 4142 2118 4146 2122
rect 3930 2103 3934 2107
rect 3937 2103 3941 2107
rect 3822 2078 3826 2082
rect 3798 2068 3802 2072
rect 3966 2068 3970 2072
rect 3438 2058 3442 2062
rect 3438 2048 3442 2052
rect 3414 2038 3418 2042
rect 3406 2028 3410 2032
rect 3454 2028 3458 2032
rect 3418 2003 3422 2007
rect 3425 2003 3429 2007
rect 3406 1958 3410 1962
rect 3550 2058 3554 2062
rect 3574 2058 3578 2062
rect 3470 2048 3474 2052
rect 3558 2048 3562 2052
rect 3590 2048 3594 2052
rect 3606 2048 3610 2052
rect 3534 2038 3538 2042
rect 3462 2018 3466 2022
rect 3478 2018 3482 2022
rect 3542 2018 3546 2022
rect 3654 2018 3658 2022
rect 3606 1988 3610 1992
rect 3534 1968 3538 1972
rect 3398 1948 3402 1952
rect 3510 1948 3514 1952
rect 3294 1938 3298 1942
rect 3334 1938 3338 1942
rect 3358 1938 3362 1942
rect 3278 1928 3282 1932
rect 3398 1908 3402 1912
rect 3534 1928 3538 1932
rect 3486 1918 3490 1922
rect 3510 1918 3514 1922
rect 3566 1918 3570 1922
rect 3582 1918 3586 1922
rect 3598 1918 3602 1922
rect 3486 1908 3490 1912
rect 3542 1908 3546 1912
rect 3838 2048 3842 2052
rect 3734 2038 3738 2042
rect 3686 2028 3690 2032
rect 3750 2028 3754 2032
rect 3750 1998 3754 2002
rect 3678 1988 3682 1992
rect 3902 1958 3906 1962
rect 3694 1948 3698 1952
rect 3750 1948 3754 1952
rect 3326 1888 3330 1892
rect 3350 1888 3354 1892
rect 3390 1888 3394 1892
rect 3406 1888 3410 1892
rect 3478 1888 3482 1892
rect 3158 1868 3162 1872
rect 3102 1848 3106 1852
rect 3150 1848 3154 1852
rect 3190 1868 3194 1872
rect 3254 1868 3258 1872
rect 3214 1858 3218 1862
rect 3198 1848 3202 1852
rect 3206 1848 3210 1852
rect 3134 1818 3138 1822
rect 3174 1818 3178 1822
rect 3190 1818 3194 1822
rect 3270 1808 3274 1812
rect 3190 1778 3194 1782
rect 3182 1768 3186 1772
rect 3166 1758 3170 1762
rect 3094 1748 3098 1752
rect 3110 1718 3114 1722
rect 3078 1708 3082 1712
rect 3054 1698 3058 1702
rect 3078 1698 3082 1702
rect 3046 1678 3050 1682
rect 3022 1658 3026 1662
rect 3078 1658 3082 1662
rect 2910 1648 2914 1652
rect 2918 1618 2922 1622
rect 2790 1608 2794 1612
rect 2766 1568 2770 1572
rect 2606 1548 2610 1552
rect 2670 1548 2674 1552
rect 2702 1548 2706 1552
rect 2750 1548 2754 1552
rect 2974 1588 2978 1592
rect 2822 1548 2826 1552
rect 2718 1528 2722 1532
rect 2606 1488 2610 1492
rect 2654 1488 2658 1492
rect 2670 1488 2674 1492
rect 2718 1478 2722 1482
rect 2710 1468 2714 1472
rect 2758 1468 2762 1472
rect 2878 1528 2882 1532
rect 2998 1558 3002 1562
rect 3094 1608 3098 1612
rect 3086 1558 3090 1562
rect 3038 1548 3042 1552
rect 2974 1538 2978 1542
rect 3038 1538 3042 1542
rect 2918 1518 2922 1522
rect 2906 1503 2910 1507
rect 2913 1503 2917 1507
rect 2846 1498 2850 1502
rect 2950 1518 2954 1522
rect 2982 1518 2986 1522
rect 3006 1518 3010 1522
rect 2974 1498 2978 1502
rect 2902 1488 2906 1492
rect 2926 1488 2930 1492
rect 2862 1478 2866 1482
rect 3086 1488 3090 1492
rect 2998 1478 3002 1482
rect 3022 1478 3026 1482
rect 2926 1468 2930 1472
rect 3014 1468 3018 1472
rect 3046 1468 3050 1472
rect 2774 1458 2778 1462
rect 2462 1448 2466 1452
rect 2630 1448 2634 1452
rect 2694 1448 2698 1452
rect 2710 1448 2714 1452
rect 2750 1448 2754 1452
rect 2454 1438 2458 1442
rect 2654 1438 2658 1442
rect 2438 1428 2442 1432
rect 2638 1428 2642 1432
rect 2526 1418 2530 1422
rect 2550 1418 2554 1422
rect 2230 1378 2234 1382
rect 2246 1378 2250 1382
rect 2342 1378 2346 1382
rect 2394 1403 2398 1407
rect 2401 1403 2405 1407
rect 2470 1378 2474 1382
rect 2198 1358 2202 1362
rect 2246 1358 2250 1362
rect 2270 1358 2274 1362
rect 2326 1358 2330 1362
rect 2350 1358 2354 1362
rect 2382 1358 2386 1362
rect 2398 1358 2402 1362
rect 2182 1348 2186 1352
rect 2190 1348 2194 1352
rect 2246 1348 2250 1352
rect 2110 1338 2114 1342
rect 2046 1298 2050 1302
rect 2054 1278 2058 1282
rect 2070 1278 2074 1282
rect 2126 1328 2130 1332
rect 1854 1268 1858 1272
rect 1942 1268 1946 1272
rect 2054 1268 2058 1272
rect 1878 1258 1882 1262
rect 1766 1248 1770 1252
rect 1782 1248 1786 1252
rect 1822 1248 1826 1252
rect 1694 1228 1698 1232
rect 1758 1228 1762 1232
rect 1910 1258 1914 1262
rect 1998 1259 2002 1263
rect 1894 1208 1898 1212
rect 1782 1178 1786 1182
rect 1902 1178 1906 1182
rect 1686 1158 1690 1162
rect 1670 1148 1674 1152
rect 1702 1148 1706 1152
rect 1638 1138 1642 1142
rect 1662 1138 1666 1142
rect 1654 1108 1658 1112
rect 1774 1138 1778 1142
rect 1694 1098 1698 1102
rect 1622 1088 1626 1092
rect 1630 1088 1634 1092
rect 1654 1088 1658 1092
rect 1902 1168 1906 1172
rect 1958 1208 1962 1212
rect 2406 1348 2410 1352
rect 2422 1348 2426 1352
rect 2214 1338 2218 1342
rect 2238 1338 2242 1342
rect 2286 1338 2290 1342
rect 2166 1328 2170 1332
rect 2182 1328 2186 1332
rect 2262 1328 2266 1332
rect 2150 1278 2154 1282
rect 2182 1278 2186 1282
rect 2998 1458 3002 1462
rect 3038 1458 3042 1462
rect 3094 1458 3098 1462
rect 3142 1718 3146 1722
rect 3254 1748 3258 1752
rect 3238 1728 3242 1732
rect 3334 1868 3338 1872
rect 3342 1858 3346 1862
rect 3358 1858 3362 1862
rect 3422 1868 3426 1872
rect 3566 1868 3570 1872
rect 3390 1858 3394 1862
rect 3406 1858 3410 1862
rect 3334 1848 3338 1852
rect 3366 1848 3370 1852
rect 3398 1838 3402 1842
rect 3302 1738 3306 1742
rect 3334 1738 3338 1742
rect 3438 1848 3442 1852
rect 3418 1803 3422 1807
rect 3425 1803 3429 1807
rect 3742 1928 3746 1932
rect 3630 1918 3634 1922
rect 3694 1918 3698 1922
rect 3702 1918 3706 1922
rect 3686 1878 3690 1882
rect 3878 1947 3882 1951
rect 3934 1948 3938 1952
rect 3950 1948 3954 1952
rect 3742 1908 3746 1912
rect 3790 1908 3794 1912
rect 3930 1903 3934 1907
rect 3937 1903 3941 1907
rect 3950 1898 3954 1902
rect 3774 1888 3778 1892
rect 3846 1888 3850 1892
rect 3622 1858 3626 1862
rect 3502 1748 3506 1752
rect 3590 1748 3594 1752
rect 3494 1738 3498 1742
rect 3510 1738 3514 1742
rect 3518 1738 3522 1742
rect 3534 1738 3538 1742
rect 3558 1738 3562 1742
rect 3566 1738 3570 1742
rect 3462 1728 3466 1732
rect 3486 1728 3490 1732
rect 3462 1718 3466 1722
rect 3342 1708 3346 1712
rect 3390 1708 3394 1712
rect 3422 1698 3426 1702
rect 3334 1688 3338 1692
rect 3374 1688 3378 1692
rect 3318 1678 3322 1682
rect 3366 1678 3370 1682
rect 3294 1668 3298 1672
rect 3302 1668 3306 1672
rect 3246 1659 3250 1663
rect 3118 1618 3122 1622
rect 3190 1648 3194 1652
rect 3134 1588 3138 1592
rect 3254 1608 3258 1612
rect 3150 1568 3154 1572
rect 3302 1648 3306 1652
rect 3318 1638 3322 1642
rect 3134 1558 3138 1562
rect 3190 1558 3194 1562
rect 3150 1548 3154 1552
rect 3254 1548 3258 1552
rect 3110 1498 3114 1502
rect 3246 1538 3250 1542
rect 3262 1538 3266 1542
rect 3230 1508 3234 1512
rect 3222 1498 3226 1502
rect 3278 1488 3282 1492
rect 3190 1478 3194 1482
rect 3286 1478 3290 1482
rect 3214 1468 3218 1472
rect 3246 1468 3250 1472
rect 3174 1458 3178 1462
rect 2958 1448 2962 1452
rect 3102 1448 3106 1452
rect 3158 1448 3162 1452
rect 2790 1438 2794 1442
rect 2846 1438 2850 1442
rect 3014 1438 3018 1442
rect 3046 1438 3050 1442
rect 2678 1408 2682 1412
rect 2726 1398 2730 1402
rect 2870 1418 2874 1422
rect 2862 1408 2866 1412
rect 2686 1378 2690 1382
rect 2750 1378 2754 1382
rect 2806 1378 2810 1382
rect 2606 1358 2610 1362
rect 2662 1358 2666 1362
rect 2550 1348 2554 1352
rect 2374 1338 2378 1342
rect 2390 1338 2394 1342
rect 2534 1338 2538 1342
rect 2710 1338 2714 1342
rect 2310 1318 2314 1322
rect 2294 1308 2298 1312
rect 2198 1278 2202 1282
rect 2286 1278 2290 1282
rect 2310 1278 2314 1282
rect 2086 1268 2090 1272
rect 2102 1268 2106 1272
rect 2110 1268 2114 1272
rect 2126 1268 2130 1272
rect 2158 1268 2162 1272
rect 2254 1268 2258 1272
rect 2294 1268 2298 1272
rect 2310 1268 2314 1272
rect 2046 1258 2050 1262
rect 2046 1248 2050 1252
rect 2086 1248 2090 1252
rect 2086 1228 2090 1232
rect 2022 1188 2026 1192
rect 2070 1178 2074 1182
rect 1806 1158 1810 1162
rect 1830 1158 1834 1162
rect 1854 1158 1858 1162
rect 1990 1158 1994 1162
rect 2054 1158 2058 1162
rect 1798 1128 1802 1132
rect 1814 1128 1818 1132
rect 1846 1148 1850 1152
rect 1862 1138 1866 1142
rect 1790 1118 1794 1122
rect 1814 1118 1818 1122
rect 1830 1118 1834 1122
rect 1874 1103 1878 1107
rect 1881 1103 1885 1107
rect 2094 1168 2098 1172
rect 2094 1158 2098 1162
rect 2038 1148 2042 1152
rect 1910 1138 1914 1142
rect 1942 1138 1946 1142
rect 1966 1138 1970 1142
rect 1934 1128 1938 1132
rect 2134 1248 2138 1252
rect 2150 1158 2154 1162
rect 2110 1148 2114 1152
rect 2142 1148 2146 1152
rect 2054 1138 2058 1142
rect 2110 1138 2114 1142
rect 2134 1138 2138 1142
rect 1982 1128 1986 1132
rect 1958 1118 1962 1122
rect 1950 1108 1954 1112
rect 2038 1128 2042 1132
rect 2014 1108 2018 1112
rect 2006 1088 2010 1092
rect 1742 1078 1746 1082
rect 1758 1078 1762 1082
rect 1846 1078 1850 1082
rect 1966 1078 1970 1082
rect 1990 1078 1994 1082
rect 1814 1068 1818 1072
rect 1830 1068 1834 1072
rect 1854 1068 1858 1072
rect 1606 1038 1610 1042
rect 1598 1028 1602 1032
rect 1534 1018 1538 1022
rect 1494 1008 1498 1012
rect 1478 988 1482 992
rect 1494 958 1498 962
rect 1470 928 1474 932
rect 1422 918 1426 922
rect 1486 918 1490 922
rect 1390 888 1394 892
rect 1414 878 1418 882
rect 1590 998 1594 1002
rect 1534 978 1538 982
rect 1566 968 1570 972
rect 1534 958 1538 962
rect 1542 958 1546 962
rect 1510 928 1514 932
rect 1558 928 1562 932
rect 1582 928 1586 932
rect 1510 878 1514 882
rect 1342 868 1346 872
rect 1382 858 1386 862
rect 1502 858 1506 862
rect 1294 848 1298 852
rect 1302 848 1306 852
rect 1086 838 1090 842
rect 1110 838 1114 842
rect 1134 838 1138 842
rect 1342 838 1346 842
rect 1078 828 1082 832
rect 1166 828 1170 832
rect 1254 828 1258 832
rect 1334 828 1338 832
rect 1094 818 1098 822
rect 1142 798 1146 802
rect 1230 808 1234 812
rect 1126 768 1130 772
rect 1150 768 1154 772
rect 1166 768 1170 772
rect 1118 758 1122 762
rect 1014 748 1018 752
rect 1046 748 1050 752
rect 990 728 994 732
rect 1030 728 1034 732
rect 1086 728 1090 732
rect 982 718 986 722
rect 1022 698 1026 702
rect 1182 758 1186 762
rect 1310 798 1314 802
rect 1342 768 1346 772
rect 1262 758 1266 762
rect 1150 748 1154 752
rect 1142 738 1146 742
rect 1174 738 1178 742
rect 1182 738 1186 742
rect 1134 698 1138 702
rect 1166 698 1170 702
rect 1030 688 1034 692
rect 1078 688 1082 692
rect 1094 688 1098 692
rect 1006 678 1010 682
rect 1310 748 1314 752
rect 1302 738 1306 742
rect 1438 828 1442 832
rect 1430 818 1434 822
rect 1370 803 1374 807
rect 1377 803 1381 807
rect 1358 798 1362 802
rect 1430 798 1434 802
rect 1406 758 1410 762
rect 1446 798 1450 802
rect 1606 958 1610 962
rect 1614 938 1618 942
rect 1606 928 1610 932
rect 1622 928 1626 932
rect 1726 1048 1730 1052
rect 1942 1068 1946 1072
rect 2110 1118 2114 1122
rect 2126 1098 2130 1102
rect 2054 1088 2058 1092
rect 1846 1058 1850 1062
rect 1878 1058 1882 1062
rect 1926 1058 1930 1062
rect 1942 1058 1946 1062
rect 1838 1048 1842 1052
rect 1910 1048 1914 1052
rect 1966 1048 1970 1052
rect 1742 1038 1746 1042
rect 2038 1038 2042 1042
rect 1718 988 1722 992
rect 1702 978 1706 982
rect 1750 978 1754 982
rect 1758 978 1762 982
rect 1686 958 1690 962
rect 1718 958 1722 962
rect 1838 958 1842 962
rect 2022 958 2026 962
rect 1686 948 1690 952
rect 1702 948 1706 952
rect 1734 948 1738 952
rect 1846 948 1850 952
rect 1886 948 1890 952
rect 2142 1088 2146 1092
rect 2142 1078 2146 1082
rect 2070 1058 2074 1062
rect 1782 938 1786 942
rect 1670 928 1674 932
rect 1758 928 1762 932
rect 1654 918 1658 922
rect 1726 898 1730 902
rect 1790 928 1794 932
rect 1814 918 1818 922
rect 1870 938 1874 942
rect 1934 938 1938 942
rect 2134 1058 2138 1062
rect 2102 1008 2106 1012
rect 2126 958 2130 962
rect 2142 958 2146 962
rect 2094 948 2098 952
rect 2134 948 2138 952
rect 2102 938 2106 942
rect 2118 938 2122 942
rect 2166 1178 2170 1182
rect 2190 1168 2194 1172
rect 2270 1258 2274 1262
rect 2302 1258 2306 1262
rect 2214 1248 2218 1252
rect 2254 1238 2258 1242
rect 2198 1158 2202 1162
rect 2206 1158 2210 1162
rect 2230 1158 2234 1162
rect 2174 1148 2178 1152
rect 2286 1198 2290 1202
rect 2310 1188 2314 1192
rect 2270 1158 2274 1162
rect 2182 1138 2186 1142
rect 2166 1108 2170 1112
rect 2158 1098 2162 1102
rect 2166 1088 2170 1092
rect 2174 1078 2178 1082
rect 2214 1078 2218 1082
rect 2190 1068 2194 1072
rect 2270 1148 2274 1152
rect 2262 1108 2266 1112
rect 2294 1078 2298 1082
rect 2230 1058 2234 1062
rect 2310 1058 2314 1062
rect 2174 1048 2178 1052
rect 2278 1048 2282 1052
rect 2302 1048 2306 1052
rect 2214 1038 2218 1042
rect 2270 1038 2274 1042
rect 2190 1018 2194 1022
rect 2166 978 2170 982
rect 2054 928 2058 932
rect 2078 928 2082 932
rect 1918 908 1922 912
rect 1874 903 1878 907
rect 1881 903 1885 907
rect 1774 898 1778 902
rect 1846 898 1850 902
rect 1878 888 1882 892
rect 1950 888 1954 892
rect 1902 878 1906 882
rect 1974 878 1978 882
rect 1990 868 1994 872
rect 1606 858 1610 862
rect 1542 848 1546 852
rect 1558 848 1562 852
rect 1630 848 1634 852
rect 1606 838 1610 842
rect 1454 768 1458 772
rect 1462 768 1466 772
rect 1502 768 1506 772
rect 1518 768 1522 772
rect 1526 768 1530 772
rect 1550 768 1554 772
rect 1574 768 1578 772
rect 1478 758 1482 762
rect 1510 758 1514 762
rect 1542 758 1546 762
rect 1374 748 1378 752
rect 1446 748 1450 752
rect 1470 748 1474 752
rect 1486 748 1490 752
rect 1334 738 1338 742
rect 1558 748 1562 752
rect 1590 748 1594 752
rect 1542 738 1546 742
rect 1582 738 1586 742
rect 1206 728 1210 732
rect 1326 728 1330 732
rect 1366 728 1370 732
rect 1382 728 1386 732
rect 1414 728 1418 732
rect 1438 728 1442 732
rect 1446 728 1450 732
rect 1486 728 1490 732
rect 1590 728 1594 732
rect 1598 728 1602 732
rect 1318 718 1322 722
rect 1470 718 1474 722
rect 1150 688 1154 692
rect 1246 688 1250 692
rect 1310 678 1314 682
rect 1022 668 1026 672
rect 1038 668 1042 672
rect 910 658 914 662
rect 966 658 970 662
rect 990 658 994 662
rect 1022 658 1026 662
rect 1046 658 1050 662
rect 982 648 986 652
rect 902 638 906 642
rect 942 628 946 632
rect 742 568 746 572
rect 814 568 818 572
rect 710 558 714 562
rect 718 548 722 552
rect 838 558 842 562
rect 774 548 778 552
rect 830 548 834 552
rect 710 538 714 542
rect 750 538 754 542
rect 782 538 786 542
rect 726 528 730 532
rect 758 528 762 532
rect 662 508 666 512
rect 686 508 690 512
rect 798 528 802 532
rect 766 498 770 502
rect 790 498 794 502
rect 886 618 890 622
rect 902 618 906 622
rect 886 598 890 602
rect 1046 608 1050 612
rect 1022 598 1026 602
rect 1038 598 1042 602
rect 990 588 994 592
rect 862 568 866 572
rect 966 568 970 572
rect 870 548 874 552
rect 910 548 914 552
rect 886 528 890 532
rect 902 528 906 532
rect 910 528 914 532
rect 1030 558 1034 562
rect 1022 548 1026 552
rect 966 538 970 542
rect 982 538 986 542
rect 1014 538 1018 542
rect 934 518 938 522
rect 958 518 962 522
rect 858 503 862 507
rect 865 503 869 507
rect 886 498 890 502
rect 822 488 826 492
rect 670 478 674 482
rect 798 478 802 482
rect 838 478 842 482
rect 654 418 658 422
rect 678 468 682 472
rect 734 468 738 472
rect 686 448 690 452
rect 710 438 714 442
rect 774 468 778 472
rect 790 468 794 472
rect 766 458 770 462
rect 862 468 866 472
rect 798 458 802 462
rect 822 458 826 462
rect 870 448 874 452
rect 758 438 762 442
rect 718 428 722 432
rect 742 428 746 432
rect 830 418 834 422
rect 846 418 850 422
rect 718 368 722 372
rect 750 368 754 372
rect 662 358 666 362
rect 710 358 714 362
rect 662 348 666 352
rect 694 348 698 352
rect 702 338 706 342
rect 782 358 786 362
rect 798 358 802 362
rect 830 358 834 362
rect 854 358 858 362
rect 750 348 754 352
rect 734 340 738 344
rect 910 458 914 462
rect 942 458 946 462
rect 950 458 954 462
rect 958 448 962 452
rect 926 438 930 442
rect 990 438 994 442
rect 950 428 954 432
rect 894 418 898 422
rect 910 418 914 422
rect 966 418 970 422
rect 974 418 978 422
rect 982 378 986 382
rect 926 368 930 372
rect 878 348 882 352
rect 1014 448 1018 452
rect 1006 438 1010 442
rect 998 428 1002 432
rect 1030 528 1034 532
rect 1102 618 1106 622
rect 1118 648 1122 652
rect 1150 648 1154 652
rect 1126 638 1130 642
rect 1134 638 1138 642
rect 1126 628 1130 632
rect 1102 608 1106 612
rect 1070 568 1074 572
rect 1574 708 1578 712
rect 1766 858 1770 862
rect 1798 858 1802 862
rect 1846 848 1850 852
rect 1646 838 1650 842
rect 1742 828 1746 832
rect 1830 798 1834 802
rect 1870 838 1874 842
rect 1894 838 1898 842
rect 1710 788 1714 792
rect 1862 788 1866 792
rect 1662 748 1666 752
rect 1686 748 1690 752
rect 1718 778 1722 782
rect 1862 768 1866 772
rect 1790 758 1794 762
rect 1814 748 1818 752
rect 1710 738 1714 742
rect 1686 718 1690 722
rect 1806 728 1810 732
rect 1854 718 1858 722
rect 1886 718 1890 722
rect 1774 698 1778 702
rect 1366 688 1370 692
rect 1606 688 1610 692
rect 1750 688 1754 692
rect 1502 678 1506 682
rect 1254 668 1258 672
rect 1166 658 1170 662
rect 1182 648 1186 652
rect 1158 558 1162 562
rect 1222 648 1226 652
rect 1198 638 1202 642
rect 1230 638 1234 642
rect 1390 658 1394 662
rect 1278 648 1282 652
rect 1422 648 1426 652
rect 1238 608 1242 612
rect 1334 638 1338 642
rect 1438 638 1442 642
rect 1254 568 1258 572
rect 1230 558 1234 562
rect 1182 548 1186 552
rect 1342 598 1346 602
rect 1078 538 1082 542
rect 1070 508 1074 512
rect 1086 508 1090 512
rect 1110 498 1114 502
rect 1158 498 1162 502
rect 1566 658 1570 662
rect 1478 628 1482 632
rect 1494 628 1498 632
rect 1446 608 1450 612
rect 1370 603 1374 607
rect 1377 603 1381 607
rect 1446 598 1450 602
rect 1350 588 1354 592
rect 1406 568 1410 572
rect 1726 678 1730 682
rect 1874 703 1878 707
rect 1881 703 1885 707
rect 1830 678 1834 682
rect 1910 758 1914 762
rect 1902 728 1906 732
rect 1998 858 2002 862
rect 1974 848 1978 852
rect 1966 828 1970 832
rect 1934 778 1938 782
rect 1926 758 1930 762
rect 1950 768 1954 772
rect 1958 768 1962 772
rect 1614 668 1618 672
rect 1670 668 1674 672
rect 1902 668 1906 672
rect 1630 659 1634 663
rect 1806 658 1810 662
rect 1726 598 1730 602
rect 1574 568 1578 572
rect 1494 558 1498 562
rect 1550 558 1554 562
rect 1662 558 1666 562
rect 1414 548 1418 552
rect 1214 538 1218 542
rect 1486 548 1490 552
rect 1542 538 1546 542
rect 1630 538 1634 542
rect 1694 538 1698 542
rect 1190 488 1194 492
rect 1166 478 1170 482
rect 1206 478 1210 482
rect 1142 468 1146 472
rect 1174 468 1178 472
rect 1078 458 1082 462
rect 1070 418 1074 422
rect 1174 438 1178 442
rect 1094 348 1098 352
rect 806 338 810 342
rect 838 338 842 342
rect 926 338 930 342
rect 1046 338 1050 342
rect 1102 338 1106 342
rect 606 328 610 332
rect 646 328 650 332
rect 662 328 666 332
rect 694 328 698 332
rect 726 328 730 332
rect 758 328 762 332
rect 750 308 754 312
rect 694 298 698 302
rect 726 298 730 302
rect 526 268 530 272
rect 622 238 626 242
rect 582 208 586 212
rect 558 178 562 182
rect 574 178 578 182
rect 470 168 474 172
rect 542 168 546 172
rect 374 158 378 162
rect 398 158 402 162
rect 334 148 338 152
rect 414 148 418 152
rect 342 138 346 142
rect 174 118 178 122
rect 126 78 130 82
rect 246 98 250 102
rect 110 68 114 72
rect 142 66 146 70
rect 238 68 242 72
rect 62 58 66 62
rect 94 58 98 62
rect 166 58 170 62
rect 174 58 178 62
rect 446 138 450 142
rect 438 128 442 132
rect 302 98 306 102
rect 262 88 266 92
rect 294 88 298 92
rect 262 68 266 72
rect 422 88 426 92
rect 502 158 506 162
rect 518 158 522 162
rect 486 148 490 152
rect 494 138 498 142
rect 534 148 538 152
rect 566 168 570 172
rect 590 168 594 172
rect 678 258 682 262
rect 710 258 714 262
rect 670 248 674 252
rect 766 308 770 312
rect 766 298 770 302
rect 758 278 762 282
rect 750 258 754 262
rect 814 328 818 332
rect 862 328 866 332
rect 638 238 642 242
rect 686 238 690 242
rect 718 238 722 242
rect 750 238 754 242
rect 782 238 786 242
rect 798 238 802 242
rect 726 228 730 232
rect 726 208 730 212
rect 750 198 754 202
rect 806 198 810 202
rect 638 178 642 182
rect 654 178 658 182
rect 790 178 794 182
rect 702 168 706 172
rect 790 168 794 172
rect 574 158 578 162
rect 582 158 586 162
rect 598 158 602 162
rect 630 158 634 162
rect 558 148 562 152
rect 630 148 634 152
rect 646 148 650 152
rect 710 148 714 152
rect 534 138 538 142
rect 542 138 546 142
rect 478 118 482 122
rect 470 88 474 92
rect 510 88 514 92
rect 318 78 322 82
rect 366 78 370 82
rect 454 78 458 82
rect 462 78 466 82
rect 598 138 602 142
rect 654 138 658 142
rect 558 128 562 132
rect 582 128 586 132
rect 598 128 602 132
rect 566 88 570 92
rect 654 88 658 92
rect 494 78 498 82
rect 550 78 554 82
rect 838 318 842 322
rect 858 303 862 307
rect 865 303 869 307
rect 838 298 842 302
rect 1046 298 1050 302
rect 1078 298 1082 302
rect 886 288 890 292
rect 1262 528 1266 532
rect 1222 518 1226 522
rect 1286 518 1290 522
rect 1310 518 1314 522
rect 1406 528 1410 532
rect 1366 518 1370 522
rect 1318 508 1322 512
rect 1342 508 1346 512
rect 1494 528 1498 532
rect 1462 518 1466 522
rect 1462 498 1466 502
rect 1438 488 1442 492
rect 1222 468 1226 472
rect 1254 468 1258 472
rect 1230 448 1234 452
rect 1454 468 1458 472
rect 1294 458 1298 462
rect 1350 458 1354 462
rect 1246 438 1250 442
rect 1270 438 1274 442
rect 1406 448 1410 452
rect 1422 448 1426 452
rect 1374 428 1378 432
rect 1390 408 1394 412
rect 1370 403 1374 407
rect 1377 403 1381 407
rect 1198 388 1202 392
rect 1574 528 1578 532
rect 1622 528 1626 532
rect 1590 518 1594 522
rect 1526 478 1530 482
rect 1558 478 1562 482
rect 1542 468 1546 472
rect 1550 468 1554 472
rect 1526 448 1530 452
rect 1534 448 1538 452
rect 1502 388 1506 392
rect 1390 378 1394 382
rect 1542 378 1546 382
rect 1550 378 1554 382
rect 1358 368 1362 372
rect 1270 348 1274 352
rect 1302 348 1306 352
rect 1374 348 1378 352
rect 1326 338 1330 342
rect 1334 338 1338 342
rect 1382 338 1386 342
rect 1422 338 1426 342
rect 1438 338 1442 342
rect 1142 328 1146 332
rect 1110 318 1114 322
rect 1174 318 1178 322
rect 1190 318 1194 322
rect 1198 308 1202 312
rect 1238 298 1242 302
rect 1206 288 1210 292
rect 982 278 986 282
rect 1038 278 1042 282
rect 1086 278 1090 282
rect 1134 278 1138 282
rect 1022 268 1026 272
rect 814 178 818 182
rect 934 258 938 262
rect 958 258 962 262
rect 974 258 978 262
rect 918 238 922 242
rect 942 238 946 242
rect 830 168 834 172
rect 910 168 914 172
rect 798 148 802 152
rect 910 148 914 152
rect 918 148 922 152
rect 998 228 1002 232
rect 958 218 962 222
rect 950 208 954 212
rect 1038 258 1042 262
rect 1030 228 1034 232
rect 1022 218 1026 222
rect 1038 218 1042 222
rect 1014 188 1018 192
rect 1046 198 1050 202
rect 1262 328 1266 332
rect 1270 328 1274 332
rect 1350 328 1354 332
rect 1206 268 1210 272
rect 1078 208 1082 212
rect 1078 198 1082 202
rect 1094 238 1098 242
rect 1118 208 1122 212
rect 670 128 674 132
rect 822 138 826 142
rect 838 138 842 142
rect 894 138 898 142
rect 934 138 938 142
rect 958 138 962 142
rect 1030 138 1034 142
rect 1070 138 1074 142
rect 782 128 786 132
rect 846 128 850 132
rect 918 128 922 132
rect 942 128 946 132
rect 1030 128 1034 132
rect 718 118 722 122
rect 854 118 858 122
rect 702 78 706 82
rect 310 68 314 72
rect 414 68 418 72
rect 446 68 450 72
rect 486 68 490 72
rect 510 68 514 72
rect 382 58 386 62
rect 422 58 426 62
rect 518 58 522 62
rect 526 58 530 62
rect 566 58 570 62
rect 590 58 594 62
rect 630 58 634 62
rect 654 58 658 62
rect 758 108 762 112
rect 742 98 746 102
rect 766 98 770 102
rect 766 78 770 82
rect 798 78 802 82
rect 806 78 810 82
rect 782 68 786 72
rect 750 58 754 62
rect 790 58 794 62
rect 858 103 862 107
rect 865 103 869 107
rect 846 98 850 102
rect 830 88 834 92
rect 878 88 882 92
rect 830 78 834 82
rect 902 78 906 82
rect 942 88 946 92
rect 950 78 954 82
rect 998 118 1002 122
rect 1038 108 1042 112
rect 990 88 994 92
rect 1054 88 1058 92
rect 1014 78 1018 82
rect 1030 78 1034 82
rect 1070 78 1074 82
rect 1126 198 1130 202
rect 1174 228 1178 232
rect 1270 318 1274 322
rect 1334 318 1338 322
rect 1246 258 1250 262
rect 1318 308 1322 312
rect 1302 298 1306 302
rect 1310 278 1314 282
rect 1286 268 1290 272
rect 1334 268 1338 272
rect 1230 248 1234 252
rect 1262 248 1266 252
rect 1246 238 1250 242
rect 1214 228 1218 232
rect 1190 208 1194 212
rect 1102 148 1106 152
rect 1134 148 1138 152
rect 1190 148 1194 152
rect 1094 138 1098 142
rect 1126 138 1130 142
rect 1286 218 1290 222
rect 1270 188 1274 192
rect 1286 147 1290 151
rect 1166 138 1170 142
rect 1286 138 1290 142
rect 1190 128 1194 132
rect 1230 128 1234 132
rect 1166 118 1170 122
rect 1182 118 1186 122
rect 1238 118 1242 122
rect 1246 118 1250 122
rect 1142 108 1146 112
rect 1150 108 1154 112
rect 1094 88 1098 92
rect 1094 78 1098 82
rect 1134 78 1138 82
rect 974 68 978 72
rect 1014 68 1018 72
rect 1078 68 1082 72
rect 966 58 970 62
rect 990 58 994 62
rect 1038 58 1042 62
rect 1110 68 1114 72
rect 1134 68 1138 72
rect 1222 108 1226 112
rect 1430 318 1434 322
rect 1486 328 1490 332
rect 1582 368 1586 372
rect 1518 348 1522 352
rect 1534 348 1538 352
rect 1542 348 1546 352
rect 1566 338 1570 342
rect 1574 338 1578 342
rect 1542 328 1546 332
rect 1582 328 1586 332
rect 1646 458 1650 462
rect 1710 538 1714 542
rect 1702 528 1706 532
rect 1694 478 1698 482
rect 1702 468 1706 472
rect 1838 618 1842 622
rect 1950 628 1954 632
rect 1958 608 1962 612
rect 1950 598 1954 602
rect 1798 568 1802 572
rect 1830 568 1834 572
rect 1886 568 1890 572
rect 1814 558 1818 562
rect 1862 558 1866 562
rect 1846 548 1850 552
rect 1854 548 1858 552
rect 1886 548 1890 552
rect 1774 508 1778 512
rect 1734 488 1738 492
rect 1726 468 1730 472
rect 1702 458 1706 462
rect 1710 448 1714 452
rect 1726 448 1730 452
rect 1702 438 1706 442
rect 1742 438 1746 442
rect 1678 428 1682 432
rect 1654 408 1658 412
rect 1694 398 1698 402
rect 1622 378 1626 382
rect 1678 378 1682 382
rect 1654 348 1658 352
rect 1686 348 1690 352
rect 1606 338 1610 342
rect 1670 338 1674 342
rect 1686 338 1690 342
rect 1750 428 1754 432
rect 1838 478 1842 482
rect 1798 398 1802 402
rect 1814 398 1818 402
rect 1790 388 1794 392
rect 1742 378 1746 382
rect 1750 378 1754 382
rect 1710 348 1714 352
rect 1734 348 1738 352
rect 1766 348 1770 352
rect 1806 348 1810 352
rect 1702 338 1706 342
rect 1726 338 1730 342
rect 1598 328 1602 332
rect 1630 328 1634 332
rect 1510 318 1514 322
rect 1518 318 1522 322
rect 1590 318 1594 322
rect 1622 318 1626 322
rect 1470 308 1474 312
rect 1494 308 1498 312
rect 1414 288 1418 292
rect 1390 278 1394 282
rect 1422 278 1426 282
rect 1614 298 1618 302
rect 1638 318 1642 322
rect 1718 318 1722 322
rect 1758 338 1762 342
rect 1742 318 1746 322
rect 1710 288 1714 292
rect 1566 278 1570 282
rect 1606 278 1610 282
rect 1678 278 1682 282
rect 1542 268 1546 272
rect 1558 268 1562 272
rect 1342 238 1346 242
rect 1398 248 1402 252
rect 1398 238 1402 242
rect 1326 218 1330 222
rect 1358 218 1362 222
rect 1326 208 1330 212
rect 1370 203 1374 207
rect 1377 203 1381 207
rect 1462 258 1466 262
rect 1478 258 1482 262
rect 1446 238 1450 242
rect 1462 238 1466 242
rect 1406 218 1410 222
rect 1478 198 1482 202
rect 1390 188 1394 192
rect 1462 188 1466 192
rect 1350 178 1354 182
rect 1334 148 1338 152
rect 1390 138 1394 142
rect 1446 138 1450 142
rect 1414 128 1418 132
rect 1446 128 1450 132
rect 1874 503 1878 507
rect 1881 503 1885 507
rect 1878 488 1882 492
rect 1846 468 1850 472
rect 1854 468 1858 472
rect 1878 458 1882 462
rect 1854 418 1858 422
rect 1862 418 1866 422
rect 1886 418 1890 422
rect 1830 378 1834 382
rect 1846 378 1850 382
rect 1830 368 1834 372
rect 1854 348 1858 352
rect 1886 348 1890 352
rect 1822 338 1826 342
rect 1790 318 1794 322
rect 1838 318 1842 322
rect 1886 318 1890 322
rect 1758 308 1762 312
rect 1874 303 1878 307
rect 1881 303 1885 307
rect 1774 288 1778 292
rect 1750 278 1754 282
rect 1574 268 1578 272
rect 1590 268 1594 272
rect 1606 268 1610 272
rect 1614 268 1618 272
rect 1686 268 1690 272
rect 1702 268 1706 272
rect 1574 248 1578 252
rect 1526 238 1530 242
rect 1558 238 1562 242
rect 1494 218 1498 222
rect 1582 238 1586 242
rect 1558 188 1562 192
rect 1486 158 1490 162
rect 1494 158 1498 162
rect 1462 138 1466 142
rect 1406 118 1410 122
rect 1454 118 1458 122
rect 1662 258 1666 262
rect 1942 578 1946 582
rect 1926 558 1930 562
rect 1918 548 1922 552
rect 2014 858 2018 862
rect 2006 848 2010 852
rect 2070 918 2074 922
rect 2094 908 2098 912
rect 2054 898 2058 902
rect 2134 898 2138 902
rect 2278 1018 2282 1022
rect 2230 968 2234 972
rect 2278 948 2282 952
rect 2214 938 2218 942
rect 2262 938 2266 942
rect 2110 888 2114 892
rect 2190 888 2194 892
rect 2262 918 2266 922
rect 2182 878 2186 882
rect 2214 878 2218 882
rect 2222 878 2226 882
rect 2294 898 2298 902
rect 2550 1328 2554 1332
rect 2574 1318 2578 1322
rect 2342 1308 2346 1312
rect 2382 1308 2386 1312
rect 2470 1308 2474 1312
rect 2334 1298 2338 1302
rect 2326 1278 2330 1282
rect 2366 1288 2370 1292
rect 2342 1218 2346 1222
rect 2390 1258 2394 1262
rect 2406 1248 2410 1252
rect 2454 1248 2458 1252
rect 2394 1203 2398 1207
rect 2401 1203 2405 1207
rect 2478 1288 2482 1292
rect 2494 1268 2498 1272
rect 2422 1178 2426 1182
rect 2470 1178 2474 1182
rect 2326 1168 2330 1172
rect 2446 1168 2450 1172
rect 2478 1168 2482 1172
rect 2342 1148 2346 1152
rect 2438 1148 2442 1152
rect 2454 1128 2458 1132
rect 2662 1328 2666 1332
rect 2710 1328 2714 1332
rect 2630 1318 2634 1322
rect 2654 1318 2658 1322
rect 2598 1298 2602 1302
rect 2630 1298 2634 1302
rect 2694 1288 2698 1292
rect 2670 1268 2674 1272
rect 2614 1258 2618 1262
rect 2558 1248 2562 1252
rect 2638 1248 2642 1252
rect 2526 1238 2530 1242
rect 2518 1218 2522 1222
rect 2670 1248 2674 1252
rect 2694 1228 2698 1232
rect 2662 1208 2666 1212
rect 2678 1208 2682 1212
rect 2502 1158 2506 1162
rect 2566 1158 2570 1162
rect 2606 1158 2610 1162
rect 2622 1158 2626 1162
rect 2486 1138 2490 1142
rect 2502 1128 2506 1132
rect 2326 1118 2330 1122
rect 2398 1118 2402 1122
rect 2454 1118 2458 1122
rect 2478 1118 2482 1122
rect 2382 1108 2386 1112
rect 2366 1098 2370 1102
rect 2614 1138 2618 1142
rect 2630 1138 2634 1142
rect 2646 1138 2650 1142
rect 2574 1098 2578 1102
rect 2606 1128 2610 1132
rect 2630 1128 2634 1132
rect 2638 1118 2642 1122
rect 2670 1118 2674 1122
rect 2670 1108 2674 1112
rect 2558 1078 2562 1082
rect 2598 1078 2602 1082
rect 2622 1078 2626 1082
rect 2350 1068 2354 1072
rect 2358 1068 2362 1072
rect 2494 1068 2498 1072
rect 2526 1068 2530 1072
rect 2342 1058 2346 1062
rect 2382 1058 2386 1062
rect 2438 1058 2442 1062
rect 2478 1058 2482 1062
rect 2502 1058 2506 1062
rect 2542 1058 2546 1062
rect 2350 1038 2354 1042
rect 2326 1018 2330 1022
rect 2318 998 2322 1002
rect 2318 988 2322 992
rect 2462 1038 2466 1042
rect 2358 1018 2362 1022
rect 2358 1008 2362 1012
rect 2394 1003 2398 1007
rect 2401 1003 2405 1007
rect 2494 1018 2498 1022
rect 2518 1018 2522 1022
rect 2478 978 2482 982
rect 2342 968 2346 972
rect 2366 968 2370 972
rect 2374 968 2378 972
rect 2654 1058 2658 1062
rect 2574 1048 2578 1052
rect 2606 1048 2610 1052
rect 2550 1038 2554 1042
rect 2582 1018 2586 1022
rect 2326 958 2330 962
rect 2390 958 2394 962
rect 2462 958 2466 962
rect 2494 958 2498 962
rect 2342 938 2346 942
rect 2358 938 2362 942
rect 2358 908 2362 912
rect 2414 938 2418 942
rect 2430 938 2434 942
rect 2542 948 2546 952
rect 2558 948 2562 952
rect 2606 948 2610 952
rect 2494 938 2498 942
rect 2518 938 2522 942
rect 2542 938 2546 942
rect 2438 928 2442 932
rect 2366 898 2370 902
rect 2406 898 2410 902
rect 2030 868 2034 872
rect 2166 868 2170 872
rect 2182 868 2186 872
rect 2294 868 2298 872
rect 2366 868 2370 872
rect 2094 858 2098 862
rect 2126 858 2130 862
rect 2142 858 2146 862
rect 2038 848 2042 852
rect 2046 848 2050 852
rect 2038 828 2042 832
rect 2006 798 2010 802
rect 2022 798 2026 802
rect 2150 848 2154 852
rect 2214 858 2218 862
rect 2254 858 2258 862
rect 2166 848 2170 852
rect 2142 838 2146 842
rect 2158 838 2162 842
rect 2270 838 2274 842
rect 2286 838 2290 842
rect 2270 818 2274 822
rect 2222 808 2226 812
rect 2038 768 2042 772
rect 2134 768 2138 772
rect 2078 758 2082 762
rect 2110 758 2114 762
rect 2086 748 2090 752
rect 2182 748 2186 752
rect 2206 748 2210 752
rect 2070 728 2074 732
rect 2110 728 2114 732
rect 2158 728 2162 732
rect 2182 728 2186 732
rect 2030 688 2034 692
rect 2150 718 2154 722
rect 2214 718 2218 722
rect 2182 708 2186 712
rect 2174 698 2178 702
rect 2102 688 2106 692
rect 2078 678 2082 682
rect 2062 638 2066 642
rect 2006 598 2010 602
rect 1982 578 1986 582
rect 1974 568 1978 572
rect 1958 558 1962 562
rect 2134 658 2138 662
rect 2102 608 2106 612
rect 2126 608 2130 612
rect 2070 558 2074 562
rect 2086 558 2090 562
rect 1974 548 1978 552
rect 1926 528 1930 532
rect 1950 527 1954 531
rect 1982 528 1986 532
rect 2022 528 2026 532
rect 1942 518 1946 522
rect 1982 518 1986 522
rect 1918 478 1922 482
rect 1934 478 1938 482
rect 1974 468 1978 472
rect 1998 498 2002 502
rect 1990 478 1994 482
rect 2014 478 2018 482
rect 2118 598 2122 602
rect 2174 568 2178 572
rect 2070 478 2074 482
rect 2390 858 2394 862
rect 2414 878 2418 882
rect 2470 928 2474 932
rect 2486 928 2490 932
rect 2462 918 2466 922
rect 2430 898 2434 902
rect 2446 878 2450 882
rect 2686 1168 2690 1172
rect 2702 1208 2706 1212
rect 2718 1278 2722 1282
rect 2718 1258 2722 1262
rect 2686 1138 2690 1142
rect 2822 1338 2826 1342
rect 2766 1328 2770 1332
rect 2774 1298 2778 1302
rect 2806 1328 2810 1332
rect 2830 1328 2834 1332
rect 2798 1298 2802 1302
rect 2782 1288 2786 1292
rect 2822 1278 2826 1282
rect 2758 1268 2762 1272
rect 2782 1268 2786 1272
rect 2750 1258 2754 1262
rect 2750 1238 2754 1242
rect 2790 1258 2794 1262
rect 2814 1258 2818 1262
rect 2982 1398 2986 1402
rect 2934 1358 2938 1362
rect 2942 1358 2946 1362
rect 2910 1328 2914 1332
rect 2942 1328 2946 1332
rect 2990 1328 2994 1332
rect 3062 1378 3066 1382
rect 3102 1378 3106 1382
rect 3142 1378 3146 1382
rect 3182 1448 3186 1452
rect 3302 1548 3306 1552
rect 3310 1538 3314 1542
rect 3310 1498 3314 1502
rect 3502 1718 3506 1722
rect 3478 1688 3482 1692
rect 3438 1668 3442 1672
rect 3462 1658 3466 1662
rect 3478 1658 3482 1662
rect 3526 1698 3530 1702
rect 3526 1688 3530 1692
rect 3510 1658 3514 1662
rect 3446 1648 3450 1652
rect 3486 1648 3490 1652
rect 3510 1648 3514 1652
rect 3518 1648 3522 1652
rect 3550 1728 3554 1732
rect 3614 1748 3618 1752
rect 3606 1698 3610 1702
rect 3662 1688 3666 1692
rect 3598 1678 3602 1682
rect 3662 1678 3666 1682
rect 3550 1658 3554 1662
rect 3382 1638 3386 1642
rect 3494 1638 3498 1642
rect 3398 1608 3402 1612
rect 3406 1608 3410 1612
rect 3342 1558 3346 1562
rect 3366 1558 3370 1562
rect 3342 1548 3346 1552
rect 3358 1538 3362 1542
rect 3390 1538 3394 1542
rect 3358 1528 3362 1532
rect 3350 1508 3354 1512
rect 3390 1488 3394 1492
rect 3334 1478 3338 1482
rect 3342 1478 3346 1482
rect 3382 1478 3386 1482
rect 3326 1448 3330 1452
rect 3230 1438 3234 1442
rect 3294 1438 3298 1442
rect 3190 1428 3194 1432
rect 3214 1428 3218 1432
rect 3190 1388 3194 1392
rect 3318 1388 3322 1392
rect 3246 1358 3250 1362
rect 3030 1348 3034 1352
rect 3150 1348 3154 1352
rect 3054 1338 3058 1342
rect 3094 1338 3098 1342
rect 3118 1338 3122 1342
rect 3174 1338 3178 1342
rect 3006 1328 3010 1332
rect 3014 1318 3018 1322
rect 2974 1308 2978 1312
rect 2998 1308 3002 1312
rect 2906 1303 2910 1307
rect 2913 1303 2917 1307
rect 2886 1298 2890 1302
rect 2862 1288 2866 1292
rect 2958 1278 2962 1282
rect 2846 1248 2850 1252
rect 2878 1268 2882 1272
rect 2910 1268 2914 1272
rect 2886 1258 2890 1262
rect 2902 1258 2906 1262
rect 2942 1258 2946 1262
rect 2886 1238 2890 1242
rect 2838 1228 2842 1232
rect 2854 1228 2858 1232
rect 2774 1218 2778 1222
rect 2782 1218 2786 1222
rect 2758 1208 2762 1212
rect 2774 1208 2778 1212
rect 2734 1168 2738 1172
rect 2710 1138 2714 1142
rect 2702 1128 2706 1132
rect 2718 1128 2722 1132
rect 2966 1268 2970 1272
rect 2982 1278 2986 1282
rect 3038 1268 3042 1272
rect 3054 1268 3058 1272
rect 3006 1258 3010 1262
rect 3022 1258 3026 1262
rect 3046 1258 3050 1262
rect 3102 1288 3106 1292
rect 3070 1268 3074 1272
rect 3094 1258 3098 1262
rect 3158 1268 3162 1272
rect 3158 1258 3162 1262
rect 2950 1248 2954 1252
rect 2974 1248 2978 1252
rect 3030 1248 3034 1252
rect 3062 1248 3066 1252
rect 2918 1208 2922 1212
rect 2902 1168 2906 1172
rect 2966 1168 2970 1172
rect 2822 1158 2826 1162
rect 2734 1138 2738 1142
rect 2766 1138 2770 1142
rect 2958 1158 2962 1162
rect 2750 1128 2754 1132
rect 2726 1118 2730 1122
rect 2838 1108 2842 1112
rect 2862 1118 2866 1122
rect 2870 1108 2874 1112
rect 2910 1128 2914 1132
rect 2934 1128 2938 1132
rect 2906 1103 2910 1107
rect 2913 1103 2917 1107
rect 2774 1078 2778 1082
rect 2806 1078 2810 1082
rect 2854 1078 2858 1082
rect 2886 1078 2890 1082
rect 2926 1078 2930 1082
rect 2686 1066 2690 1070
rect 2734 1068 2738 1072
rect 2742 1068 2746 1072
rect 2750 1058 2754 1062
rect 2662 1048 2666 1052
rect 2702 1048 2706 1052
rect 2742 1048 2746 1052
rect 2646 1038 2650 1042
rect 2782 1068 2786 1072
rect 2766 1038 2770 1042
rect 2814 1068 2818 1072
rect 2838 1058 2842 1062
rect 2854 1058 2858 1062
rect 2886 1058 2890 1062
rect 2918 1058 2922 1062
rect 2838 1048 2842 1052
rect 2854 1048 2858 1052
rect 2886 1048 2890 1052
rect 2798 1038 2802 1042
rect 2814 1038 2818 1042
rect 2790 1018 2794 1022
rect 2742 998 2746 1002
rect 2862 1018 2866 1022
rect 2734 988 2738 992
rect 2798 968 2802 972
rect 2870 968 2874 972
rect 2678 958 2682 962
rect 2654 948 2658 952
rect 2710 948 2714 952
rect 2822 938 2826 942
rect 2614 928 2618 932
rect 2622 928 2626 932
rect 2758 928 2762 932
rect 2606 918 2610 922
rect 2582 908 2586 912
rect 2742 908 2746 912
rect 2582 898 2586 902
rect 2614 898 2618 902
rect 2726 888 2730 892
rect 2558 878 2562 882
rect 2566 878 2570 882
rect 2638 878 2642 882
rect 2646 878 2650 882
rect 2494 868 2498 872
rect 2518 868 2522 872
rect 2542 868 2546 872
rect 2862 918 2866 922
rect 2870 918 2874 922
rect 2774 888 2778 892
rect 2830 878 2834 882
rect 2582 868 2586 872
rect 2710 868 2714 872
rect 2830 868 2834 872
rect 2422 858 2426 862
rect 2438 858 2442 862
rect 2462 858 2466 862
rect 2566 858 2570 862
rect 2334 848 2338 852
rect 2422 848 2426 852
rect 2454 848 2458 852
rect 2526 848 2530 852
rect 2790 848 2794 852
rect 2310 838 2314 842
rect 2414 838 2418 842
rect 2766 828 2770 832
rect 2294 818 2298 822
rect 2358 818 2362 822
rect 2614 818 2618 822
rect 2394 803 2398 807
rect 2401 803 2405 807
rect 2294 778 2298 782
rect 2502 778 2506 782
rect 2286 768 2290 772
rect 2326 768 2330 772
rect 2478 768 2482 772
rect 2670 768 2674 772
rect 2814 838 2818 842
rect 2942 1068 2946 1072
rect 2974 1128 2978 1132
rect 3102 1238 3106 1242
rect 2998 1228 3002 1232
rect 3006 1228 3010 1232
rect 3054 1218 3058 1222
rect 3006 1208 3010 1212
rect 3198 1328 3202 1332
rect 3230 1328 3234 1332
rect 3230 1278 3234 1282
rect 3262 1288 3266 1292
rect 3294 1268 3298 1272
rect 3246 1258 3250 1262
rect 3182 1198 3186 1202
rect 3198 1188 3202 1192
rect 2990 1178 2994 1182
rect 2998 1168 3002 1172
rect 2990 1158 2994 1162
rect 3198 1158 3202 1162
rect 2982 1118 2986 1122
rect 2998 1118 3002 1122
rect 2966 1078 2970 1082
rect 2950 1058 2954 1062
rect 2934 1038 2938 1042
rect 2958 978 2962 982
rect 2990 968 2994 972
rect 2974 948 2978 952
rect 2966 908 2970 912
rect 2906 903 2910 907
rect 2913 903 2917 907
rect 3086 1138 3090 1142
rect 3134 1138 3138 1142
rect 3062 1118 3066 1122
rect 3006 928 3010 932
rect 2894 888 2898 892
rect 3102 1038 3106 1042
rect 3182 1088 3186 1092
rect 3150 1078 3154 1082
rect 3158 1058 3162 1062
rect 3310 1088 3314 1092
rect 3310 1078 3314 1082
rect 3214 1068 3218 1072
rect 3350 1438 3354 1442
rect 3418 1603 3422 1607
rect 3425 1603 3429 1607
rect 3422 1548 3426 1552
rect 3414 1538 3418 1542
rect 3462 1538 3466 1542
rect 3414 1508 3418 1512
rect 3406 1468 3410 1472
rect 3382 1438 3386 1442
rect 3366 1418 3370 1422
rect 3366 1318 3370 1322
rect 3454 1438 3458 1442
rect 3502 1508 3506 1512
rect 3494 1488 3498 1492
rect 3478 1468 3482 1472
rect 3462 1428 3466 1432
rect 3470 1428 3474 1432
rect 3494 1428 3498 1432
rect 3418 1403 3422 1407
rect 3425 1403 3429 1407
rect 3574 1658 3578 1662
rect 3638 1668 3642 1672
rect 3566 1648 3570 1652
rect 3590 1648 3594 1652
rect 3614 1648 3618 1652
rect 3558 1638 3562 1642
rect 3582 1638 3586 1642
rect 3566 1628 3570 1632
rect 3518 1548 3522 1552
rect 3550 1498 3554 1502
rect 3934 1878 3938 1882
rect 3806 1868 3810 1872
rect 3718 1858 3722 1862
rect 3742 1858 3746 1862
rect 3854 1858 3858 1862
rect 3718 1838 3722 1842
rect 3870 1818 3874 1822
rect 3758 1758 3762 1762
rect 3790 1758 3794 1762
rect 3894 1758 3898 1762
rect 3718 1748 3722 1752
rect 3726 1748 3730 1752
rect 3718 1738 3722 1742
rect 3678 1718 3682 1722
rect 3694 1708 3698 1712
rect 3710 1698 3714 1702
rect 3734 1718 3738 1722
rect 3718 1688 3722 1692
rect 3750 1748 3754 1752
rect 3758 1738 3762 1742
rect 3782 1748 3786 1752
rect 3862 1748 3866 1752
rect 3806 1738 3810 1742
rect 4006 2098 4010 2102
rect 4022 2088 4026 2092
rect 4070 2098 4074 2102
rect 4062 2078 4066 2082
rect 4102 2078 4106 2082
rect 4062 2068 4066 2072
rect 3990 2058 3994 2062
rect 4094 2058 4098 2062
rect 3982 2038 3986 2042
rect 4070 1988 4074 1992
rect 4022 1968 4026 1972
rect 3974 1958 3978 1962
rect 4006 1958 4010 1962
rect 4038 1958 4042 1962
rect 4054 1958 4058 1962
rect 4030 1948 4034 1952
rect 4046 1938 4050 1942
rect 4062 1948 4066 1952
rect 3974 1928 3978 1932
rect 3982 1898 3986 1902
rect 4078 1968 4082 1972
rect 4118 2058 4122 2062
rect 4142 2058 4146 2062
rect 4134 2048 4138 2052
rect 4102 2038 4106 2042
rect 4118 2018 4122 2022
rect 4222 2258 4226 2262
rect 4222 2248 4226 2252
rect 4270 2248 4274 2252
rect 4214 2238 4218 2242
rect 4190 2218 4194 2222
rect 4350 2358 4354 2362
rect 4310 2288 4314 2292
rect 4334 2288 4338 2292
rect 4350 2288 4354 2292
rect 4326 2278 4330 2282
rect 4342 2278 4346 2282
rect 4334 2268 4338 2272
rect 4302 2258 4306 2262
rect 4310 2258 4314 2262
rect 4294 2238 4298 2242
rect 4278 2228 4282 2232
rect 4270 2208 4274 2212
rect 4254 2198 4258 2202
rect 4230 2178 4234 2182
rect 4262 2178 4266 2182
rect 4278 2178 4282 2182
rect 4238 2168 4242 2172
rect 4254 2168 4258 2172
rect 4214 2158 4218 2162
rect 4222 2158 4226 2162
rect 4246 2148 4250 2152
rect 4278 2148 4282 2152
rect 4206 2128 4210 2132
rect 4158 2108 4162 2112
rect 4310 2238 4314 2242
rect 4294 2218 4298 2222
rect 4302 2218 4306 2222
rect 4294 2188 4298 2192
rect 4582 2478 4586 2482
rect 4598 2478 4602 2482
rect 4638 2478 4642 2482
rect 4590 2468 4594 2472
rect 4614 2468 4618 2472
rect 4566 2458 4570 2462
rect 4598 2458 4602 2462
rect 4638 2458 4642 2462
rect 4630 2448 4634 2452
rect 4534 2438 4538 2442
rect 4558 2438 4562 2442
rect 4398 2418 4402 2422
rect 4442 2403 4446 2407
rect 4449 2403 4453 2407
rect 4542 2378 4546 2382
rect 4494 2368 4498 2372
rect 4534 2368 4538 2372
rect 4366 2358 4370 2362
rect 4398 2358 4402 2362
rect 4422 2338 4426 2342
rect 4470 2338 4474 2342
rect 4470 2328 4474 2332
rect 4510 2328 4514 2332
rect 4574 2358 4578 2362
rect 4582 2358 4586 2362
rect 4662 2578 4666 2582
rect 4670 2568 4674 2572
rect 4670 2558 4674 2562
rect 4710 2558 4714 2562
rect 4686 2548 4690 2552
rect 4678 2538 4682 2542
rect 4798 2598 4802 2602
rect 4758 2588 4762 2592
rect 4790 2538 4794 2542
rect 4702 2528 4706 2532
rect 4742 2528 4746 2532
rect 4702 2498 4706 2502
rect 4734 2508 4738 2512
rect 4662 2478 4666 2482
rect 4726 2478 4730 2482
rect 4670 2468 4674 2472
rect 4678 2468 4682 2472
rect 4766 2518 4770 2522
rect 4790 2498 4794 2502
rect 4766 2488 4770 2492
rect 4846 2598 4850 2602
rect 4862 2558 4866 2562
rect 5038 2868 5042 2872
rect 5118 2918 5122 2922
rect 5126 2918 5130 2922
rect 5062 2858 5066 2862
rect 4942 2848 4946 2852
rect 4950 2848 4954 2852
rect 4998 2848 5002 2852
rect 5022 2848 5026 2852
rect 5046 2838 5050 2842
rect 4990 2768 4994 2772
rect 5006 2748 5010 2752
rect 5022 2748 5026 2752
rect 4966 2738 4970 2742
rect 4942 2728 4946 2732
rect 5006 2728 5010 2732
rect 5022 2728 5026 2732
rect 4974 2718 4978 2722
rect 4954 2703 4958 2707
rect 4961 2703 4965 2707
rect 4910 2668 4914 2672
rect 4894 2648 4898 2652
rect 4910 2648 4914 2652
rect 4894 2638 4898 2642
rect 4902 2618 4906 2622
rect 4886 2608 4890 2612
rect 5030 2718 5034 2722
rect 5006 2698 5010 2702
rect 5006 2688 5010 2692
rect 4990 2668 4994 2672
rect 4998 2648 5002 2652
rect 5086 2758 5090 2762
rect 5070 2738 5074 2742
rect 5038 2688 5042 2692
rect 5046 2688 5050 2692
rect 5038 2678 5042 2682
rect 5070 2678 5074 2682
rect 5046 2668 5050 2672
rect 5054 2668 5058 2672
rect 5094 2748 5098 2752
rect 5182 2928 5186 2932
rect 5174 2868 5178 2872
rect 5230 2908 5234 2912
rect 5262 3078 5266 3082
rect 5270 3078 5274 3082
rect 5278 3058 5282 3062
rect 5270 3048 5274 3052
rect 5286 3028 5290 3032
rect 5262 3018 5266 3022
rect 5294 3018 5298 3022
rect 5286 2948 5290 2952
rect 5294 2938 5298 2942
rect 5262 2928 5266 2932
rect 5254 2918 5258 2922
rect 5270 2918 5274 2922
rect 5222 2868 5226 2872
rect 5222 2828 5226 2832
rect 5214 2758 5218 2762
rect 5134 2698 5138 2702
rect 5142 2688 5146 2692
rect 5182 2668 5186 2672
rect 5070 2648 5074 2652
rect 5190 2658 5194 2662
rect 5126 2648 5130 2652
rect 5022 2638 5026 2642
rect 5030 2638 5034 2642
rect 5054 2638 5058 2642
rect 5110 2638 5114 2642
rect 5134 2638 5138 2642
rect 5190 2638 5194 2642
rect 5286 2908 5290 2912
rect 5310 3068 5314 3072
rect 5310 3048 5314 3052
rect 5310 2968 5314 2972
rect 5310 2948 5314 2952
rect 5302 2898 5306 2902
rect 5358 2898 5362 2902
rect 5286 2848 5290 2852
rect 5278 2768 5282 2772
rect 5270 2758 5274 2762
rect 5254 2738 5258 2742
rect 5302 2738 5306 2742
rect 5262 2688 5266 2692
rect 4990 2628 4994 2632
rect 5158 2628 5162 2632
rect 5230 2628 5234 2632
rect 4982 2598 4986 2602
rect 4886 2568 4890 2572
rect 4942 2568 4946 2572
rect 4982 2568 4986 2572
rect 4998 2568 5002 2572
rect 4894 2558 4898 2562
rect 4934 2558 4938 2562
rect 4830 2548 4834 2552
rect 4846 2548 4850 2552
rect 4870 2548 4874 2552
rect 4814 2538 4818 2542
rect 4822 2538 4826 2542
rect 4838 2538 4842 2542
rect 4806 2498 4810 2502
rect 4814 2488 4818 2492
rect 4782 2468 4786 2472
rect 4814 2468 4818 2472
rect 5238 2608 5242 2612
rect 5102 2578 5106 2582
rect 4966 2558 4970 2562
rect 5022 2558 5026 2562
rect 5094 2558 5098 2562
rect 4990 2548 4994 2552
rect 4934 2538 4938 2542
rect 5014 2538 5018 2542
rect 4870 2528 4874 2532
rect 4926 2518 4930 2522
rect 4982 2518 4986 2522
rect 4854 2478 4858 2482
rect 4878 2508 4882 2512
rect 4894 2478 4898 2482
rect 4886 2468 4890 2472
rect 4694 2458 4698 2462
rect 4758 2458 4762 2462
rect 4766 2458 4770 2462
rect 4830 2458 4834 2462
rect 4954 2503 4958 2507
rect 4961 2503 4965 2507
rect 4934 2478 4938 2482
rect 5022 2528 5026 2532
rect 5022 2508 5026 2512
rect 5134 2568 5138 2572
rect 5198 2568 5202 2572
rect 5182 2548 5186 2552
rect 5254 2548 5258 2552
rect 5102 2518 5106 2522
rect 5102 2508 5106 2512
rect 5094 2498 5098 2502
rect 5038 2478 5042 2482
rect 5078 2478 5082 2482
rect 5278 2698 5282 2702
rect 5270 2638 5274 2642
rect 5270 2608 5274 2612
rect 5158 2528 5162 2532
rect 5246 2528 5250 2532
rect 5262 2528 5266 2532
rect 5110 2488 5114 2492
rect 5158 2478 5162 2482
rect 4918 2468 4922 2472
rect 4958 2468 4962 2472
rect 5038 2468 5042 2472
rect 5094 2468 5098 2472
rect 5126 2468 5130 2472
rect 5030 2458 5034 2462
rect 5054 2458 5058 2462
rect 5086 2458 5090 2462
rect 5102 2458 5106 2462
rect 5150 2458 5154 2462
rect 4726 2448 4730 2452
rect 4750 2448 4754 2452
rect 5078 2448 5082 2452
rect 5142 2448 5146 2452
rect 5150 2448 5154 2452
rect 4686 2388 4690 2392
rect 4670 2378 4674 2382
rect 4758 2378 4762 2382
rect 4766 2378 4770 2382
rect 4734 2368 4738 2372
rect 4750 2368 4754 2372
rect 4734 2358 4738 2362
rect 4766 2358 4770 2362
rect 4790 2358 4794 2362
rect 4822 2358 4826 2362
rect 4566 2338 4570 2342
rect 4590 2338 4594 2342
rect 4654 2338 4658 2342
rect 4550 2328 4554 2332
rect 4574 2328 4578 2332
rect 4462 2318 4466 2322
rect 4502 2318 4506 2322
rect 4518 2318 4522 2322
rect 4526 2318 4530 2322
rect 4366 2288 4370 2292
rect 4398 2278 4402 2282
rect 4470 2278 4474 2282
rect 4718 2338 4722 2342
rect 5062 2438 5066 2442
rect 5078 2438 5082 2442
rect 5094 2438 5098 2442
rect 5110 2438 5114 2442
rect 5054 2418 5058 2422
rect 4910 2378 4914 2382
rect 4918 2368 4922 2372
rect 4958 2368 4962 2372
rect 4822 2348 4826 2352
rect 4846 2348 4850 2352
rect 4862 2348 4866 2352
rect 4886 2348 4890 2352
rect 4894 2348 4898 2352
rect 4798 2338 4802 2342
rect 4814 2338 4818 2342
rect 4830 2338 4834 2342
rect 4846 2338 4850 2342
rect 4902 2338 4906 2342
rect 4982 2338 4986 2342
rect 4678 2328 4682 2332
rect 4742 2328 4746 2332
rect 4790 2328 4794 2332
rect 4542 2308 4546 2312
rect 4614 2308 4618 2312
rect 4590 2298 4594 2302
rect 4526 2288 4530 2292
rect 4574 2288 4578 2292
rect 4550 2278 4554 2282
rect 4374 2268 4378 2272
rect 4430 2268 4434 2272
rect 4486 2268 4490 2272
rect 4406 2258 4410 2262
rect 4422 2258 4426 2262
rect 4502 2258 4506 2262
rect 4414 2248 4418 2252
rect 4534 2268 4538 2272
rect 4390 2238 4394 2242
rect 4446 2238 4450 2242
rect 4398 2228 4402 2232
rect 4430 2218 4434 2222
rect 4422 2198 4426 2202
rect 4310 2168 4314 2172
rect 4342 2168 4346 2172
rect 4302 2158 4306 2162
rect 4334 2158 4338 2162
rect 4294 2148 4298 2152
rect 4414 2148 4418 2152
rect 4310 2108 4314 2112
rect 4350 2118 4354 2122
rect 4414 2118 4418 2122
rect 4342 2108 4346 2112
rect 4334 2098 4338 2102
rect 4442 2203 4446 2207
rect 4449 2203 4453 2207
rect 4638 2288 4642 2292
rect 4686 2318 4690 2322
rect 4654 2278 4658 2282
rect 4934 2328 4938 2332
rect 4838 2318 4842 2322
rect 4694 2288 4698 2292
rect 4774 2288 4778 2292
rect 4686 2278 4690 2282
rect 4742 2278 4746 2282
rect 4758 2278 4762 2282
rect 4670 2268 4674 2272
rect 4734 2268 4738 2272
rect 4766 2268 4770 2272
rect 4566 2258 4570 2262
rect 4638 2258 4642 2262
rect 4718 2258 4722 2262
rect 4574 2248 4578 2252
rect 4590 2248 4594 2252
rect 4526 2228 4530 2232
rect 4558 2228 4562 2232
rect 4606 2238 4610 2242
rect 4854 2278 4858 2282
rect 4910 2278 4914 2282
rect 4954 2303 4958 2307
rect 4961 2303 4965 2307
rect 5046 2398 5050 2402
rect 5022 2368 5026 2372
rect 5062 2378 5066 2382
rect 5102 2378 5106 2382
rect 5078 2368 5082 2372
rect 5006 2358 5010 2362
rect 5014 2358 5018 2362
rect 5062 2358 5066 2362
rect 5046 2348 5050 2352
rect 5070 2348 5074 2352
rect 5086 2348 5090 2352
rect 5102 2348 5106 2352
rect 5022 2338 5026 2342
rect 4990 2298 4994 2302
rect 4982 2278 4986 2282
rect 5094 2338 5098 2342
rect 5062 2308 5066 2312
rect 5086 2298 5090 2302
rect 5046 2288 5050 2292
rect 5022 2278 5026 2282
rect 4942 2268 4946 2272
rect 4966 2268 4970 2272
rect 4798 2258 4802 2262
rect 4846 2258 4850 2262
rect 4902 2258 4906 2262
rect 4926 2258 4930 2262
rect 5134 2398 5138 2402
rect 5126 2368 5130 2372
rect 5118 2338 5122 2342
rect 5150 2358 5154 2362
rect 5270 2518 5274 2522
rect 5174 2508 5178 2512
rect 5206 2508 5210 2512
rect 5182 2478 5186 2482
rect 5262 2508 5266 2512
rect 5270 2508 5274 2512
rect 5214 2498 5218 2502
rect 5214 2478 5218 2482
rect 5190 2458 5194 2462
rect 5206 2408 5210 2412
rect 5182 2398 5186 2402
rect 5214 2388 5218 2392
rect 5190 2358 5194 2362
rect 5182 2338 5186 2342
rect 5190 2328 5194 2332
rect 5166 2318 5170 2322
rect 5134 2308 5138 2312
rect 5174 2308 5178 2312
rect 5126 2298 5130 2302
rect 5166 2298 5170 2302
rect 5110 2288 5114 2292
rect 5150 2278 5154 2282
rect 5214 2338 5218 2342
rect 5222 2328 5226 2332
rect 5294 2678 5298 2682
rect 5286 2668 5290 2672
rect 5302 2658 5306 2662
rect 5286 2558 5290 2562
rect 5286 2538 5290 2542
rect 5310 2538 5314 2542
rect 5294 2518 5298 2522
rect 5302 2478 5306 2482
rect 5286 2458 5290 2462
rect 5286 2348 5290 2352
rect 5278 2338 5282 2342
rect 5294 2338 5298 2342
rect 5206 2288 5210 2292
rect 5246 2278 5250 2282
rect 5062 2268 5066 2272
rect 5134 2268 5138 2272
rect 5174 2268 5178 2272
rect 5222 2268 5226 2272
rect 4998 2258 5002 2262
rect 5006 2258 5010 2262
rect 4750 2248 4754 2252
rect 4886 2248 4890 2252
rect 4998 2248 5002 2252
rect 4774 2238 4778 2242
rect 4598 2228 4602 2232
rect 4622 2228 4626 2232
rect 4734 2198 4738 2202
rect 4638 2188 4642 2192
rect 4726 2188 4730 2192
rect 4502 2168 4506 2172
rect 4550 2168 4554 2172
rect 4598 2168 4602 2172
rect 4630 2168 4634 2172
rect 4566 2158 4570 2162
rect 4438 2148 4442 2152
rect 4526 2148 4530 2152
rect 4438 2128 4442 2132
rect 4470 2128 4474 2132
rect 4550 2148 4554 2152
rect 4590 2158 4594 2162
rect 4582 2148 4586 2152
rect 4598 2148 4602 2152
rect 4654 2178 4658 2182
rect 4678 2178 4682 2182
rect 4662 2158 4666 2162
rect 4718 2148 4722 2152
rect 4606 2138 4610 2142
rect 4614 2138 4618 2142
rect 4646 2138 4650 2142
rect 4686 2138 4690 2142
rect 4558 2128 4562 2132
rect 4606 2128 4610 2132
rect 4542 2118 4546 2122
rect 4622 2118 4626 2122
rect 4486 2108 4490 2112
rect 4518 2108 4522 2112
rect 4734 2158 4738 2162
rect 4766 2158 4770 2162
rect 4758 2148 4762 2152
rect 4862 2188 4866 2192
rect 4790 2178 4794 2182
rect 4830 2168 4834 2172
rect 4870 2178 4874 2182
rect 4790 2148 4794 2152
rect 4902 2158 4906 2162
rect 5086 2248 5090 2252
rect 5030 2238 5034 2242
rect 5062 2238 5066 2242
rect 4990 2208 4994 2212
rect 4934 2188 4938 2192
rect 4950 2178 4954 2182
rect 4982 2168 4986 2172
rect 5078 2168 5082 2172
rect 4926 2158 4930 2162
rect 5022 2158 5026 2162
rect 5030 2158 5034 2162
rect 4966 2148 4970 2152
rect 4822 2138 4826 2142
rect 4846 2138 4850 2142
rect 4926 2138 4930 2142
rect 4950 2138 4954 2142
rect 4742 2128 4746 2132
rect 4694 2118 4698 2122
rect 4702 2118 4706 2122
rect 4750 2118 4754 2122
rect 4174 2078 4178 2082
rect 4198 2078 4202 2082
rect 4422 2078 4426 2082
rect 4550 2078 4554 2082
rect 4598 2078 4602 2082
rect 4166 2058 4170 2062
rect 4230 2068 4234 2072
rect 4246 2058 4250 2062
rect 4214 2048 4218 2052
rect 4222 2048 4226 2052
rect 4790 2098 4794 2102
rect 4654 2088 4658 2092
rect 4686 2088 4690 2092
rect 4854 2088 4858 2092
rect 4902 2128 4906 2132
rect 4886 2078 4890 2082
rect 4270 2068 4274 2072
rect 4486 2068 4490 2072
rect 4774 2068 4778 2072
rect 4334 2058 4338 2062
rect 4254 2038 4258 2042
rect 4278 2038 4282 2042
rect 4166 2028 4170 2032
rect 4270 1998 4274 2002
rect 4150 1978 4154 1982
rect 4118 1958 4122 1962
rect 4182 1948 4186 1952
rect 4542 2058 4546 2062
rect 4406 2048 4410 2052
rect 4686 2048 4690 2052
rect 4574 2038 4578 2042
rect 4442 2003 4446 2007
rect 4449 2003 4453 2007
rect 4382 1948 4386 1952
rect 4422 1948 4426 1952
rect 4510 1948 4514 1952
rect 4102 1938 4106 1942
rect 4350 1938 4354 1942
rect 4414 1938 4418 1942
rect 4438 1938 4442 1942
rect 4094 1918 4098 1922
rect 4142 1918 4146 1922
rect 4190 1918 4194 1922
rect 4238 1908 4242 1912
rect 4390 1928 4394 1932
rect 4254 1898 4258 1902
rect 4342 1898 4346 1902
rect 4190 1888 4194 1892
rect 4110 1878 4114 1882
rect 4158 1878 4162 1882
rect 4182 1878 4186 1882
rect 4270 1888 4274 1892
rect 4302 1888 4306 1892
rect 4366 1888 4370 1892
rect 4198 1878 4202 1882
rect 4238 1878 4242 1882
rect 4190 1868 4194 1872
rect 4046 1848 4050 1852
rect 4054 1838 4058 1842
rect 4014 1828 4018 1832
rect 3982 1788 3986 1792
rect 3862 1728 3866 1732
rect 3798 1708 3802 1712
rect 3830 1698 3834 1702
rect 3774 1688 3778 1692
rect 3806 1688 3810 1692
rect 3678 1668 3682 1672
rect 3710 1668 3714 1672
rect 3742 1668 3746 1672
rect 3702 1638 3706 1642
rect 3678 1608 3682 1612
rect 3670 1598 3674 1602
rect 3670 1558 3674 1562
rect 3686 1558 3690 1562
rect 3646 1548 3650 1552
rect 3718 1548 3722 1552
rect 3630 1538 3634 1542
rect 3622 1518 3626 1522
rect 3550 1488 3554 1492
rect 3550 1478 3554 1482
rect 3518 1468 3522 1472
rect 3574 1468 3578 1472
rect 3582 1468 3586 1472
rect 3558 1418 3562 1422
rect 3510 1398 3514 1402
rect 3526 1388 3530 1392
rect 3566 1388 3570 1392
rect 3438 1348 3442 1352
rect 3406 1328 3410 1332
rect 3390 1278 3394 1282
rect 3462 1278 3466 1282
rect 3534 1348 3538 1352
rect 3494 1338 3498 1342
rect 3358 1268 3362 1272
rect 3390 1268 3394 1272
rect 3478 1268 3482 1272
rect 3342 1258 3346 1262
rect 3334 1208 3338 1212
rect 3206 1058 3210 1062
rect 3198 1048 3202 1052
rect 3166 1038 3170 1042
rect 3126 978 3130 982
rect 3198 1038 3202 1042
rect 3158 968 3162 972
rect 3182 968 3186 972
rect 3150 958 3154 962
rect 3086 948 3090 952
rect 3134 948 3138 952
rect 3182 948 3186 952
rect 3222 1028 3226 1032
rect 3262 1048 3266 1052
rect 3230 1018 3234 1022
rect 3358 1108 3362 1112
rect 3406 1258 3410 1262
rect 3382 1218 3386 1222
rect 3334 1078 3338 1082
rect 3326 1028 3330 1032
rect 3318 1018 3322 1022
rect 3214 948 3218 952
rect 3230 948 3234 952
rect 3238 948 3242 952
rect 3294 948 3298 952
rect 3046 938 3050 942
rect 3054 938 3058 942
rect 3150 938 3154 942
rect 3198 938 3202 942
rect 3270 938 3274 942
rect 3094 928 3098 932
rect 3118 928 3122 932
rect 3142 928 3146 932
rect 3134 918 3138 922
rect 3022 908 3026 912
rect 3030 888 3034 892
rect 3054 888 3058 892
rect 3078 888 3082 892
rect 2974 878 2978 882
rect 3030 878 3034 882
rect 3038 878 3042 882
rect 3118 878 3122 882
rect 3126 878 3130 882
rect 2942 868 2946 872
rect 2974 868 2978 872
rect 3158 878 3162 882
rect 3078 868 3082 872
rect 3110 868 3114 872
rect 2958 858 2962 862
rect 2990 848 2994 852
rect 3038 848 3042 852
rect 3054 848 3058 852
rect 3054 818 3058 822
rect 2934 798 2938 802
rect 2942 798 2946 802
rect 2886 788 2890 792
rect 2910 788 2914 792
rect 2774 778 2778 782
rect 2238 758 2242 762
rect 2246 758 2250 762
rect 2270 758 2274 762
rect 2318 748 2322 752
rect 2230 738 2234 742
rect 2278 738 2282 742
rect 2310 738 2314 742
rect 2198 638 2202 642
rect 2182 498 2186 502
rect 2438 758 2442 762
rect 2470 758 2474 762
rect 2534 758 2538 762
rect 2606 758 2610 762
rect 2350 748 2354 752
rect 2430 748 2434 752
rect 2462 748 2466 752
rect 2374 738 2378 742
rect 2446 738 2450 742
rect 2238 728 2242 732
rect 2254 728 2258 732
rect 2438 728 2442 732
rect 2454 728 2458 732
rect 2462 728 2466 732
rect 2502 728 2506 732
rect 2318 718 2322 722
rect 2374 718 2378 722
rect 2302 698 2306 702
rect 2286 688 2290 692
rect 2278 668 2282 672
rect 2294 648 2298 652
rect 2286 628 2290 632
rect 2262 548 2266 552
rect 2294 548 2298 552
rect 2270 498 2274 502
rect 2182 488 2186 492
rect 2222 488 2226 492
rect 2222 478 2226 482
rect 1998 458 2002 462
rect 2014 458 2018 462
rect 2206 458 2210 462
rect 2278 458 2282 462
rect 1950 448 1954 452
rect 1998 448 2002 452
rect 2038 448 2042 452
rect 1958 438 1962 442
rect 1918 428 1922 432
rect 1974 428 1978 432
rect 1958 418 1962 422
rect 1918 398 1922 402
rect 1910 388 1914 392
rect 1926 388 1930 392
rect 1934 368 1938 372
rect 1950 368 1954 372
rect 2086 378 2090 382
rect 2094 378 2098 382
rect 2030 348 2034 352
rect 2062 348 2066 352
rect 1966 328 1970 332
rect 1766 268 1770 272
rect 1782 268 1786 272
rect 1830 268 1834 272
rect 1870 268 1874 272
rect 1814 258 1818 262
rect 1854 258 1858 262
rect 1654 248 1658 252
rect 1726 248 1730 252
rect 1814 248 1818 252
rect 1846 248 1850 252
rect 1638 238 1642 242
rect 1654 198 1658 202
rect 1662 198 1666 202
rect 1710 198 1714 202
rect 1686 188 1690 192
rect 1782 188 1786 192
rect 1838 188 1842 192
rect 1846 188 1850 192
rect 1878 168 1882 172
rect 1622 158 1626 162
rect 1518 138 1522 142
rect 1534 138 1538 142
rect 1550 138 1554 142
rect 1582 138 1586 142
rect 1510 128 1514 132
rect 1486 98 1490 102
rect 1334 88 1338 92
rect 1358 88 1362 92
rect 1406 88 1410 92
rect 1502 88 1506 92
rect 1302 78 1306 82
rect 1310 78 1314 82
rect 1478 78 1482 82
rect 1526 128 1530 132
rect 1558 128 1562 132
rect 1582 128 1586 132
rect 1598 128 1602 132
rect 1606 118 1610 122
rect 1654 158 1658 162
rect 1686 158 1690 162
rect 1718 158 1722 162
rect 1758 158 1762 162
rect 1766 158 1770 162
rect 1694 138 1698 142
rect 1726 138 1730 142
rect 1742 138 1746 142
rect 1702 128 1706 132
rect 1742 128 1746 132
rect 1646 118 1650 122
rect 1702 118 1706 122
rect 1726 118 1730 122
rect 1630 108 1634 112
rect 1734 108 1738 112
rect 1790 138 1794 142
rect 1806 138 1810 142
rect 1822 138 1826 142
rect 1774 108 1778 112
rect 1814 108 1818 112
rect 1782 98 1786 102
rect 1630 88 1634 92
rect 1678 88 1682 92
rect 1766 88 1770 92
rect 1782 88 1786 92
rect 1806 88 1810 92
rect 1646 78 1650 82
rect 1670 78 1674 82
rect 1726 78 1730 82
rect 1758 78 1762 82
rect 1766 78 1770 82
rect 1214 68 1218 72
rect 1438 68 1442 72
rect 1534 68 1538 72
rect 1590 68 1594 72
rect 1102 58 1106 62
rect 1278 58 1282 62
rect 1382 58 1386 62
rect 1446 58 1450 62
rect 1486 58 1490 62
rect 270 48 274 52
rect 278 48 282 52
rect 478 48 482 52
rect 686 48 690 52
rect 718 48 722 52
rect 734 48 738 52
rect 958 48 962 52
rect 982 48 986 52
rect 1078 48 1082 52
rect 1150 48 1154 52
rect 1206 48 1210 52
rect 1238 48 1242 52
rect 1278 48 1282 52
rect 1310 48 1314 52
rect 1574 58 1578 62
rect 1622 58 1626 62
rect 1630 58 1634 62
rect 1686 68 1690 72
rect 1718 68 1722 72
rect 1750 68 1754 72
rect 1766 68 1770 72
rect 1790 68 1794 72
rect 1814 78 1818 82
rect 1854 128 1858 132
rect 1830 118 1834 122
rect 1838 118 1842 122
rect 1678 58 1682 62
rect 1686 58 1690 62
rect 1734 58 1738 62
rect 1846 108 1850 112
rect 1878 138 1882 142
rect 1862 118 1866 122
rect 1874 103 1878 107
rect 1881 103 1885 107
rect 1614 48 1618 52
rect 1654 48 1658 52
rect 1670 48 1674 52
rect 1782 48 1786 52
rect 702 38 706 42
rect 1134 38 1138 42
rect 1550 38 1554 42
rect 1582 38 1586 42
rect 1614 38 1618 42
rect 1230 18 1234 22
rect 486 8 490 12
rect 526 8 530 12
rect 558 8 562 12
rect 798 8 802 12
rect 1078 8 1082 12
rect 1110 8 1114 12
rect 1174 8 1178 12
rect 346 3 350 7
rect 353 3 357 7
rect 1254 8 1258 12
rect 1278 8 1282 12
rect 1294 8 1298 12
rect 1358 8 1362 12
rect 1390 8 1394 12
rect 1462 8 1466 12
rect 1478 8 1482 12
rect 1638 8 1642 12
rect 1678 8 1682 12
rect 1734 8 1738 12
rect 1798 8 1802 12
rect 1370 3 1374 7
rect 1377 3 1381 7
rect 2054 308 2058 312
rect 1982 278 1986 282
rect 2014 298 2018 302
rect 2086 308 2090 312
rect 2078 298 2082 302
rect 2030 288 2034 292
rect 2102 368 2106 372
rect 2126 368 2130 372
rect 2174 368 2178 372
rect 2246 368 2250 372
rect 2254 368 2258 372
rect 2182 348 2186 352
rect 2214 348 2218 352
rect 2142 338 2146 342
rect 2190 338 2194 342
rect 2134 318 2138 322
rect 2118 308 2122 312
rect 2110 298 2114 302
rect 2238 348 2242 352
rect 2222 338 2226 342
rect 2254 338 2258 342
rect 2230 328 2234 332
rect 2214 298 2218 302
rect 2222 288 2226 292
rect 2206 278 2210 282
rect 2230 278 2234 282
rect 1974 268 1978 272
rect 2150 268 2154 272
rect 2182 268 2186 272
rect 1958 258 1962 262
rect 1990 258 1994 262
rect 2038 258 2042 262
rect 1926 238 1930 242
rect 1918 218 1922 222
rect 1902 148 1906 152
rect 2086 208 2090 212
rect 1942 188 1946 192
rect 1982 188 1986 192
rect 2086 188 2090 192
rect 2110 188 2114 192
rect 1918 138 1922 142
rect 1910 118 1914 122
rect 2038 138 2042 142
rect 2510 718 2514 722
rect 2422 708 2426 712
rect 2462 698 2466 702
rect 2502 698 2506 702
rect 2510 698 2514 702
rect 2350 688 2354 692
rect 2438 688 2442 692
rect 2486 688 2490 692
rect 2318 678 2322 682
rect 2342 668 2346 672
rect 2430 668 2434 672
rect 2486 668 2490 672
rect 2326 658 2330 662
rect 2350 658 2354 662
rect 2366 658 2370 662
rect 2510 668 2514 672
rect 2438 658 2442 662
rect 2462 658 2466 662
rect 2494 658 2498 662
rect 2502 658 2506 662
rect 2518 658 2522 662
rect 2358 648 2362 652
rect 2374 648 2378 652
rect 2390 648 2394 652
rect 2438 648 2442 652
rect 2318 638 2322 642
rect 2374 638 2378 642
rect 2518 638 2522 642
rect 2310 628 2314 632
rect 2390 628 2394 632
rect 2318 618 2322 622
rect 2310 588 2314 592
rect 2462 608 2466 612
rect 2394 603 2398 607
rect 2401 603 2405 607
rect 2582 718 2586 722
rect 2550 708 2554 712
rect 2590 698 2594 702
rect 2646 738 2650 742
rect 2662 738 2666 742
rect 2630 718 2634 722
rect 2694 748 2698 752
rect 2718 748 2722 752
rect 2838 748 2842 752
rect 2902 748 2906 752
rect 3030 758 3034 762
rect 3158 858 3162 862
rect 3134 838 3138 842
rect 3150 838 3154 842
rect 3102 828 3106 832
rect 3094 818 3098 822
rect 3118 798 3122 802
rect 3062 758 3066 762
rect 3110 748 3114 752
rect 3134 748 3138 752
rect 2726 728 2730 732
rect 2782 728 2786 732
rect 2766 718 2770 722
rect 2758 708 2762 712
rect 2614 698 2618 702
rect 2630 698 2634 702
rect 2638 698 2642 702
rect 2718 698 2722 702
rect 2726 698 2730 702
rect 2606 678 2610 682
rect 2934 728 2938 732
rect 2814 718 2818 722
rect 2830 718 2834 722
rect 2854 708 2858 712
rect 2822 698 2826 702
rect 2662 688 2666 692
rect 2678 688 2682 692
rect 2718 688 2722 692
rect 2782 688 2786 692
rect 2654 678 2658 682
rect 2542 658 2546 662
rect 2542 648 2546 652
rect 2574 648 2578 652
rect 2558 638 2562 642
rect 2566 628 2570 632
rect 2654 658 2658 662
rect 2606 638 2610 642
rect 2582 608 2586 612
rect 2334 588 2338 592
rect 2374 588 2378 592
rect 2430 578 2434 582
rect 2654 628 2658 632
rect 2630 608 2634 612
rect 2534 568 2538 572
rect 2654 598 2658 602
rect 2358 558 2362 562
rect 2518 558 2522 562
rect 2574 558 2578 562
rect 2614 558 2618 562
rect 2622 558 2626 562
rect 2414 548 2418 552
rect 2422 548 2426 552
rect 2454 548 2458 552
rect 2534 548 2538 552
rect 2542 548 2546 552
rect 2318 538 2322 542
rect 2350 538 2354 542
rect 2398 538 2402 542
rect 2446 538 2450 542
rect 2486 538 2490 542
rect 2414 528 2418 532
rect 2454 528 2458 532
rect 2526 538 2530 542
rect 2366 518 2370 522
rect 2510 518 2514 522
rect 2590 538 2594 542
rect 2630 548 2634 552
rect 2782 678 2786 682
rect 2798 678 2802 682
rect 2670 668 2674 672
rect 2686 668 2690 672
rect 2718 668 2722 672
rect 2734 668 2738 672
rect 2766 668 2770 672
rect 2906 703 2910 707
rect 2913 703 2917 707
rect 3206 888 3210 892
rect 3286 928 3290 932
rect 3254 918 3258 922
rect 3230 898 3234 902
rect 3262 898 3266 902
rect 3286 898 3290 902
rect 3222 868 3226 872
rect 3334 918 3338 922
rect 3350 1018 3354 1022
rect 3366 968 3370 972
rect 3418 1203 3422 1207
rect 3425 1203 3429 1207
rect 3398 1158 3402 1162
rect 3430 1148 3434 1152
rect 3470 1148 3474 1152
rect 3470 1138 3474 1142
rect 3446 1098 3450 1102
rect 3406 1078 3410 1082
rect 3382 948 3386 952
rect 3342 898 3346 902
rect 3358 888 3362 892
rect 3222 858 3226 862
rect 3254 858 3258 862
rect 3294 858 3298 862
rect 3278 838 3282 842
rect 3278 828 3282 832
rect 3214 788 3218 792
rect 3198 758 3202 762
rect 3166 748 3170 752
rect 3150 738 3154 742
rect 3158 738 3162 742
rect 2966 698 2970 702
rect 3126 728 3130 732
rect 3142 728 3146 732
rect 3086 718 3090 722
rect 3126 708 3130 712
rect 3150 698 3154 702
rect 3158 698 3162 702
rect 2838 688 2842 692
rect 3054 688 3058 692
rect 2862 678 2866 682
rect 3086 678 3090 682
rect 2886 668 2890 672
rect 3030 668 3034 672
rect 2678 658 2682 662
rect 2710 658 2714 662
rect 2726 658 2730 662
rect 2766 658 2770 662
rect 2790 658 2794 662
rect 2878 658 2882 662
rect 2910 658 2914 662
rect 2974 658 2978 662
rect 2734 648 2738 652
rect 2822 648 2826 652
rect 2830 648 2834 652
rect 2686 638 2690 642
rect 2758 638 2762 642
rect 2742 608 2746 612
rect 3022 658 3026 662
rect 2942 648 2946 652
rect 2998 648 3002 652
rect 3022 648 3026 652
rect 2870 638 2874 642
rect 2766 598 2770 602
rect 2814 598 2818 602
rect 2862 588 2866 592
rect 2694 558 2698 562
rect 2846 558 2850 562
rect 2726 548 2730 552
rect 2774 548 2778 552
rect 2726 538 2730 542
rect 2734 538 2738 542
rect 2790 538 2794 542
rect 2566 518 2570 522
rect 2606 518 2610 522
rect 2646 518 2650 522
rect 2670 518 2674 522
rect 2558 508 2562 512
rect 2574 508 2578 512
rect 2358 468 2362 472
rect 2462 468 2466 472
rect 2334 458 2338 462
rect 2414 458 2418 462
rect 2446 458 2450 462
rect 2542 458 2546 462
rect 2262 258 2266 262
rect 2278 258 2282 262
rect 2174 238 2178 242
rect 2246 208 2250 212
rect 2062 138 2066 142
rect 2118 138 2122 142
rect 2166 138 2170 142
rect 2190 138 2194 142
rect 2046 128 2050 132
rect 2134 128 2138 132
rect 2142 128 2146 132
rect 2182 128 2186 132
rect 2030 108 2034 112
rect 1958 98 1962 102
rect 2086 108 2090 112
rect 2118 108 2122 112
rect 1942 78 1946 82
rect 2070 78 2074 82
rect 2102 78 2106 82
rect 1918 68 1922 72
rect 1958 58 1962 62
rect 2014 59 2018 63
rect 2038 58 2042 62
rect 2158 68 2162 72
rect 2190 68 2194 72
rect 2270 198 2274 202
rect 2262 68 2266 72
rect 2078 48 2082 52
rect 2094 48 2098 52
rect 2094 38 2098 42
rect 2078 28 2082 32
rect 2062 18 2066 22
rect 2046 8 2050 12
rect 2214 28 2218 32
rect 2126 8 2130 12
rect 2150 8 2154 12
rect 2182 8 2186 12
rect 2198 8 2202 12
rect 2246 18 2250 22
rect 2246 8 2250 12
rect 2270 8 2274 12
rect 2558 448 2562 452
rect 2526 438 2530 442
rect 2394 403 2398 407
rect 2401 403 2405 407
rect 2414 398 2418 402
rect 2374 348 2378 352
rect 2398 348 2402 352
rect 2406 338 2410 342
rect 2310 308 2314 312
rect 2350 288 2354 292
rect 2350 278 2354 282
rect 2446 378 2450 382
rect 2486 368 2490 372
rect 2510 348 2514 352
rect 2422 338 2426 342
rect 2470 328 2474 332
rect 2470 318 2474 322
rect 2478 318 2482 322
rect 2518 318 2522 322
rect 2462 288 2466 292
rect 2542 428 2546 432
rect 2622 498 2626 502
rect 2606 388 2610 392
rect 2534 368 2538 372
rect 2606 368 2610 372
rect 2566 348 2570 352
rect 2558 338 2562 342
rect 2542 328 2546 332
rect 2726 508 2730 512
rect 2718 488 2722 492
rect 2662 468 2666 472
rect 2638 388 2642 392
rect 2630 378 2634 382
rect 2654 378 2658 382
rect 2694 468 2698 472
rect 2702 458 2706 462
rect 2678 378 2682 382
rect 2670 368 2674 372
rect 2798 518 2802 522
rect 2734 488 2738 492
rect 2750 488 2754 492
rect 2782 488 2786 492
rect 2758 468 2762 472
rect 2766 468 2770 472
rect 2830 528 2834 532
rect 2838 488 2842 492
rect 2822 468 2826 472
rect 2718 438 2722 442
rect 2758 438 2762 442
rect 2694 428 2698 432
rect 2734 428 2738 432
rect 2774 458 2778 462
rect 2798 458 2802 462
rect 2806 448 2810 452
rect 2838 458 2842 462
rect 2830 448 2834 452
rect 2814 438 2818 442
rect 2806 428 2810 432
rect 2902 638 2906 642
rect 2950 638 2954 642
rect 2886 628 2890 632
rect 2982 628 2986 632
rect 3094 658 3098 662
rect 3038 608 3042 612
rect 3030 598 3034 602
rect 2998 578 3002 582
rect 3118 618 3122 622
rect 3046 588 3050 592
rect 2894 568 2898 572
rect 2958 558 2962 562
rect 2974 558 2978 562
rect 2990 558 2994 562
rect 2878 548 2882 552
rect 2950 548 2954 552
rect 2998 548 3002 552
rect 3014 548 3018 552
rect 2878 528 2882 532
rect 2926 528 2930 532
rect 2906 503 2910 507
rect 2913 503 2917 507
rect 2870 488 2874 492
rect 2878 488 2882 492
rect 2870 478 2874 482
rect 2910 478 2914 482
rect 3110 568 3114 572
rect 3062 558 3066 562
rect 3054 538 3058 542
rect 3022 528 3026 532
rect 3078 528 3082 532
rect 3102 548 3106 552
rect 3094 538 3098 542
rect 3094 518 3098 522
rect 3086 488 3090 492
rect 2878 468 2882 472
rect 2958 468 2962 472
rect 2974 468 2978 472
rect 3190 738 3194 742
rect 3230 738 3234 742
rect 3342 868 3346 872
rect 3318 858 3322 862
rect 3302 848 3306 852
rect 3310 848 3314 852
rect 3326 828 3330 832
rect 3326 818 3330 822
rect 3310 768 3314 772
rect 3342 838 3346 842
rect 3478 1118 3482 1122
rect 3470 1078 3474 1082
rect 3430 1068 3434 1072
rect 3542 1338 3546 1342
rect 3606 1488 3610 1492
rect 3606 1468 3610 1472
rect 3630 1498 3634 1502
rect 3678 1528 3682 1532
rect 3670 1518 3674 1522
rect 3702 1538 3706 1542
rect 3686 1508 3690 1512
rect 3630 1478 3634 1482
rect 3622 1418 3626 1422
rect 3590 1358 3594 1362
rect 3590 1338 3594 1342
rect 3550 1328 3554 1332
rect 3598 1328 3602 1332
rect 3542 1298 3546 1302
rect 3550 1288 3554 1292
rect 3566 1288 3570 1292
rect 3542 1278 3546 1282
rect 3558 1278 3562 1282
rect 3558 1268 3562 1272
rect 3678 1468 3682 1472
rect 3654 1448 3658 1452
rect 3686 1448 3690 1452
rect 3654 1438 3658 1442
rect 3646 1418 3650 1422
rect 3718 1518 3722 1522
rect 3702 1428 3706 1432
rect 3654 1358 3658 1362
rect 3726 1468 3730 1472
rect 3854 1668 3858 1672
rect 3758 1558 3762 1562
rect 3782 1548 3786 1552
rect 3822 1538 3826 1542
rect 3750 1508 3754 1512
rect 3774 1488 3778 1492
rect 3782 1478 3786 1482
rect 3838 1628 3842 1632
rect 3886 1688 3890 1692
rect 3862 1508 3866 1512
rect 3838 1498 3842 1502
rect 3902 1628 3906 1632
rect 3930 1703 3934 1707
rect 3937 1703 3941 1707
rect 3966 1668 3970 1672
rect 3950 1648 3954 1652
rect 3966 1598 3970 1602
rect 3918 1548 3922 1552
rect 3902 1538 3906 1542
rect 3894 1468 3898 1472
rect 3930 1503 3934 1507
rect 3937 1503 3941 1507
rect 4006 1718 4010 1722
rect 4070 1818 4074 1822
rect 4062 1808 4066 1812
rect 4278 1878 4282 1882
rect 4398 1878 4402 1882
rect 4254 1868 4258 1872
rect 4294 1868 4298 1872
rect 4310 1868 4314 1872
rect 4358 1868 4362 1872
rect 4382 1868 4386 1872
rect 4182 1858 4186 1862
rect 4238 1858 4242 1862
rect 4262 1858 4266 1862
rect 4326 1858 4330 1862
rect 4342 1858 4346 1862
rect 4358 1858 4362 1862
rect 4182 1838 4186 1842
rect 4214 1838 4218 1842
rect 4230 1838 4234 1842
rect 4102 1788 4106 1792
rect 4214 1798 4218 1802
rect 4238 1798 4242 1802
rect 4278 1798 4282 1802
rect 4198 1788 4202 1792
rect 4214 1788 4218 1792
rect 4190 1758 4194 1762
rect 4086 1748 4090 1752
rect 4182 1748 4186 1752
rect 4198 1748 4202 1752
rect 4262 1768 4266 1772
rect 4254 1748 4258 1752
rect 4286 1748 4290 1752
rect 4334 1798 4338 1802
rect 4350 1778 4354 1782
rect 4382 1798 4386 1802
rect 4366 1768 4370 1772
rect 4358 1758 4362 1762
rect 4310 1748 4314 1752
rect 4342 1748 4346 1752
rect 4366 1748 4370 1752
rect 4486 1918 4490 1922
rect 4518 1918 4522 1922
rect 4534 1918 4538 1922
rect 4422 1898 4426 1902
rect 4470 1898 4474 1902
rect 4454 1858 4458 1862
rect 4574 1918 4578 1922
rect 4598 1898 4602 1902
rect 4486 1858 4490 1862
rect 4494 1858 4498 1862
rect 4558 1868 4562 1872
rect 4590 1868 4594 1872
rect 4582 1858 4586 1862
rect 4534 1848 4538 1852
rect 4574 1848 4578 1852
rect 4598 1848 4602 1852
rect 4494 1838 4498 1842
rect 4574 1838 4578 1842
rect 4606 1838 4610 1842
rect 4502 1828 4506 1832
rect 4414 1768 4418 1772
rect 4442 1803 4446 1807
rect 4449 1803 4453 1807
rect 4478 1778 4482 1782
rect 4486 1768 4490 1772
rect 4542 1768 4546 1772
rect 4438 1758 4442 1762
rect 4542 1758 4546 1762
rect 4230 1738 4234 1742
rect 4294 1738 4298 1742
rect 4382 1738 4386 1742
rect 4406 1738 4410 1742
rect 4446 1738 4450 1742
rect 4510 1738 4514 1742
rect 4582 1768 4586 1772
rect 4718 2058 4722 2062
rect 4766 2058 4770 2062
rect 4774 2048 4778 2052
rect 4822 2038 4826 2042
rect 4954 2103 4958 2107
rect 4961 2103 4965 2107
rect 4958 2088 4962 2092
rect 5014 2128 5018 2132
rect 4998 2108 5002 2112
rect 5062 2138 5066 2142
rect 5150 2258 5154 2262
rect 5214 2258 5218 2262
rect 5142 2198 5146 2202
rect 5150 2188 5154 2192
rect 5246 2248 5250 2252
rect 5206 2238 5210 2242
rect 5262 2228 5266 2232
rect 5222 2208 5226 2212
rect 5262 2208 5266 2212
rect 5118 2178 5122 2182
rect 5190 2178 5194 2182
rect 5214 2178 5218 2182
rect 5094 2168 5098 2172
rect 5102 2168 5106 2172
rect 5078 2138 5082 2142
rect 5030 2118 5034 2122
rect 5078 2118 5082 2122
rect 5062 2098 5066 2102
rect 5086 2098 5090 2102
rect 5198 2168 5202 2172
rect 5198 2148 5202 2152
rect 5214 2138 5218 2142
rect 5102 2128 5106 2132
rect 5158 2128 5162 2132
rect 5182 2128 5186 2132
rect 5110 2108 5114 2112
rect 5046 2078 5050 2082
rect 5094 2078 5098 2082
rect 5174 2078 5178 2082
rect 4982 2068 4986 2072
rect 4990 2068 4994 2072
rect 4998 2068 5002 2072
rect 5078 2068 5082 2072
rect 5094 2068 5098 2072
rect 4830 2028 4834 2032
rect 5022 2028 5026 2032
rect 5054 2018 5058 2022
rect 5254 2168 5258 2172
rect 5230 2148 5234 2152
rect 5246 2148 5250 2152
rect 5254 2148 5258 2152
rect 5246 2138 5250 2142
rect 5230 2128 5234 2132
rect 5246 2128 5250 2132
rect 5142 2028 5146 2032
rect 5078 2018 5082 2022
rect 5094 2018 5098 2022
rect 5118 2018 5122 2022
rect 4798 2008 4802 2012
rect 5014 2008 5018 2012
rect 5038 2008 5042 2012
rect 5070 2008 5074 2012
rect 4710 1978 4714 1982
rect 5006 1998 5010 2002
rect 4886 1988 4890 1992
rect 4942 1988 4946 1992
rect 4838 1968 4842 1972
rect 4806 1948 4810 1952
rect 5038 1958 5042 1962
rect 5054 1958 5058 1962
rect 4910 1948 4914 1952
rect 5022 1938 5026 1942
rect 4742 1928 4746 1932
rect 4774 1918 4778 1922
rect 4686 1908 4690 1912
rect 4654 1878 4658 1882
rect 4954 1903 4958 1907
rect 4961 1903 4965 1907
rect 5246 2058 5250 2062
rect 5230 2048 5234 2052
rect 5254 2048 5258 2052
rect 5198 2038 5202 2042
rect 5230 2038 5234 2042
rect 5198 2018 5202 2022
rect 5166 1998 5170 2002
rect 5166 1988 5170 1992
rect 5214 1958 5218 1962
rect 5094 1948 5098 1952
rect 5062 1928 5066 1932
rect 5110 1918 5114 1922
rect 4774 1888 4778 1892
rect 4806 1888 4810 1892
rect 4918 1888 4922 1892
rect 4974 1888 4978 1892
rect 5046 1888 5050 1892
rect 4894 1878 4898 1882
rect 5014 1878 5018 1882
rect 5022 1878 5026 1882
rect 5078 1878 5082 1882
rect 4662 1868 4666 1872
rect 4678 1868 4682 1872
rect 4830 1868 4834 1872
rect 4638 1858 4642 1862
rect 4694 1858 4698 1862
rect 4630 1848 4634 1852
rect 4678 1848 4682 1852
rect 4838 1858 4842 1862
rect 4886 1858 4890 1862
rect 4942 1858 4946 1862
rect 4710 1848 4714 1852
rect 4694 1838 4698 1842
rect 4638 1798 4642 1802
rect 4710 1798 4714 1802
rect 4718 1798 4722 1802
rect 4662 1778 4666 1782
rect 4694 1778 4698 1782
rect 4622 1768 4626 1772
rect 4630 1758 4634 1762
rect 4686 1758 4690 1762
rect 4598 1748 4602 1752
rect 4574 1738 4578 1742
rect 4590 1738 4594 1742
rect 4614 1738 4618 1742
rect 4126 1728 4130 1732
rect 4302 1728 4306 1732
rect 4430 1728 4434 1732
rect 4486 1728 4490 1732
rect 4542 1728 4546 1732
rect 4558 1728 4562 1732
rect 4054 1718 4058 1722
rect 4118 1718 4122 1722
rect 4142 1708 4146 1712
rect 4086 1698 4090 1702
rect 4110 1678 4114 1682
rect 4166 1678 4170 1682
rect 4006 1668 4010 1672
rect 4046 1668 4050 1672
rect 3974 1538 3978 1542
rect 3990 1538 3994 1542
rect 4214 1658 4218 1662
rect 4254 1678 4258 1682
rect 4230 1668 4234 1672
rect 4286 1678 4290 1682
rect 4294 1668 4298 1672
rect 4270 1658 4274 1662
rect 4382 1718 4386 1722
rect 4462 1718 4466 1722
rect 4334 1698 4338 1702
rect 4310 1658 4314 1662
rect 4462 1708 4466 1712
rect 4470 1698 4474 1702
rect 4558 1688 4562 1692
rect 4350 1678 4354 1682
rect 4358 1678 4362 1682
rect 4422 1678 4426 1682
rect 4526 1678 4530 1682
rect 4350 1668 4354 1672
rect 4390 1668 4394 1672
rect 4414 1668 4418 1672
rect 4526 1668 4530 1672
rect 4534 1668 4538 1672
rect 4262 1648 4266 1652
rect 4286 1648 4290 1652
rect 4342 1648 4346 1652
rect 4158 1638 4162 1642
rect 4246 1638 4250 1642
rect 4366 1638 4370 1642
rect 4446 1638 4450 1642
rect 4022 1548 4026 1552
rect 4014 1538 4018 1542
rect 4006 1488 4010 1492
rect 4070 1478 4074 1482
rect 3766 1448 3770 1452
rect 3822 1448 3826 1452
rect 3782 1438 3786 1442
rect 3766 1428 3770 1432
rect 3806 1428 3810 1432
rect 3718 1358 3722 1362
rect 3758 1358 3762 1362
rect 3790 1398 3794 1402
rect 3846 1398 3850 1402
rect 3822 1358 3826 1362
rect 3886 1358 3890 1362
rect 3790 1338 3794 1342
rect 3710 1328 3714 1332
rect 3646 1308 3650 1312
rect 3662 1308 3666 1312
rect 3694 1308 3698 1312
rect 3590 1288 3594 1292
rect 3622 1288 3626 1292
rect 3654 1288 3658 1292
rect 3614 1268 3618 1272
rect 3638 1268 3642 1272
rect 3654 1268 3658 1272
rect 3502 1248 3506 1252
rect 3582 1248 3586 1252
rect 3606 1248 3610 1252
rect 3526 1228 3530 1232
rect 3502 1158 3506 1162
rect 3494 1128 3498 1132
rect 3622 1218 3626 1222
rect 3558 1158 3562 1162
rect 3590 1158 3594 1162
rect 3606 1158 3610 1162
rect 3542 1148 3546 1152
rect 3582 1148 3586 1152
rect 3622 1148 3626 1152
rect 3534 1138 3538 1142
rect 3614 1128 3618 1132
rect 3502 1108 3506 1112
rect 3526 1108 3530 1112
rect 3558 1078 3562 1082
rect 3418 1003 3422 1007
rect 3425 1003 3429 1007
rect 3574 1108 3578 1112
rect 3582 1098 3586 1102
rect 3638 1088 3642 1092
rect 3670 1298 3674 1302
rect 3686 1278 3690 1282
rect 3702 1278 3706 1282
rect 3678 1258 3682 1262
rect 3814 1338 3818 1342
rect 3822 1338 3826 1342
rect 3774 1328 3778 1332
rect 3806 1328 3810 1332
rect 3734 1288 3738 1292
rect 3798 1288 3802 1292
rect 3718 1278 3722 1282
rect 3782 1258 3786 1262
rect 3742 1158 3746 1162
rect 3774 1158 3778 1162
rect 3686 1147 3690 1151
rect 3726 1148 3730 1152
rect 3726 1118 3730 1122
rect 3710 1098 3714 1102
rect 3742 1088 3746 1092
rect 3614 1078 3618 1082
rect 3630 1078 3634 1082
rect 3638 1078 3642 1082
rect 3662 1078 3666 1082
rect 3678 1078 3682 1082
rect 3566 1068 3570 1072
rect 3598 1068 3602 1072
rect 3622 1068 3626 1072
rect 3494 1038 3498 1042
rect 3574 1018 3578 1022
rect 3478 968 3482 972
rect 3422 958 3426 962
rect 3470 938 3474 942
rect 3494 938 3498 942
rect 3462 928 3466 932
rect 3390 918 3394 922
rect 3382 878 3386 882
rect 3422 898 3426 902
rect 3398 878 3402 882
rect 3526 948 3530 952
rect 3502 928 3506 932
rect 3510 918 3514 922
rect 3518 908 3522 912
rect 3518 898 3522 902
rect 3478 888 3482 892
rect 3494 888 3498 892
rect 3510 888 3514 892
rect 3430 878 3434 882
rect 3454 878 3458 882
rect 3478 878 3482 882
rect 3430 868 3434 872
rect 3478 868 3482 872
rect 3462 858 3466 862
rect 3374 828 3378 832
rect 3418 803 3422 807
rect 3425 803 3429 807
rect 3350 788 3354 792
rect 3366 788 3370 792
rect 3454 788 3458 792
rect 3470 768 3474 772
rect 3502 768 3506 772
rect 3390 758 3394 762
rect 3430 758 3434 762
rect 3462 758 3466 762
rect 3334 748 3338 752
rect 3382 748 3386 752
rect 3278 738 3282 742
rect 3310 738 3314 742
rect 3262 718 3266 722
rect 3254 698 3258 702
rect 3174 688 3178 692
rect 3214 678 3218 682
rect 3302 688 3306 692
rect 3414 748 3418 752
rect 3446 748 3450 752
rect 3454 748 3458 752
rect 3374 738 3378 742
rect 3398 738 3402 742
rect 3398 728 3402 732
rect 3430 728 3434 732
rect 3350 718 3354 722
rect 3150 658 3154 662
rect 3230 658 3234 662
rect 3318 658 3322 662
rect 3142 588 3146 592
rect 3534 928 3538 932
rect 3566 908 3570 912
rect 3542 898 3546 902
rect 3646 1048 3650 1052
rect 3590 1028 3594 1032
rect 3726 1058 3730 1062
rect 3702 1048 3706 1052
rect 3758 1048 3762 1052
rect 3654 1038 3658 1042
rect 3694 1038 3698 1042
rect 3710 1038 3714 1042
rect 3614 968 3618 972
rect 3630 968 3634 972
rect 3646 968 3650 972
rect 3590 948 3594 952
rect 3614 948 3618 952
rect 3590 938 3594 942
rect 3622 938 3626 942
rect 3694 988 3698 992
rect 3670 958 3674 962
rect 3638 898 3642 902
rect 3614 878 3618 882
rect 3782 1128 3786 1132
rect 3798 1108 3802 1112
rect 3774 1018 3778 1022
rect 3726 988 3730 992
rect 3774 968 3778 972
rect 3718 948 3722 952
rect 3758 948 3762 952
rect 3726 928 3730 932
rect 3718 898 3722 902
rect 3830 1318 3834 1322
rect 3974 1468 3978 1472
rect 4190 1618 4194 1622
rect 4302 1618 4306 1622
rect 4150 1608 4154 1612
rect 4126 1588 4130 1592
rect 4142 1588 4146 1592
rect 4094 1578 4098 1582
rect 4246 1558 4250 1562
rect 4206 1547 4210 1551
rect 4246 1548 4250 1552
rect 4442 1603 4446 1607
rect 4449 1603 4453 1607
rect 4502 1658 4506 1662
rect 4518 1658 4522 1662
rect 4574 1678 4578 1682
rect 4598 1678 4602 1682
rect 4598 1668 4602 1672
rect 4582 1658 4586 1662
rect 4510 1648 4514 1652
rect 4502 1638 4506 1642
rect 4494 1568 4498 1572
rect 4422 1558 4426 1562
rect 4478 1558 4482 1562
rect 4358 1548 4362 1552
rect 4382 1548 4386 1552
rect 4406 1548 4410 1552
rect 4510 1548 4514 1552
rect 4534 1558 4538 1562
rect 4558 1558 4562 1562
rect 4542 1548 4546 1552
rect 4574 1548 4578 1552
rect 4414 1538 4418 1542
rect 4486 1538 4490 1542
rect 4518 1538 4522 1542
rect 4086 1508 4090 1512
rect 4102 1508 4106 1512
rect 4086 1478 4090 1482
rect 4174 1488 4178 1492
rect 4134 1478 4138 1482
rect 4086 1448 4090 1452
rect 4046 1418 4050 1422
rect 4014 1398 4018 1402
rect 4078 1358 4082 1362
rect 3966 1348 3970 1352
rect 3930 1303 3934 1307
rect 3937 1303 3941 1307
rect 4030 1348 4034 1352
rect 4086 1348 4090 1352
rect 3982 1338 3986 1342
rect 4014 1338 4018 1342
rect 3934 1288 3938 1292
rect 3958 1288 3962 1292
rect 3894 1278 3898 1282
rect 3894 1268 3898 1272
rect 4270 1518 4274 1522
rect 4286 1508 4290 1512
rect 4342 1518 4346 1522
rect 4318 1498 4322 1502
rect 4262 1488 4266 1492
rect 4446 1528 4450 1532
rect 4494 1528 4498 1532
rect 4486 1518 4490 1522
rect 4502 1518 4506 1522
rect 4350 1508 4354 1512
rect 4374 1508 4378 1512
rect 4414 1508 4418 1512
rect 4406 1498 4410 1502
rect 4374 1488 4378 1492
rect 4150 1468 4154 1472
rect 4118 1458 4122 1462
rect 4206 1458 4210 1462
rect 4150 1448 4154 1452
rect 4158 1448 4162 1452
rect 4142 1438 4146 1442
rect 4126 1388 4130 1392
rect 4102 1378 4106 1382
rect 4094 1338 4098 1342
rect 4094 1288 4098 1292
rect 4150 1408 4154 1412
rect 4150 1398 4154 1402
rect 4294 1458 4298 1462
rect 4262 1428 4266 1432
rect 4198 1408 4202 1412
rect 4174 1358 4178 1362
rect 4294 1428 4298 1432
rect 4270 1388 4274 1392
rect 4222 1368 4226 1372
rect 4318 1458 4322 1462
rect 4414 1488 4418 1492
rect 4470 1488 4474 1492
rect 4454 1468 4458 1472
rect 4494 1478 4498 1482
rect 4478 1468 4482 1472
rect 4510 1508 4514 1512
rect 4526 1498 4530 1502
rect 4510 1468 4514 1472
rect 4470 1458 4474 1462
rect 4438 1448 4442 1452
rect 4310 1418 4314 1422
rect 4334 1388 4338 1392
rect 4350 1388 4354 1392
rect 4318 1378 4322 1382
rect 4214 1358 4218 1362
rect 4262 1358 4266 1362
rect 4302 1358 4306 1362
rect 4198 1348 4202 1352
rect 4230 1348 4234 1352
rect 4286 1348 4290 1352
rect 4238 1338 4242 1342
rect 4262 1338 4266 1342
rect 4214 1328 4218 1332
rect 4262 1328 4266 1332
rect 4166 1308 4170 1312
rect 4158 1298 4162 1302
rect 4246 1308 4250 1312
rect 4246 1288 4250 1292
rect 4134 1268 4138 1272
rect 3950 1258 3954 1262
rect 3830 1148 3834 1152
rect 3998 1158 4002 1162
rect 3958 1148 3962 1152
rect 3990 1148 3994 1152
rect 3862 1138 3866 1142
rect 3974 1138 3978 1142
rect 4006 1138 4010 1142
rect 3846 1098 3850 1102
rect 3830 1088 3834 1092
rect 3822 1078 3826 1082
rect 3854 1008 3858 1012
rect 3822 968 3826 972
rect 3846 968 3850 972
rect 3854 968 3858 972
rect 3806 958 3810 962
rect 3814 958 3818 962
rect 3830 958 3834 962
rect 3862 948 3866 952
rect 3790 938 3794 942
rect 3910 1128 3914 1132
rect 3958 1128 3962 1132
rect 3886 1088 3890 1092
rect 3930 1103 3934 1107
rect 3937 1103 3941 1107
rect 3998 1128 4002 1132
rect 4062 1218 4066 1222
rect 4110 1218 4114 1222
rect 4054 1188 4058 1192
rect 4038 1158 4042 1162
rect 4094 1178 4098 1182
rect 3974 1088 3978 1092
rect 3990 1088 3994 1092
rect 4022 1088 4026 1092
rect 3966 1078 3970 1082
rect 3934 1068 3938 1072
rect 3886 1058 3890 1062
rect 3902 1038 3906 1042
rect 3958 1058 3962 1062
rect 3934 1018 3938 1022
rect 3910 1008 3914 1012
rect 4046 1128 4050 1132
rect 4102 1158 4106 1162
rect 4310 1338 4314 1342
rect 4302 1328 4306 1332
rect 4390 1438 4394 1442
rect 4442 1403 4446 1407
rect 4449 1403 4453 1407
rect 4486 1448 4490 1452
rect 4510 1448 4514 1452
rect 4470 1418 4474 1422
rect 4502 1388 4506 1392
rect 4462 1368 4466 1372
rect 4470 1368 4474 1372
rect 4486 1368 4490 1372
rect 4342 1358 4346 1362
rect 4366 1358 4370 1362
rect 4502 1358 4506 1362
rect 4510 1358 4514 1362
rect 4406 1348 4410 1352
rect 4622 1658 4626 1662
rect 4638 1658 4642 1662
rect 4606 1638 4610 1642
rect 4622 1638 4626 1642
rect 4598 1568 4602 1572
rect 4582 1538 4586 1542
rect 4702 1768 4706 1772
rect 4742 1788 4746 1792
rect 4742 1778 4746 1782
rect 4766 1768 4770 1772
rect 4750 1758 4754 1762
rect 4814 1758 4818 1762
rect 4830 1758 4834 1762
rect 4734 1748 4738 1752
rect 4750 1748 4754 1752
rect 4814 1748 4818 1752
rect 4822 1748 4826 1752
rect 4670 1738 4674 1742
rect 4726 1738 4730 1742
rect 4766 1738 4770 1742
rect 4662 1688 4666 1692
rect 4662 1668 4666 1672
rect 4702 1718 4706 1722
rect 4678 1678 4682 1682
rect 4686 1658 4690 1662
rect 4686 1648 4690 1652
rect 4694 1638 4698 1642
rect 4678 1628 4682 1632
rect 4654 1618 4658 1622
rect 4662 1588 4666 1592
rect 5070 1858 5074 1862
rect 5126 1858 5130 1862
rect 5134 1848 5138 1852
rect 4950 1818 4954 1822
rect 5046 1808 5050 1812
rect 4910 1798 4914 1802
rect 4878 1778 4882 1782
rect 4862 1768 4866 1772
rect 4894 1768 4898 1772
rect 4926 1768 4930 1772
rect 4942 1768 4946 1772
rect 4854 1758 4858 1762
rect 4894 1758 4898 1762
rect 4846 1738 4850 1742
rect 4958 1758 4962 1762
rect 5014 1758 5018 1762
rect 4878 1748 4882 1752
rect 4902 1748 4906 1752
rect 4926 1748 4930 1752
rect 4942 1748 4946 1752
rect 4798 1688 4802 1692
rect 4822 1688 4826 1692
rect 4886 1738 4890 1742
rect 4766 1678 4770 1682
rect 4806 1678 4810 1682
rect 4830 1678 4834 1682
rect 4838 1678 4842 1682
rect 4870 1678 4874 1682
rect 4718 1668 4722 1672
rect 4726 1658 4730 1662
rect 4782 1668 4786 1672
rect 5070 1758 5074 1762
rect 4966 1748 4970 1752
rect 5014 1738 5018 1742
rect 4950 1728 4954 1732
rect 5006 1708 5010 1712
rect 5038 1708 5042 1712
rect 4954 1703 4958 1707
rect 4961 1703 4965 1707
rect 4950 1688 4954 1692
rect 5166 1888 5170 1892
rect 5214 1938 5218 1942
rect 5198 1878 5202 1882
rect 5278 2278 5282 2282
rect 5278 2258 5282 2262
rect 5278 2208 5282 2212
rect 5278 2178 5282 2182
rect 5270 2158 5274 2162
rect 5286 2148 5290 2152
rect 5302 2328 5306 2332
rect 5302 2278 5306 2282
rect 5302 2158 5306 2162
rect 5302 2138 5306 2142
rect 5294 2128 5298 2132
rect 5310 2128 5314 2132
rect 5278 2088 5282 2092
rect 5262 1968 5266 1972
rect 5238 1958 5242 1962
rect 5262 1948 5266 1952
rect 5238 1888 5242 1892
rect 5214 1868 5218 1872
rect 5246 1868 5250 1872
rect 5198 1858 5202 1862
rect 5206 1858 5210 1862
rect 5230 1858 5234 1862
rect 5182 1848 5186 1852
rect 5222 1838 5226 1842
rect 5158 1828 5162 1832
rect 5142 1808 5146 1812
rect 5214 1768 5218 1772
rect 5214 1758 5218 1762
rect 5238 1758 5242 1762
rect 5110 1748 5114 1752
rect 5094 1738 5098 1742
rect 5238 1738 5242 1742
rect 5158 1728 5162 1732
rect 5102 1718 5106 1722
rect 5046 1688 5050 1692
rect 5078 1688 5082 1692
rect 5006 1678 5010 1682
rect 4758 1658 4762 1662
rect 4798 1658 4802 1662
rect 4750 1648 4754 1652
rect 4774 1648 4778 1652
rect 4646 1568 4650 1572
rect 4686 1548 4690 1552
rect 4614 1528 4618 1532
rect 4630 1528 4634 1532
rect 4574 1508 4578 1512
rect 4598 1508 4602 1512
rect 4542 1488 4546 1492
rect 4566 1488 4570 1492
rect 4590 1478 4594 1482
rect 4606 1488 4610 1492
rect 4542 1468 4546 1472
rect 4550 1468 4554 1472
rect 4582 1468 4586 1472
rect 4694 1518 4698 1522
rect 4742 1568 4746 1572
rect 4790 1618 4794 1622
rect 4886 1668 4890 1672
rect 4918 1668 4922 1672
rect 4942 1668 4946 1672
rect 4846 1648 4850 1652
rect 4886 1638 4890 1642
rect 4806 1598 4810 1602
rect 4822 1598 4826 1602
rect 4798 1588 4802 1592
rect 4814 1588 4818 1592
rect 4782 1568 4786 1572
rect 4806 1568 4810 1572
rect 4710 1558 4714 1562
rect 4734 1558 4738 1562
rect 4758 1558 4762 1562
rect 4766 1558 4770 1562
rect 4798 1558 4802 1562
rect 4766 1548 4770 1552
rect 4798 1548 4802 1552
rect 4814 1548 4818 1552
rect 4894 1558 4898 1562
rect 4822 1538 4826 1542
rect 4734 1508 4738 1512
rect 4710 1498 4714 1502
rect 4862 1518 4866 1522
rect 4702 1488 4706 1492
rect 4766 1488 4770 1492
rect 4806 1478 4810 1482
rect 4846 1478 4850 1482
rect 4886 1478 4890 1482
rect 4782 1468 4786 1472
rect 4814 1468 4818 1472
rect 4846 1468 4850 1472
rect 4662 1458 4666 1462
rect 4678 1458 4682 1462
rect 4694 1458 4698 1462
rect 4750 1458 4754 1462
rect 4774 1458 4778 1462
rect 4790 1448 4794 1452
rect 4814 1448 4818 1452
rect 4558 1438 4562 1442
rect 4638 1438 4642 1442
rect 4894 1458 4898 1462
rect 4886 1448 4890 1452
rect 4910 1588 4914 1592
rect 4934 1578 4938 1582
rect 4918 1558 4922 1562
rect 4918 1538 4922 1542
rect 4926 1528 4930 1532
rect 4918 1478 4922 1482
rect 4918 1468 4922 1472
rect 5014 1568 5018 1572
rect 5038 1568 5042 1572
rect 5062 1568 5066 1572
rect 5110 1688 5114 1692
rect 5102 1658 5106 1662
rect 4974 1558 4978 1562
rect 5030 1558 5034 1562
rect 5054 1548 5058 1552
rect 5014 1538 5018 1542
rect 5054 1538 5058 1542
rect 4942 1518 4946 1522
rect 4954 1503 4958 1507
rect 4961 1503 4965 1507
rect 4942 1468 4946 1472
rect 4974 1468 4978 1472
rect 4798 1428 4802 1432
rect 4822 1428 4826 1432
rect 4830 1428 4834 1432
rect 4654 1368 4658 1372
rect 4678 1368 4682 1372
rect 4766 1368 4770 1372
rect 4598 1358 4602 1362
rect 4550 1348 4554 1352
rect 4566 1338 4570 1342
rect 4622 1348 4626 1352
rect 4702 1358 4706 1362
rect 4686 1348 4690 1352
rect 4846 1428 4850 1432
rect 4854 1388 4858 1392
rect 4846 1358 4850 1362
rect 4350 1328 4354 1332
rect 4486 1328 4490 1332
rect 4518 1328 4522 1332
rect 4606 1328 4610 1332
rect 4334 1298 4338 1302
rect 4382 1298 4386 1302
rect 4326 1288 4330 1292
rect 4310 1268 4314 1272
rect 4246 1258 4250 1262
rect 4270 1258 4274 1262
rect 4198 1178 4202 1182
rect 4150 1168 4154 1172
rect 4166 1168 4170 1172
rect 4230 1168 4234 1172
rect 4118 1148 4122 1152
rect 4206 1148 4210 1152
rect 4238 1148 4242 1152
rect 4190 1138 4194 1142
rect 4222 1138 4226 1142
rect 4126 1088 4130 1092
rect 4070 1078 4074 1082
rect 4030 1068 4034 1072
rect 4078 1058 4082 1062
rect 4110 1058 4114 1062
rect 4006 1038 4010 1042
rect 4022 1038 4026 1042
rect 3990 1008 3994 1012
rect 4062 1008 4066 1012
rect 3990 988 3994 992
rect 3982 968 3986 972
rect 4022 968 4026 972
rect 3878 948 3882 952
rect 3894 948 3898 952
rect 3958 948 3962 952
rect 3886 938 3890 942
rect 3950 938 3954 942
rect 3870 888 3874 892
rect 3694 878 3698 882
rect 3734 878 3738 882
rect 3838 878 3842 882
rect 3942 918 3946 922
rect 3930 903 3934 907
rect 3937 903 3941 907
rect 3718 868 3722 872
rect 3662 858 3666 862
rect 3630 848 3634 852
rect 3574 818 3578 822
rect 3558 758 3562 762
rect 3526 748 3530 752
rect 3614 808 3618 812
rect 3686 848 3690 852
rect 3694 848 3698 852
rect 3694 828 3698 832
rect 3638 798 3642 802
rect 3726 798 3730 802
rect 3766 868 3770 872
rect 3854 868 3858 872
rect 3870 868 3874 872
rect 3886 868 3890 872
rect 3790 858 3794 862
rect 3862 858 3866 862
rect 3918 858 3922 862
rect 4038 948 4042 952
rect 3974 938 3978 942
rect 3998 938 4002 942
rect 4094 938 4098 942
rect 4030 928 4034 932
rect 4046 928 4050 932
rect 3966 898 3970 902
rect 4078 898 4082 902
rect 3966 888 3970 892
rect 4038 888 4042 892
rect 3990 878 3994 882
rect 4054 878 4058 882
rect 4022 868 4026 872
rect 4038 868 4042 872
rect 4054 868 4058 872
rect 4070 868 4074 872
rect 3958 848 3962 852
rect 3838 838 3842 842
rect 3854 838 3858 842
rect 3934 838 3938 842
rect 3718 788 3722 792
rect 3734 788 3738 792
rect 4118 978 4122 982
rect 4182 1128 4186 1132
rect 4206 1128 4210 1132
rect 4230 1128 4234 1132
rect 4214 1098 4218 1102
rect 4206 1088 4210 1092
rect 4238 1088 4242 1092
rect 4150 1048 4154 1052
rect 4182 1048 4186 1052
rect 4142 988 4146 992
rect 4134 968 4138 972
rect 4150 958 4154 962
rect 4166 948 4170 952
rect 4118 938 4122 942
rect 4134 938 4138 942
rect 4182 938 4186 942
rect 4238 1058 4242 1062
rect 4222 1048 4226 1052
rect 4262 1148 4266 1152
rect 4262 1138 4266 1142
rect 4350 1288 4354 1292
rect 4710 1318 4714 1322
rect 4694 1308 4698 1312
rect 4654 1288 4658 1292
rect 4494 1278 4498 1282
rect 4646 1278 4650 1282
rect 4790 1328 4794 1332
rect 4830 1338 4834 1342
rect 4846 1338 4850 1342
rect 4870 1368 4874 1372
rect 4966 1428 4970 1432
rect 4910 1408 4914 1412
rect 4902 1358 4906 1362
rect 4870 1338 4874 1342
rect 4846 1328 4850 1332
rect 4862 1328 4866 1332
rect 4798 1318 4802 1322
rect 4742 1308 4746 1312
rect 4886 1328 4890 1332
rect 4774 1278 4778 1282
rect 4790 1278 4794 1282
rect 4830 1278 4834 1282
rect 4342 1268 4346 1272
rect 4358 1268 4362 1272
rect 4638 1268 4642 1272
rect 4662 1268 4666 1272
rect 4774 1268 4778 1272
rect 4318 1258 4322 1262
rect 4294 1158 4298 1162
rect 4318 1178 4322 1182
rect 4302 1148 4306 1152
rect 4310 1138 4314 1142
rect 4366 1258 4370 1262
rect 4518 1258 4522 1262
rect 4438 1248 4442 1252
rect 4442 1203 4446 1207
rect 4449 1203 4453 1207
rect 4502 1188 4506 1192
rect 4430 1178 4434 1182
rect 4446 1178 4450 1182
rect 4342 1158 4346 1162
rect 4334 1148 4338 1152
rect 4374 1148 4378 1152
rect 4430 1148 4434 1152
rect 4382 1138 4386 1142
rect 4438 1128 4442 1132
rect 4350 1118 4354 1122
rect 4326 1088 4330 1092
rect 4478 1088 4482 1092
rect 4502 1088 4506 1092
rect 4350 1078 4354 1082
rect 4358 1078 4362 1082
rect 4558 1228 4562 1232
rect 4718 1258 4722 1262
rect 4582 1248 4586 1252
rect 4638 1248 4642 1252
rect 4750 1248 4754 1252
rect 4614 1218 4618 1222
rect 4574 1188 4578 1192
rect 4566 1128 4570 1132
rect 4558 1118 4562 1122
rect 4590 1118 4594 1122
rect 4622 1108 4626 1112
rect 4678 1188 4682 1192
rect 4678 1168 4682 1172
rect 4742 1158 4746 1162
rect 4686 1088 4690 1092
rect 4974 1348 4978 1352
rect 4926 1328 4930 1332
rect 4950 1318 4954 1322
rect 4954 1303 4958 1307
rect 4961 1303 4965 1307
rect 4990 1528 4994 1532
rect 5006 1528 5010 1532
rect 5142 1688 5146 1692
rect 5150 1678 5154 1682
rect 5134 1588 5138 1592
rect 5126 1578 5130 1582
rect 5166 1718 5170 1722
rect 5238 1708 5242 1712
rect 5190 1698 5194 1702
rect 5174 1688 5178 1692
rect 5198 1688 5202 1692
rect 5214 1688 5218 1692
rect 5190 1678 5194 1682
rect 5174 1668 5178 1672
rect 5230 1678 5234 1682
rect 5302 2088 5306 2092
rect 5294 1868 5298 1872
rect 5262 1858 5266 1862
rect 5262 1848 5266 1852
rect 5262 1778 5266 1782
rect 5270 1758 5274 1762
rect 5294 1758 5298 1762
rect 5286 1728 5290 1732
rect 5270 1718 5274 1722
rect 5278 1718 5282 1722
rect 5262 1708 5266 1712
rect 5294 1698 5298 1702
rect 5262 1688 5266 1692
rect 5182 1658 5186 1662
rect 5198 1658 5202 1662
rect 5222 1658 5226 1662
rect 5214 1648 5218 1652
rect 5214 1598 5218 1602
rect 5270 1658 5274 1662
rect 5174 1558 5178 1562
rect 5214 1558 5218 1562
rect 5230 1558 5234 1562
rect 5086 1548 5090 1552
rect 5158 1548 5162 1552
rect 5078 1538 5082 1542
rect 5070 1518 5074 1522
rect 5014 1508 5018 1512
rect 4990 1478 4994 1482
rect 5094 1528 5098 1532
rect 5102 1518 5106 1522
rect 5174 1518 5178 1522
rect 5150 1508 5154 1512
rect 5206 1518 5210 1522
rect 5270 1548 5274 1552
rect 5110 1488 5114 1492
rect 5062 1478 5066 1482
rect 5134 1478 5138 1482
rect 5150 1478 5154 1482
rect 5190 1478 5194 1482
rect 4998 1458 5002 1462
rect 5006 1428 5010 1432
rect 4998 1418 5002 1422
rect 5030 1468 5034 1472
rect 5046 1468 5050 1472
rect 5054 1468 5058 1472
rect 5102 1468 5106 1472
rect 5110 1458 5114 1462
rect 5102 1438 5106 1442
rect 5126 1438 5130 1442
rect 5110 1428 5114 1432
rect 5062 1418 5066 1422
rect 5038 1348 5042 1352
rect 5006 1338 5010 1342
rect 5014 1338 5018 1342
rect 5054 1328 5058 1332
rect 5070 1308 5074 1312
rect 5062 1298 5066 1302
rect 5014 1278 5018 1282
rect 5062 1278 5066 1282
rect 4934 1268 4938 1272
rect 5006 1268 5010 1272
rect 4806 1258 4810 1262
rect 4782 1248 4786 1252
rect 4798 1248 4802 1252
rect 4830 1248 4834 1252
rect 4838 1248 4842 1252
rect 4886 1248 4890 1252
rect 4846 1238 4850 1242
rect 4902 1238 4906 1242
rect 5094 1338 5098 1342
rect 5110 1338 5114 1342
rect 5158 1468 5162 1472
rect 5174 1468 5178 1472
rect 5142 1458 5146 1462
rect 5150 1458 5154 1462
rect 5174 1458 5178 1462
rect 5182 1438 5186 1442
rect 5174 1418 5178 1422
rect 5150 1348 5154 1352
rect 5182 1348 5186 1352
rect 5142 1338 5146 1342
rect 5166 1338 5170 1342
rect 5134 1328 5138 1332
rect 5126 1308 5130 1312
rect 5134 1298 5138 1302
rect 5150 1328 5154 1332
rect 5238 1538 5242 1542
rect 5246 1528 5250 1532
rect 5270 1518 5274 1522
rect 5278 1518 5282 1522
rect 5302 1498 5306 1502
rect 5278 1488 5282 1492
rect 5294 1488 5298 1492
rect 5246 1478 5250 1482
rect 5278 1478 5282 1482
rect 5230 1468 5234 1472
rect 5246 1468 5250 1472
rect 5270 1468 5274 1472
rect 5206 1458 5210 1462
rect 5230 1448 5234 1452
rect 5214 1418 5218 1422
rect 5214 1378 5218 1382
rect 5206 1358 5210 1362
rect 5198 1348 5202 1352
rect 5254 1458 5258 1462
rect 5238 1378 5242 1382
rect 5230 1358 5234 1362
rect 5182 1328 5186 1332
rect 5246 1328 5250 1332
rect 5222 1298 5226 1302
rect 5158 1288 5162 1292
rect 5190 1288 5194 1292
rect 5142 1278 5146 1282
rect 5150 1278 5154 1282
rect 5222 1278 5226 1282
rect 5070 1268 5074 1272
rect 5070 1258 5074 1262
rect 4990 1248 4994 1252
rect 4974 1228 4978 1232
rect 5014 1218 5018 1222
rect 4814 1168 4818 1172
rect 4902 1168 4906 1172
rect 4814 1128 4818 1132
rect 4766 1118 4770 1122
rect 4942 1148 4946 1152
rect 4982 1148 4986 1152
rect 4910 1138 4914 1142
rect 5062 1248 5066 1252
rect 5174 1268 5178 1272
rect 5198 1268 5202 1272
rect 5150 1258 5154 1262
rect 5190 1258 5194 1262
rect 5174 1248 5178 1252
rect 5046 1238 5050 1242
rect 5062 1238 5066 1242
rect 5142 1238 5146 1242
rect 5102 1208 5106 1212
rect 5102 1168 5106 1172
rect 5126 1168 5130 1172
rect 5118 1158 5122 1162
rect 5086 1148 5090 1152
rect 5142 1158 5146 1162
rect 5158 1158 5162 1162
rect 5174 1158 5178 1162
rect 5182 1158 5186 1162
rect 5102 1138 5106 1142
rect 5118 1138 5122 1142
rect 4910 1118 4914 1122
rect 4518 1078 4522 1082
rect 4662 1078 4666 1082
rect 4286 1058 4290 1062
rect 4286 1048 4290 1052
rect 4334 1038 4338 1042
rect 4318 1018 4322 1022
rect 4254 978 4258 982
rect 4350 1048 4354 1052
rect 4374 1058 4378 1062
rect 4390 1058 4394 1062
rect 4406 1058 4410 1062
rect 4398 1048 4402 1052
rect 4382 1038 4386 1042
rect 4494 1068 4498 1072
rect 4422 1048 4426 1052
rect 4414 1018 4418 1022
rect 4430 1038 4434 1042
rect 4486 1008 4490 1012
rect 4442 1003 4446 1007
rect 4449 1003 4453 1007
rect 4318 968 4322 972
rect 4214 948 4218 952
rect 4222 938 4226 942
rect 4126 928 4130 932
rect 4182 928 4186 932
rect 4190 928 4194 932
rect 4222 928 4226 932
rect 4174 918 4178 922
rect 4126 898 4130 902
rect 4126 878 4130 882
rect 4062 848 4066 852
rect 4254 918 4258 922
rect 4206 878 4210 882
rect 4254 868 4258 872
rect 4102 858 4106 862
rect 4182 858 4186 862
rect 4086 838 4090 842
rect 3742 768 3746 772
rect 3822 768 3826 772
rect 3662 758 3666 762
rect 3678 758 3682 762
rect 3702 758 3706 762
rect 3726 758 3730 762
rect 3638 748 3642 752
rect 3454 738 3458 742
rect 3518 738 3522 742
rect 3478 728 3482 732
rect 3582 728 3586 732
rect 3574 708 3578 712
rect 3478 698 3482 702
rect 3510 698 3514 702
rect 3710 748 3714 752
rect 3838 748 3842 752
rect 3870 748 3874 752
rect 3902 748 3906 752
rect 4022 748 4026 752
rect 4062 758 4066 762
rect 4102 758 4106 762
rect 4262 828 4266 832
rect 4302 928 4306 932
rect 4318 928 4322 932
rect 4278 918 4282 922
rect 4342 958 4346 962
rect 4398 958 4402 962
rect 4478 958 4482 962
rect 4366 938 4370 942
rect 4302 908 4306 912
rect 4334 848 4338 852
rect 4358 848 4362 852
rect 4318 828 4322 832
rect 4438 948 4442 952
rect 4470 948 4474 952
rect 4550 1068 4554 1072
rect 4566 1068 4570 1072
rect 4590 1068 4594 1072
rect 4742 1068 4746 1072
rect 4502 1058 4506 1062
rect 4518 1048 4522 1052
rect 4574 1058 4578 1062
rect 4582 1008 4586 1012
rect 4654 1038 4658 1042
rect 4606 1008 4610 1012
rect 4638 988 4642 992
rect 4614 978 4618 982
rect 4542 968 4546 972
rect 4574 968 4578 972
rect 4502 948 4506 952
rect 4518 948 4522 952
rect 4494 938 4498 942
rect 4382 928 4386 932
rect 4614 948 4618 952
rect 4654 958 4658 962
rect 4566 938 4570 942
rect 4598 928 4602 932
rect 4630 928 4634 932
rect 4646 928 4650 932
rect 4542 918 4546 922
rect 4670 1038 4674 1042
rect 4830 1058 4834 1062
rect 4862 1058 4866 1062
rect 4774 1038 4778 1042
rect 4894 1048 4898 1052
rect 4966 1128 4970 1132
rect 4954 1103 4958 1107
rect 4961 1103 4965 1107
rect 5030 1118 5034 1122
rect 5150 1148 5154 1152
rect 5158 1148 5162 1152
rect 5078 1068 5082 1072
rect 4918 1058 4922 1062
rect 4942 1058 4946 1062
rect 4982 1058 4986 1062
rect 4990 1058 4994 1062
rect 5022 1058 5026 1062
rect 5046 1058 5050 1062
rect 5158 1138 5162 1142
rect 5190 1148 5194 1152
rect 5262 1408 5266 1412
rect 5278 1368 5282 1372
rect 5262 1358 5266 1362
rect 5278 1328 5282 1332
rect 5278 1308 5282 1312
rect 5254 1298 5258 1302
rect 5262 1268 5266 1272
rect 5246 1258 5250 1262
rect 5206 1238 5210 1242
rect 5214 1208 5218 1212
rect 5262 1238 5266 1242
rect 5278 1238 5282 1242
rect 5270 1228 5274 1232
rect 5230 1218 5234 1222
rect 5246 1218 5250 1222
rect 5206 1198 5210 1202
rect 5222 1198 5226 1202
rect 5246 1178 5250 1182
rect 5206 1138 5210 1142
rect 5198 1068 5202 1072
rect 5222 1068 5226 1072
rect 5262 1078 5266 1082
rect 5278 1068 5282 1072
rect 5150 1048 5154 1052
rect 5254 1048 5258 1052
rect 5110 1038 5114 1042
rect 4710 978 4714 982
rect 4854 978 4858 982
rect 4662 948 4666 952
rect 4678 948 4682 952
rect 4694 948 4698 952
rect 4686 938 4690 942
rect 5094 968 5098 972
rect 4750 958 4754 962
rect 4718 948 4722 952
rect 4670 918 4674 922
rect 4702 918 4706 922
rect 4726 918 4730 922
rect 4782 948 4786 952
rect 4742 938 4746 942
rect 4734 908 4738 912
rect 4718 898 4722 902
rect 4734 898 4738 902
rect 4886 958 4890 962
rect 4942 958 4946 962
rect 4934 948 4938 952
rect 4982 948 4986 952
rect 5062 948 5066 952
rect 4798 938 4802 942
rect 4862 938 4866 942
rect 4870 938 4874 942
rect 4886 938 4890 942
rect 4982 938 4986 942
rect 5046 938 5050 942
rect 4790 918 4794 922
rect 4766 908 4770 912
rect 4846 928 4850 932
rect 4870 918 4874 922
rect 4886 918 4890 922
rect 4822 898 4826 902
rect 4710 888 4714 892
rect 4814 888 4818 892
rect 4462 878 4466 882
rect 4478 878 4482 882
rect 4654 878 4658 882
rect 4702 878 4706 882
rect 4718 878 4722 882
rect 4766 878 4770 882
rect 4406 868 4410 872
rect 4398 848 4402 852
rect 4374 838 4378 842
rect 4414 838 4418 842
rect 4430 828 4434 832
rect 4422 818 4426 822
rect 4270 808 4274 812
rect 4294 808 4298 812
rect 4334 808 4338 812
rect 4366 808 4370 812
rect 4390 808 4394 812
rect 4442 803 4446 807
rect 4449 803 4453 807
rect 4478 858 4482 862
rect 4510 858 4514 862
rect 4526 848 4530 852
rect 4462 798 4466 802
rect 4454 778 4458 782
rect 4294 768 4298 772
rect 4310 768 4314 772
rect 4318 768 4322 772
rect 4414 768 4418 772
rect 4198 758 4202 762
rect 4278 758 4282 762
rect 4286 748 4290 752
rect 3774 708 3778 712
rect 3814 708 3818 712
rect 3398 658 3402 662
rect 3742 678 3746 682
rect 3774 678 3778 682
rect 3806 678 3810 682
rect 3734 668 3738 672
rect 3766 668 3770 672
rect 3782 668 3786 672
rect 3486 648 3490 652
rect 3710 658 3714 662
rect 3726 658 3730 662
rect 3782 658 3786 662
rect 3702 648 3706 652
rect 3574 638 3578 642
rect 3678 638 3682 642
rect 3686 638 3690 642
rect 3574 608 3578 612
rect 3418 603 3422 607
rect 3425 603 3429 607
rect 3350 598 3354 602
rect 3694 628 3698 632
rect 3366 588 3370 592
rect 3574 588 3578 592
rect 3582 588 3586 592
rect 3262 568 3266 572
rect 3310 568 3314 572
rect 3182 558 3186 562
rect 3238 558 3242 562
rect 3270 558 3274 562
rect 3390 558 3394 562
rect 3150 548 3154 552
rect 3174 548 3178 552
rect 3206 548 3210 552
rect 3182 528 3186 532
rect 3670 578 3674 582
rect 3630 558 3634 562
rect 3646 558 3650 562
rect 3486 548 3490 552
rect 3510 548 3514 552
rect 3198 518 3202 522
rect 3166 508 3170 512
rect 3190 508 3194 512
rect 3238 518 3242 522
rect 3334 528 3338 532
rect 3750 628 3754 632
rect 3726 578 3730 582
rect 3854 688 3858 692
rect 3814 658 3818 662
rect 3838 658 3842 662
rect 3838 648 3842 652
rect 3846 648 3850 652
rect 4102 738 4106 742
rect 4150 738 4154 742
rect 3926 728 3930 732
rect 3886 678 3890 682
rect 3902 668 3906 672
rect 4126 728 4130 732
rect 3966 718 3970 722
rect 3930 703 3934 707
rect 3937 703 3941 707
rect 3974 678 3978 682
rect 3998 678 4002 682
rect 4070 678 4074 682
rect 3966 668 3970 672
rect 3934 658 3938 662
rect 3950 658 3954 662
rect 3982 658 3986 662
rect 3886 648 3890 652
rect 3894 648 3898 652
rect 3822 618 3826 622
rect 3782 598 3786 602
rect 3742 568 3746 572
rect 3766 568 3770 572
rect 3790 568 3794 572
rect 3734 558 3738 562
rect 3750 558 3754 562
rect 3654 548 3658 552
rect 3686 548 3690 552
rect 3566 538 3570 542
rect 3614 538 3618 542
rect 3670 538 3674 542
rect 3438 528 3442 532
rect 3486 528 3490 532
rect 3262 508 3266 512
rect 3342 508 3346 512
rect 3390 508 3394 512
rect 3454 498 3458 502
rect 3470 488 3474 492
rect 3310 478 3314 482
rect 3414 478 3418 482
rect 3182 468 3186 472
rect 3470 468 3474 472
rect 3502 478 3506 482
rect 2854 458 2858 462
rect 3014 458 3018 462
rect 3238 458 3242 462
rect 3246 458 3250 462
rect 3294 458 3298 462
rect 3518 458 3522 462
rect 3526 458 3530 462
rect 2854 448 2858 452
rect 2934 448 2938 452
rect 2894 438 2898 442
rect 2814 408 2818 412
rect 2838 408 2842 412
rect 2750 378 2754 382
rect 2798 378 2802 382
rect 2934 418 2938 422
rect 2734 368 2738 372
rect 2782 368 2786 372
rect 2798 368 2802 372
rect 2822 368 2826 372
rect 2630 348 2634 352
rect 2638 348 2642 352
rect 2670 348 2674 352
rect 2750 348 2754 352
rect 2606 338 2610 342
rect 2574 328 2578 332
rect 2534 318 2538 322
rect 2566 318 2570 322
rect 2574 318 2578 322
rect 2590 308 2594 312
rect 2550 288 2554 292
rect 2582 288 2586 292
rect 2542 278 2546 282
rect 2646 288 2650 292
rect 2678 288 2682 292
rect 2702 278 2706 282
rect 2494 268 2498 272
rect 2518 268 2522 272
rect 2430 258 2434 262
rect 2454 258 2458 262
rect 2510 258 2514 262
rect 2550 258 2554 262
rect 2726 328 2730 332
rect 2790 338 2794 342
rect 2846 348 2850 352
rect 2878 348 2882 352
rect 2806 318 2810 322
rect 2830 318 2834 322
rect 2758 308 2762 312
rect 2766 308 2770 312
rect 2734 298 2738 302
rect 2750 298 2754 302
rect 2774 278 2778 282
rect 2790 278 2794 282
rect 2766 268 2770 272
rect 2758 258 2762 262
rect 2462 248 2466 252
rect 2710 248 2714 252
rect 2718 248 2722 252
rect 2906 303 2910 307
rect 2913 303 2917 307
rect 2870 278 2874 282
rect 2910 278 2914 282
rect 2806 268 2810 272
rect 2902 268 2906 272
rect 2798 258 2802 262
rect 2830 258 2834 262
rect 2894 248 2898 252
rect 2830 238 2834 242
rect 2854 238 2858 242
rect 2414 228 2418 232
rect 2614 218 2618 222
rect 2394 203 2398 207
rect 2401 203 2405 207
rect 2302 198 2306 202
rect 2318 198 2322 202
rect 2310 18 2314 22
rect 2294 8 2298 12
rect 2358 188 2362 192
rect 2542 188 2546 192
rect 2630 188 2634 192
rect 2654 188 2658 192
rect 2686 188 2690 192
rect 2430 178 2434 182
rect 2326 158 2330 162
rect 2390 138 2394 142
rect 2390 128 2394 132
rect 2366 98 2370 102
rect 2486 168 2490 172
rect 2478 148 2482 152
rect 2558 158 2562 162
rect 2590 158 2594 162
rect 2678 158 2682 162
rect 2750 188 2754 192
rect 2710 158 2714 162
rect 2742 158 2746 162
rect 2878 208 2882 212
rect 2870 188 2874 192
rect 2822 158 2826 162
rect 2862 158 2866 162
rect 2766 148 2770 152
rect 2710 138 2714 142
rect 2534 128 2538 132
rect 2598 128 2602 132
rect 2462 118 2466 122
rect 2438 108 2442 112
rect 2502 108 2506 112
rect 2526 98 2530 102
rect 2446 88 2450 92
rect 2446 78 2450 82
rect 2494 78 2498 82
rect 2614 118 2618 122
rect 2622 118 2626 122
rect 2702 118 2706 122
rect 2662 108 2666 112
rect 2734 138 2738 142
rect 2782 138 2786 142
rect 2758 128 2762 132
rect 2750 118 2754 122
rect 2790 118 2794 122
rect 2702 98 2706 102
rect 2726 98 2730 102
rect 2742 98 2746 102
rect 2670 78 2674 82
rect 2686 78 2690 82
rect 2694 78 2698 82
rect 2590 68 2594 72
rect 2678 68 2682 72
rect 2510 58 2514 62
rect 2534 59 2538 63
rect 2406 48 2410 52
rect 2358 8 2362 12
rect 2446 8 2450 12
rect 2394 3 2398 7
rect 2401 3 2405 7
rect 2670 58 2674 62
rect 2726 58 2730 62
rect 2774 108 2778 112
rect 2758 78 2762 82
rect 2646 48 2650 52
rect 2758 48 2762 52
rect 2790 98 2794 102
rect 2918 188 2922 192
rect 2886 148 2890 152
rect 2902 148 2906 152
rect 2814 138 2818 142
rect 2830 138 2834 142
rect 2838 138 2842 142
rect 2862 138 2866 142
rect 2870 138 2874 142
rect 2822 118 2826 122
rect 2846 118 2850 122
rect 2782 78 2786 82
rect 2998 388 3002 392
rect 3262 398 3266 402
rect 3446 448 3450 452
rect 3478 448 3482 452
rect 3510 448 3514 452
rect 3582 528 3586 532
rect 3598 528 3602 532
rect 3766 558 3770 562
rect 3782 548 3786 552
rect 3758 538 3762 542
rect 3678 528 3682 532
rect 3718 528 3722 532
rect 3670 518 3674 522
rect 3558 488 3562 492
rect 3574 478 3578 482
rect 3590 478 3594 482
rect 3566 458 3570 462
rect 3654 498 3658 502
rect 3638 488 3642 492
rect 3702 508 3706 512
rect 3694 468 3698 472
rect 3654 458 3658 462
rect 3662 458 3666 462
rect 3678 458 3682 462
rect 3550 448 3554 452
rect 3710 448 3714 452
rect 3486 438 3490 442
rect 3526 438 3530 442
rect 3418 403 3422 407
rect 3425 403 3429 407
rect 3342 378 3346 382
rect 3182 368 3186 372
rect 3334 368 3338 372
rect 3102 348 3106 352
rect 3134 348 3138 352
rect 3166 348 3170 352
rect 2958 328 2962 332
rect 3006 318 3010 322
rect 3078 318 3082 322
rect 3062 298 3066 302
rect 3006 288 3010 292
rect 3038 288 3042 292
rect 2974 278 2978 282
rect 3014 278 3018 282
rect 2950 268 2954 272
rect 3006 258 3010 262
rect 3086 298 3090 302
rect 3102 328 3106 332
rect 3150 318 3154 322
rect 3102 298 3106 302
rect 3070 288 3074 292
rect 3094 268 3098 272
rect 3038 258 3042 262
rect 3070 258 3074 262
rect 3086 258 3090 262
rect 3118 258 3122 262
rect 2942 248 2946 252
rect 3206 308 3210 312
rect 3142 298 3146 302
rect 3270 298 3274 302
rect 3302 298 3306 302
rect 3270 288 3274 292
rect 3310 288 3314 292
rect 3254 278 3258 282
rect 3238 258 3242 262
rect 3246 258 3250 262
rect 3246 248 3250 252
rect 3262 248 3266 252
rect 3158 238 3162 242
rect 3214 238 3218 242
rect 3126 218 3130 222
rect 3022 208 3026 212
rect 2998 198 3002 202
rect 2950 188 2954 192
rect 2958 158 2962 162
rect 3006 188 3010 192
rect 2894 128 2898 132
rect 2926 108 2930 112
rect 2906 103 2910 107
rect 2913 103 2917 107
rect 2934 98 2938 102
rect 2870 78 2874 82
rect 2798 68 2802 72
rect 2806 68 2810 72
rect 2822 68 2826 72
rect 2830 68 2834 72
rect 2846 68 2850 72
rect 2854 68 2858 72
rect 2894 68 2898 72
rect 2918 68 2922 72
rect 2854 58 2858 62
rect 2702 38 2706 42
rect 2710 28 2714 32
rect 2558 8 2562 12
rect 2926 8 2930 12
rect 2950 148 2954 152
rect 2966 148 2970 152
rect 2998 148 3002 152
rect 3062 208 3066 212
rect 3046 158 3050 162
rect 2974 138 2978 142
rect 3022 138 3026 142
rect 3142 168 3146 172
rect 3078 158 3082 162
rect 3286 278 3290 282
rect 3302 278 3306 282
rect 3334 328 3338 332
rect 3390 328 3394 332
rect 3366 318 3370 322
rect 3342 308 3346 312
rect 3510 428 3514 432
rect 3574 438 3578 442
rect 3622 438 3626 442
rect 3630 428 3634 432
rect 3566 358 3570 362
rect 3454 348 3458 352
rect 3470 348 3474 352
rect 3494 348 3498 352
rect 3542 348 3546 352
rect 3462 338 3466 342
rect 3326 288 3330 292
rect 3430 288 3434 292
rect 3318 278 3322 282
rect 3398 278 3402 282
rect 3382 268 3386 272
rect 3390 268 3394 272
rect 3342 258 3346 262
rect 3326 238 3330 242
rect 3270 218 3274 222
rect 3198 168 3202 172
rect 3222 168 3226 172
rect 3142 148 3146 152
rect 3158 148 3162 152
rect 3078 138 3082 142
rect 3102 138 3106 142
rect 2982 128 2986 132
rect 2990 118 2994 122
rect 3078 118 3082 122
rect 2974 78 2978 82
rect 3126 108 3130 112
rect 3038 88 3042 92
rect 3070 88 3074 92
rect 2990 68 2994 72
rect 2998 68 3002 72
rect 2974 58 2978 62
rect 3094 78 3098 82
rect 3230 158 3234 162
rect 3238 148 3242 152
rect 3246 148 3250 152
rect 3150 98 3154 102
rect 3230 128 3234 132
rect 3246 118 3250 122
rect 3214 98 3218 102
rect 3254 98 3258 102
rect 3174 88 3178 92
rect 3198 88 3202 92
rect 3198 78 3202 82
rect 3366 248 3370 252
rect 3534 328 3538 332
rect 3478 318 3482 322
rect 3542 318 3546 322
rect 3454 308 3458 312
rect 3518 308 3522 312
rect 3510 288 3514 292
rect 3446 278 3450 282
rect 3494 278 3498 282
rect 3438 268 3442 272
rect 3430 258 3434 262
rect 3438 248 3442 252
rect 3358 238 3362 242
rect 3390 238 3394 242
rect 3462 268 3466 272
rect 3478 268 3482 272
rect 3566 338 3570 342
rect 3726 488 3730 492
rect 3806 548 3810 552
rect 3798 538 3802 542
rect 3830 598 3834 602
rect 3902 638 3906 642
rect 3846 588 3850 592
rect 3854 588 3858 592
rect 3830 548 3834 552
rect 4006 668 4010 672
rect 4038 658 4042 662
rect 3958 648 3962 652
rect 3990 648 3994 652
rect 4014 648 4018 652
rect 4062 648 4066 652
rect 3878 568 3882 572
rect 3894 568 3898 572
rect 3918 568 3922 572
rect 3934 568 3938 572
rect 3870 548 3874 552
rect 3918 558 3922 562
rect 3910 548 3914 552
rect 4030 638 4034 642
rect 4094 658 4098 662
rect 4102 658 4106 662
rect 4102 648 4106 652
rect 4166 698 4170 702
rect 4150 688 4154 692
rect 4342 758 4346 762
rect 4374 758 4378 762
rect 4406 758 4410 762
rect 4430 758 4434 762
rect 4446 758 4450 762
rect 4318 748 4322 752
rect 4198 698 4202 702
rect 4230 698 4234 702
rect 4310 698 4314 702
rect 4166 678 4170 682
rect 4182 678 4186 682
rect 4134 658 4138 662
rect 4158 648 4162 652
rect 4166 648 4170 652
rect 4078 638 4082 642
rect 4110 638 4114 642
rect 4126 638 4130 642
rect 4006 628 4010 632
rect 4030 628 4034 632
rect 4054 628 4058 632
rect 4078 628 4082 632
rect 4070 598 4074 602
rect 3958 558 3962 562
rect 3934 548 3938 552
rect 3950 548 3954 552
rect 3990 548 3994 552
rect 4014 548 4018 552
rect 4038 548 4042 552
rect 3830 528 3834 532
rect 3822 518 3826 522
rect 3758 508 3762 512
rect 3774 508 3778 512
rect 3798 508 3802 512
rect 3774 498 3778 502
rect 3930 503 3934 507
rect 3937 503 3941 507
rect 3974 508 3978 512
rect 3814 488 3818 492
rect 3854 488 3858 492
rect 3726 468 3730 472
rect 3766 468 3770 472
rect 3790 468 3794 472
rect 3846 458 3850 462
rect 3894 468 3898 472
rect 3926 468 3930 472
rect 3902 458 3906 462
rect 3870 448 3874 452
rect 3870 398 3874 402
rect 3822 388 3826 392
rect 3846 388 3850 392
rect 3614 368 3618 372
rect 3718 368 3722 372
rect 3606 348 3610 352
rect 3638 358 3642 362
rect 3718 358 3722 362
rect 3822 358 3826 362
rect 3654 348 3658 352
rect 3662 348 3666 352
rect 3582 328 3586 332
rect 3614 328 3618 332
rect 3598 318 3602 322
rect 3542 298 3546 302
rect 3558 298 3562 302
rect 3582 298 3586 302
rect 3726 348 3730 352
rect 3774 328 3778 332
rect 3686 308 3690 312
rect 3670 298 3674 302
rect 3798 348 3802 352
rect 3862 348 3866 352
rect 3822 338 3826 342
rect 3934 458 3938 462
rect 3926 448 3930 452
rect 3910 438 3914 442
rect 3902 428 3906 432
rect 3878 338 3882 342
rect 3830 328 3834 332
rect 3862 328 3866 332
rect 3750 318 3754 322
rect 3766 318 3770 322
rect 3782 318 3786 322
rect 3774 298 3778 302
rect 3670 278 3674 282
rect 3846 298 3850 302
rect 3910 388 3914 392
rect 4102 598 4106 602
rect 4110 598 4114 602
rect 4110 568 4114 572
rect 4134 548 4138 552
rect 4046 538 4050 542
rect 3990 528 3994 532
rect 4014 528 4018 532
rect 4238 688 4242 692
rect 4206 668 4210 672
rect 4198 658 4202 662
rect 4382 748 4386 752
rect 4390 748 4394 752
rect 4374 728 4378 732
rect 4342 698 4346 702
rect 4398 738 4402 742
rect 4422 698 4426 702
rect 4254 668 4258 672
rect 4334 668 4338 672
rect 4366 668 4370 672
rect 4414 668 4418 672
rect 4630 868 4634 872
rect 4654 868 4658 872
rect 4694 868 4698 872
rect 4566 858 4570 862
rect 4606 858 4610 862
rect 4582 848 4586 852
rect 4606 848 4610 852
rect 4534 838 4538 842
rect 4542 838 4546 842
rect 4622 838 4626 842
rect 4478 778 4482 782
rect 4510 778 4514 782
rect 4494 768 4498 772
rect 4646 828 4650 832
rect 4606 818 4610 822
rect 4686 818 4690 822
rect 4566 808 4570 812
rect 4558 778 4562 782
rect 4758 868 4762 872
rect 4774 868 4778 872
rect 4710 818 4714 822
rect 4702 808 4706 812
rect 4790 848 4794 852
rect 4878 908 4882 912
rect 4966 928 4970 932
rect 5006 928 5010 932
rect 4974 918 4978 922
rect 4954 903 4958 907
rect 4961 903 4965 907
rect 4934 888 4938 892
rect 5030 888 5034 892
rect 4862 868 4866 872
rect 4902 868 4906 872
rect 4934 868 4938 872
rect 4846 858 4850 862
rect 4830 848 4834 852
rect 4846 848 4850 852
rect 4838 828 4842 832
rect 4678 778 4682 782
rect 4798 778 4802 782
rect 4582 768 4586 772
rect 4534 758 4538 762
rect 4558 758 4562 762
rect 4606 768 4610 772
rect 4630 768 4634 772
rect 4670 768 4674 772
rect 4678 768 4682 772
rect 4614 758 4618 762
rect 4486 748 4490 752
rect 4518 748 4522 752
rect 4574 748 4578 752
rect 4638 758 4642 762
rect 4654 748 4658 752
rect 4470 738 4474 742
rect 4478 738 4482 742
rect 4510 738 4514 742
rect 4566 738 4570 742
rect 4614 738 4618 742
rect 4646 738 4650 742
rect 4502 688 4506 692
rect 4486 678 4490 682
rect 4230 658 4234 662
rect 4246 658 4250 662
rect 4310 648 4314 652
rect 4222 638 4226 642
rect 4286 638 4290 642
rect 4182 568 4186 572
rect 4358 648 4362 652
rect 4390 648 4394 652
rect 4414 648 4418 652
rect 4566 668 4570 672
rect 4694 758 4698 762
rect 4790 758 4794 762
rect 4734 748 4738 752
rect 4710 738 4714 742
rect 4726 688 4730 692
rect 4814 768 4818 772
rect 4782 738 4786 742
rect 4854 748 4858 752
rect 4798 728 4802 732
rect 4766 698 4770 702
rect 4750 688 4754 692
rect 4894 858 4898 862
rect 4918 858 4922 862
rect 4878 848 4882 852
rect 4910 848 4914 852
rect 4894 838 4898 842
rect 4926 838 4930 842
rect 5014 858 5018 862
rect 5006 848 5010 852
rect 5014 848 5018 852
rect 5030 848 5034 852
rect 4990 838 4994 842
rect 4950 828 4954 832
rect 4870 818 4874 822
rect 4982 818 4986 822
rect 5046 928 5050 932
rect 5070 928 5074 932
rect 5126 948 5130 952
rect 5190 948 5194 952
rect 5142 928 5146 932
rect 5110 918 5114 922
rect 5118 918 5122 922
rect 5174 918 5178 922
rect 5270 1008 5274 1012
rect 5238 968 5242 972
rect 5254 958 5258 962
rect 5262 928 5266 932
rect 5278 948 5282 952
rect 5174 888 5178 892
rect 5206 888 5210 892
rect 5222 888 5226 892
rect 5262 888 5266 892
rect 5046 868 5050 872
rect 5070 858 5074 862
rect 5030 838 5034 842
rect 5014 788 5018 792
rect 4974 768 4978 772
rect 4982 758 4986 762
rect 4910 748 4914 752
rect 4926 748 4930 752
rect 4870 738 4874 742
rect 4862 718 4866 722
rect 4622 648 4626 652
rect 4942 738 4946 742
rect 4926 718 4930 722
rect 4954 703 4958 707
rect 4961 703 4965 707
rect 4998 758 5002 762
rect 5022 778 5026 782
rect 5038 728 5042 732
rect 5030 708 5034 712
rect 5046 708 5050 712
rect 4910 668 4914 672
rect 4822 658 4826 662
rect 4862 658 4866 662
rect 4886 658 4890 662
rect 5046 678 5050 682
rect 4974 668 4978 672
rect 5022 668 5026 672
rect 5054 668 5058 672
rect 5270 868 5274 872
rect 5262 858 5266 862
rect 5278 858 5282 862
rect 5230 798 5234 802
rect 5134 788 5138 792
rect 5110 778 5114 782
rect 5182 778 5186 782
rect 5142 768 5146 772
rect 5078 758 5082 762
rect 5102 758 5106 762
rect 5126 758 5130 762
rect 5150 758 5154 762
rect 5110 748 5114 752
rect 5078 728 5082 732
rect 5086 688 5090 692
rect 5126 738 5130 742
rect 5158 718 5162 722
rect 5102 678 5106 682
rect 5118 678 5122 682
rect 5198 748 5202 752
rect 5246 728 5250 732
rect 5206 688 5210 692
rect 5254 678 5258 682
rect 5230 668 5234 672
rect 4942 658 4946 662
rect 4982 658 4986 662
rect 5102 658 5106 662
rect 5158 658 5162 662
rect 4918 648 4922 652
rect 4966 648 4970 652
rect 4654 638 4658 642
rect 4694 638 4698 642
rect 4718 638 4722 642
rect 4742 638 4746 642
rect 4878 638 4882 642
rect 5270 618 5274 622
rect 4430 608 4434 612
rect 4442 603 4446 607
rect 4449 603 4453 607
rect 4334 598 4338 602
rect 4166 548 4170 552
rect 4190 548 4194 552
rect 4278 548 4282 552
rect 4310 548 4314 552
rect 4350 548 4354 552
rect 4190 538 4194 542
rect 4142 528 4146 532
rect 4166 528 4170 532
rect 4046 518 4050 522
rect 4054 518 4058 522
rect 3990 498 3994 502
rect 4006 498 4010 502
rect 4110 498 4114 502
rect 4046 488 4050 492
rect 4070 488 4074 492
rect 4102 488 4106 492
rect 3982 478 3986 482
rect 3998 478 4002 482
rect 4054 468 4058 472
rect 3974 448 3978 452
rect 4006 448 4010 452
rect 3966 438 3970 442
rect 3982 438 3986 442
rect 4014 438 4018 442
rect 3958 428 3962 432
rect 3974 368 3978 372
rect 3990 348 3994 352
rect 4006 348 4010 352
rect 3974 338 3978 342
rect 3998 328 4002 332
rect 4142 498 4146 502
rect 4134 488 4138 492
rect 4094 468 4098 472
rect 4134 468 4138 472
rect 4086 458 4090 462
rect 4214 538 4218 542
rect 4262 538 4266 542
rect 4278 538 4282 542
rect 4198 528 4202 532
rect 4270 528 4274 532
rect 4302 528 4306 532
rect 4326 518 4330 522
rect 4334 518 4338 522
rect 4246 508 4250 512
rect 5278 588 5282 592
rect 5078 578 5082 582
rect 5142 578 5146 582
rect 4518 568 4522 572
rect 4542 568 4546 572
rect 4566 568 4570 572
rect 4598 568 4602 572
rect 4526 548 4530 552
rect 4222 498 4226 502
rect 4158 458 4162 462
rect 4438 478 4442 482
rect 4550 548 4554 552
rect 4590 548 4594 552
rect 4814 558 4818 562
rect 4622 548 4626 552
rect 4638 548 4642 552
rect 4678 548 4682 552
rect 4694 548 4698 552
rect 4606 538 4610 542
rect 4646 528 4650 532
rect 4550 498 4554 502
rect 4502 488 4506 492
rect 4534 488 4538 492
rect 4486 478 4490 482
rect 4214 458 4218 462
rect 4126 448 4130 452
rect 4174 448 4178 452
rect 4062 438 4066 442
rect 4022 398 4026 402
rect 4166 438 4170 442
rect 4150 428 4154 432
rect 4270 418 4274 422
rect 4302 448 4306 452
rect 4382 458 4386 462
rect 4518 478 4522 482
rect 4494 458 4498 462
rect 4518 458 4522 462
rect 4382 448 4386 452
rect 4446 448 4450 452
rect 4614 488 4618 492
rect 4622 488 4626 492
rect 4638 488 4642 492
rect 4662 488 4666 492
rect 4710 488 4714 492
rect 4590 478 4594 482
rect 4606 468 4610 472
rect 4558 458 4562 462
rect 4574 458 4578 462
rect 4550 448 4554 452
rect 4358 438 4362 442
rect 4390 438 4394 442
rect 4454 438 4458 442
rect 4566 438 4570 442
rect 4318 418 4322 422
rect 4278 408 4282 412
rect 4406 408 4410 412
rect 4442 403 4446 407
rect 4449 403 4453 407
rect 4078 388 4082 392
rect 4214 388 4218 392
rect 4030 368 4034 372
rect 4086 358 4090 362
rect 4022 338 4026 342
rect 4038 338 4042 342
rect 3990 318 3994 322
rect 4014 318 4018 322
rect 4062 338 4066 342
rect 4422 378 4426 382
rect 4454 378 4458 382
rect 4238 348 4242 352
rect 4278 348 4282 352
rect 4382 368 4386 372
rect 4406 348 4410 352
rect 4542 398 4546 402
rect 4502 378 4506 382
rect 4526 378 4530 382
rect 4502 368 4506 372
rect 4518 358 4522 362
rect 4502 348 4506 352
rect 4598 448 4602 452
rect 4654 478 4658 482
rect 4670 468 4674 472
rect 4638 458 4642 462
rect 4662 458 4666 462
rect 4614 438 4618 442
rect 4598 378 4602 382
rect 4566 358 4570 362
rect 4678 448 4682 452
rect 4670 418 4674 422
rect 4646 398 4650 402
rect 4638 378 4642 382
rect 4646 378 4650 382
rect 4606 358 4610 362
rect 4102 338 4106 342
rect 4486 338 4490 342
rect 4542 338 4546 342
rect 4574 338 4578 342
rect 4622 338 4626 342
rect 4054 318 4058 322
rect 4078 318 4082 322
rect 3930 303 3934 307
rect 3937 303 3941 307
rect 4006 298 4010 302
rect 4118 318 4122 322
rect 4142 318 4146 322
rect 4334 328 4338 332
rect 4310 318 4314 322
rect 4350 318 4354 322
rect 4182 308 4186 312
rect 4134 298 4138 302
rect 4214 288 4218 292
rect 4254 288 4258 292
rect 3582 268 3586 272
rect 3638 268 3642 272
rect 3726 268 3730 272
rect 3750 268 3754 272
rect 4006 268 4010 272
rect 4118 268 4122 272
rect 4166 268 4170 272
rect 4238 268 4242 272
rect 3486 258 3490 262
rect 3670 258 3674 262
rect 3726 258 3730 262
rect 3758 258 3762 262
rect 3830 258 3834 262
rect 3870 258 3874 262
rect 3934 258 3938 262
rect 4110 258 4114 262
rect 3526 248 3530 252
rect 3630 248 3634 252
rect 3646 248 3650 252
rect 3814 248 3818 252
rect 4038 248 4042 252
rect 3910 238 3914 242
rect 3718 218 3722 222
rect 3350 198 3354 202
rect 3278 188 3282 192
rect 3310 168 3314 172
rect 3326 168 3330 172
rect 3418 203 3422 207
rect 3425 203 3429 207
rect 3358 158 3362 162
rect 3406 158 3410 162
rect 3462 158 3466 162
rect 3278 108 3282 112
rect 3622 188 3626 192
rect 3638 188 3642 192
rect 3526 168 3530 172
rect 3566 168 3570 172
rect 3438 148 3442 152
rect 3686 178 3690 182
rect 3654 168 3658 172
rect 3710 168 3714 172
rect 3574 158 3578 162
rect 3630 158 3634 162
rect 3702 158 3706 162
rect 3350 138 3354 142
rect 3374 138 3378 142
rect 3462 138 3466 142
rect 3486 138 3490 142
rect 3518 138 3522 142
rect 3558 138 3562 142
rect 3366 128 3370 132
rect 3382 128 3386 132
rect 3406 128 3410 132
rect 3326 118 3330 122
rect 3454 118 3458 122
rect 3382 98 3386 102
rect 3390 98 3394 102
rect 3430 98 3434 102
rect 3310 88 3314 92
rect 3278 78 3282 82
rect 3286 78 3290 82
rect 3358 78 3362 82
rect 3366 78 3370 82
rect 3134 68 3138 72
rect 3150 68 3154 72
rect 3174 68 3178 72
rect 3190 68 3194 72
rect 3318 68 3322 72
rect 3342 68 3346 72
rect 3422 68 3426 72
rect 3214 58 3218 62
rect 3086 48 3090 52
rect 3118 48 3122 52
rect 2982 38 2986 42
rect 3006 38 3010 42
rect 3014 38 3018 42
rect 3142 38 3146 42
rect 3438 88 3442 92
rect 3454 78 3458 82
rect 3590 138 3594 142
rect 3638 148 3642 152
rect 3702 148 3706 152
rect 3622 138 3626 142
rect 3654 138 3658 142
rect 3710 138 3714 142
rect 3486 128 3490 132
rect 3518 128 3522 132
rect 3582 128 3586 132
rect 3598 128 3602 132
rect 3470 118 3474 122
rect 3478 118 3482 122
rect 3534 118 3538 122
rect 3502 108 3506 112
rect 3502 88 3506 92
rect 3526 78 3530 82
rect 3462 68 3466 72
rect 3550 68 3554 72
rect 3886 228 3890 232
rect 3790 188 3794 192
rect 3742 178 3746 182
rect 3766 178 3770 182
rect 3750 168 3754 172
rect 3742 158 3746 162
rect 3734 138 3738 142
rect 3774 168 3778 172
rect 3798 168 3802 172
rect 3822 168 3826 172
rect 3822 158 3826 162
rect 3942 178 3946 182
rect 3790 148 3794 152
rect 3822 148 3826 152
rect 3782 138 3786 142
rect 3822 138 3826 142
rect 3886 138 3890 142
rect 3606 118 3610 122
rect 3686 118 3690 122
rect 3774 118 3778 122
rect 3718 98 3722 102
rect 3606 88 3610 92
rect 3630 88 3634 92
rect 3646 88 3650 92
rect 3574 78 3578 82
rect 3614 78 3618 82
rect 3662 78 3666 82
rect 3622 68 3626 72
rect 3646 68 3650 72
rect 3710 68 3714 72
rect 3598 58 3602 62
rect 3638 58 3642 62
rect 3694 58 3698 62
rect 3302 48 3306 52
rect 3350 48 3354 52
rect 3590 48 3594 52
rect 3734 68 3738 72
rect 3758 68 3762 72
rect 3734 48 3738 52
rect 3822 128 3826 132
rect 3798 98 3802 102
rect 3814 88 3818 92
rect 3822 88 3826 92
rect 3846 88 3850 92
rect 3822 78 3826 82
rect 3878 78 3882 82
rect 3782 66 3786 70
rect 3886 58 3890 62
rect 3758 48 3762 52
rect 3766 48 3770 52
rect 3814 48 3818 52
rect 3822 48 3826 52
rect 3854 48 3858 52
rect 3870 48 3874 52
rect 3494 38 3498 42
rect 3678 38 3682 42
rect 3702 38 3706 42
rect 3718 38 3722 42
rect 3742 38 3746 42
rect 3286 28 3290 32
rect 3006 18 3010 22
rect 3982 138 3986 142
rect 3918 128 3922 132
rect 3918 118 3922 122
rect 3910 98 3914 102
rect 3930 103 3934 107
rect 3937 103 3941 107
rect 3934 88 3938 92
rect 3982 98 3986 102
rect 3918 58 3922 62
rect 2982 8 2986 12
rect 3006 8 3010 12
rect 3086 8 3090 12
rect 3182 8 3186 12
rect 3342 8 3346 12
rect 3502 8 3506 12
rect 3558 8 3562 12
rect 3718 8 3722 12
rect 3878 8 3882 12
rect 3902 8 3906 12
rect 3418 3 3422 7
rect 3425 3 3429 7
rect 4126 258 4130 262
rect 4246 258 4250 262
rect 4102 248 4106 252
rect 4278 248 4282 252
rect 4294 248 4298 252
rect 4094 198 4098 202
rect 4350 288 4354 292
rect 4534 328 4538 332
rect 4582 328 4586 332
rect 4510 318 4514 322
rect 4614 288 4618 292
rect 4494 278 4498 282
rect 4318 258 4322 262
rect 4590 278 4594 282
rect 4638 278 4642 282
rect 4662 348 4666 352
rect 4742 478 4746 482
rect 4846 548 4850 552
rect 4862 558 4866 562
rect 4870 548 4874 552
rect 4886 548 4890 552
rect 4902 548 4906 552
rect 5006 548 5010 552
rect 4838 538 4842 542
rect 4854 538 4858 542
rect 4958 538 4962 542
rect 5118 548 5122 552
rect 5174 568 5178 572
rect 5302 1278 5306 1282
rect 5302 868 5306 872
rect 5238 558 5242 562
rect 5214 548 5218 552
rect 4862 498 4866 502
rect 4822 478 4826 482
rect 4846 478 4850 482
rect 4718 468 4722 472
rect 4766 468 4770 472
rect 4790 468 4794 472
rect 4694 418 4698 422
rect 4686 408 4690 412
rect 4702 378 4706 382
rect 4686 368 4690 372
rect 4726 458 4730 462
rect 4862 468 4866 472
rect 4894 468 4898 472
rect 4806 458 4810 462
rect 4718 448 4722 452
rect 4750 448 4754 452
rect 4798 448 4802 452
rect 4758 428 4762 432
rect 4870 428 4874 432
rect 4886 428 4890 432
rect 4854 408 4858 412
rect 4954 503 4958 507
rect 4961 503 4965 507
rect 5070 498 5074 502
rect 5094 498 5098 502
rect 5030 488 5034 492
rect 5054 478 5058 482
rect 4950 468 4954 472
rect 5006 468 5010 472
rect 5030 468 5034 472
rect 4958 458 4962 462
rect 4982 458 4986 462
rect 4926 448 4930 452
rect 4934 438 4938 442
rect 4998 438 5002 442
rect 5014 438 5018 442
rect 5038 438 5042 442
rect 5086 488 5090 492
rect 5078 478 5082 482
rect 5126 468 5130 472
rect 5278 548 5282 552
rect 5278 538 5282 542
rect 5294 538 5298 542
rect 5070 458 5074 462
rect 5174 458 5178 462
rect 5134 448 5138 452
rect 5166 448 5170 452
rect 5054 438 5058 442
rect 5142 438 5146 442
rect 4934 418 4938 422
rect 4742 388 4746 392
rect 5014 408 5018 412
rect 4910 378 4914 382
rect 4966 378 4970 382
rect 4982 378 4986 382
rect 5142 378 5146 382
rect 4934 368 4938 372
rect 4686 358 4690 362
rect 4710 358 4714 362
rect 4894 358 4898 362
rect 4902 358 4906 362
rect 4966 358 4970 362
rect 4726 348 4730 352
rect 4798 348 4802 352
rect 4678 338 4682 342
rect 4694 338 4698 342
rect 4702 328 4706 332
rect 4678 288 4682 292
rect 4686 288 4690 292
rect 4662 268 4666 272
rect 4462 258 4466 262
rect 4558 258 4562 262
rect 4614 258 4618 262
rect 4374 248 4378 252
rect 4310 238 4314 242
rect 4134 188 4138 192
rect 4158 188 4162 192
rect 4302 188 4306 192
rect 4214 168 4218 172
rect 4198 158 4202 162
rect 4094 151 4098 152
rect 4094 148 4098 151
rect 4102 148 4106 152
rect 4054 138 4058 142
rect 4166 118 4170 122
rect 4102 88 4106 92
rect 4166 78 4170 82
rect 4126 68 4130 72
rect 4214 68 4218 72
rect 4046 8 4050 12
rect 4094 8 4098 12
rect 4190 8 4194 12
rect 4342 178 4346 182
rect 4398 168 4402 172
rect 4342 148 4346 152
rect 4358 148 4362 152
rect 4502 248 4506 252
rect 4442 203 4446 207
rect 4449 203 4453 207
rect 4430 158 4434 162
rect 4646 248 4650 252
rect 4710 298 4714 302
rect 4694 268 4698 272
rect 4710 268 4714 272
rect 4838 348 4842 352
rect 4862 348 4866 352
rect 4910 348 4914 352
rect 4806 338 4810 342
rect 4822 340 4826 344
rect 4854 338 4858 342
rect 4782 328 4786 332
rect 4790 328 4794 332
rect 4774 318 4778 322
rect 4798 318 4802 322
rect 4758 298 4762 302
rect 4734 278 4738 282
rect 4726 268 4730 272
rect 4686 248 4690 252
rect 4662 238 4666 242
rect 4678 238 4682 242
rect 4590 148 4594 152
rect 4686 178 4690 182
rect 4678 168 4682 172
rect 4710 168 4714 172
rect 4798 268 4802 272
rect 4862 328 4866 332
rect 4942 348 4946 352
rect 4966 348 4970 352
rect 4990 368 4994 372
rect 5038 368 5042 372
rect 5006 358 5010 362
rect 5022 348 5026 352
rect 4982 338 4986 342
rect 5006 338 5010 342
rect 4926 328 4930 332
rect 4954 303 4958 307
rect 4961 303 4965 307
rect 4870 298 4874 302
rect 4894 288 4898 292
rect 4814 278 4818 282
rect 4862 278 4866 282
rect 4886 278 4890 282
rect 4990 278 4994 282
rect 5246 448 5250 452
rect 5270 358 5274 362
rect 5046 348 5050 352
rect 5110 348 5114 352
rect 5134 348 5138 352
rect 5174 348 5178 352
rect 5078 338 5082 342
rect 5086 328 5090 332
rect 5110 328 5114 332
rect 5142 328 5146 332
rect 5190 328 5194 332
rect 4750 258 4754 262
rect 4774 258 4778 262
rect 4822 258 4826 262
rect 4902 268 4906 272
rect 4958 268 4962 272
rect 4990 268 4994 272
rect 4758 248 4762 252
rect 4774 248 4778 252
rect 4838 248 4842 252
rect 4726 238 4730 242
rect 4702 158 4706 162
rect 4718 158 4722 162
rect 4734 178 4738 182
rect 4646 138 4650 142
rect 4262 118 4266 122
rect 4294 108 4298 112
rect 4334 98 4338 102
rect 4254 88 4258 92
rect 4318 88 4322 92
rect 4270 78 4274 82
rect 4302 78 4306 82
rect 4286 68 4290 72
rect 4318 68 4322 72
rect 4294 58 4298 62
rect 4406 118 4410 122
rect 4438 108 4442 112
rect 4486 108 4490 112
rect 4374 98 4378 102
rect 4350 88 4354 92
rect 4622 118 4626 122
rect 4558 108 4562 112
rect 4862 238 4866 242
rect 4910 258 4914 262
rect 4926 258 4930 262
rect 4926 248 4930 252
rect 5038 278 5042 282
rect 5062 278 5066 282
rect 5046 268 5050 272
rect 5078 268 5082 272
rect 5214 298 5218 302
rect 5134 288 5138 292
rect 5206 288 5210 292
rect 5214 288 5218 292
rect 5166 278 5170 282
rect 5182 278 5186 282
rect 5110 268 5114 272
rect 5134 268 5138 272
rect 5150 268 5154 272
rect 5222 268 5226 272
rect 5094 258 5098 262
rect 5126 258 5130 262
rect 5158 258 5162 262
rect 4950 238 4954 242
rect 5006 238 5010 242
rect 5014 238 5018 242
rect 4894 228 4898 232
rect 4910 228 4914 232
rect 5014 218 5018 222
rect 5086 228 5090 232
rect 5046 198 5050 202
rect 5070 198 5074 202
rect 4878 188 4882 192
rect 4798 178 4802 182
rect 5062 178 5066 182
rect 4766 168 4770 172
rect 4782 158 4786 162
rect 4846 168 4850 172
rect 5070 168 5074 172
rect 5102 238 5106 242
rect 5102 168 5106 172
rect 4814 158 4818 162
rect 4878 158 4882 162
rect 4886 158 4890 162
rect 4926 158 4930 162
rect 4942 158 4946 162
rect 4774 148 4778 152
rect 4790 148 4794 152
rect 4838 148 4842 152
rect 4678 138 4682 142
rect 4742 138 4746 142
rect 4806 138 4810 142
rect 4838 138 4842 142
rect 4862 138 4866 142
rect 4710 128 4714 132
rect 4766 128 4770 132
rect 4718 118 4722 122
rect 4774 118 4778 122
rect 4494 98 4498 102
rect 4534 98 4538 102
rect 4606 98 4610 102
rect 4982 138 4986 142
rect 4918 128 4922 132
rect 4934 128 4938 132
rect 4954 103 4958 107
rect 4961 103 4965 107
rect 5094 148 5098 152
rect 4998 138 5002 142
rect 5126 148 5130 152
rect 5142 148 5146 152
rect 5078 138 5082 142
rect 5102 138 5106 142
rect 5142 138 5146 142
rect 4998 118 5002 122
rect 4558 88 4562 92
rect 4638 88 4642 92
rect 4918 88 4922 92
rect 4982 88 4986 92
rect 4990 88 4994 92
rect 5030 88 5034 92
rect 5038 88 5042 92
rect 5086 88 5090 92
rect 4654 78 4658 82
rect 5006 78 5010 82
rect 5062 78 5066 82
rect 5094 78 5098 82
rect 4334 68 4338 72
rect 4558 68 4562 72
rect 4358 58 4362 62
rect 4414 58 4418 62
rect 4294 48 4298 52
rect 4470 48 4474 52
rect 4390 38 4394 42
rect 4422 8 4426 12
rect 4486 8 4490 12
rect 4442 3 4446 7
rect 4449 3 4453 7
rect 4766 58 4770 62
rect 4798 58 4802 62
rect 4902 48 4906 52
rect 5214 148 5218 152
rect 5174 138 5178 142
rect 5158 88 5162 92
rect 5206 68 5210 72
rect 5118 58 5122 62
rect 5030 48 5034 52
rect 5038 48 5042 52
rect 5070 48 5074 52
rect 5086 48 5090 52
rect 5358 588 5362 592
rect 5286 368 5290 372
rect 5286 348 5290 352
rect 5270 328 5274 332
rect 5278 328 5282 332
rect 5246 268 5250 272
rect 5262 268 5266 272
rect 5294 338 5298 342
rect 5294 318 5298 322
rect 5246 258 5250 262
rect 5278 238 5282 242
rect 5270 188 5274 192
rect 5270 148 5274 152
rect 5238 138 5242 142
rect 5294 78 5298 82
rect 5270 58 5274 62
rect 5294 58 5298 62
rect 5246 8 5250 12
<< metal3 >>
rect 856 3703 858 3707
rect 862 3703 865 3707
rect 870 3703 872 3707
rect 1872 3703 1874 3707
rect 1878 3703 1881 3707
rect 1886 3703 1888 3707
rect 2904 3703 2906 3707
rect 2910 3703 2913 3707
rect 2918 3703 2920 3707
rect 3928 3703 3930 3707
rect 3934 3703 3937 3707
rect 3942 3703 3944 3707
rect 4952 3703 4954 3707
rect 4958 3703 4961 3707
rect 4966 3703 4968 3707
rect 522 3698 558 3701
rect 562 3698 694 3701
rect 1954 3698 1982 3701
rect 2178 3698 2206 3701
rect 2698 3698 2718 3701
rect 3962 3698 3974 3701
rect 3994 3698 3998 3701
rect 4074 3698 4078 3701
rect 4210 3698 4214 3701
rect 4370 3698 4374 3701
rect 5242 3698 5246 3701
rect 3286 3692 3289 3698
rect 4238 3692 4241 3698
rect 4294 3692 4297 3698
rect 490 3688 1078 3691
rect 1106 3688 1214 3691
rect 1738 3688 1742 3691
rect 1778 3688 2230 3691
rect 2234 3688 2254 3691
rect 2274 3688 2278 3691
rect 2690 3688 2710 3691
rect 3810 3688 3862 3691
rect 4090 3688 4182 3691
rect 4346 3688 4374 3691
rect 5066 3688 5150 3691
rect 294 3681 297 3688
rect 294 3678 422 3681
rect 426 3678 446 3681
rect 458 3678 478 3681
rect 546 3678 566 3681
rect 834 3678 942 3681
rect 954 3678 982 3681
rect 986 3678 1046 3681
rect 1222 3681 1225 3688
rect 1222 3678 1294 3681
rect 1626 3678 1670 3681
rect 1698 3678 1742 3681
rect 1826 3678 1966 3681
rect 1986 3678 2097 3681
rect 2258 3678 2286 3681
rect 2310 3681 2313 3688
rect 2298 3678 2313 3681
rect 2458 3678 2470 3681
rect 2550 3681 2553 3688
rect 2638 3681 2641 3688
rect 2550 3678 2641 3681
rect 3066 3678 3110 3681
rect 3218 3678 3318 3681
rect 3730 3678 3854 3681
rect 4058 3678 4102 3681
rect 4194 3678 4446 3681
rect 4666 3678 4710 3681
rect 4730 3678 4734 3681
rect 4850 3678 4894 3681
rect 414 3668 465 3671
rect 622 3671 625 3678
rect 610 3668 726 3671
rect 734 3671 737 3678
rect 734 3668 782 3671
rect 786 3668 910 3671
rect 914 3668 958 3671
rect 978 3668 990 3671
rect 1370 3668 1425 3671
rect 1482 3668 1502 3671
rect 1598 3671 1601 3678
rect 2094 3672 2097 3678
rect 1598 3668 1630 3671
rect 1650 3668 1742 3671
rect 1794 3668 1801 3671
rect 1890 3668 1910 3671
rect 1914 3668 1982 3671
rect 2098 3668 2190 3671
rect 2194 3668 2214 3671
rect 2250 3668 2270 3671
rect 2274 3668 2358 3671
rect 2442 3668 2654 3671
rect 2658 3668 2678 3671
rect 2922 3668 3118 3671
rect 3122 3668 3326 3671
rect 3330 3668 3462 3671
rect 3674 3668 3742 3671
rect 3962 3668 4094 3671
rect 4306 3668 4422 3671
rect 4562 3668 4702 3671
rect 4998 3671 5001 3678
rect 4834 3668 4897 3671
rect 4998 3668 5038 3671
rect 414 3662 417 3668
rect 462 3662 465 3668
rect 618 3658 654 3661
rect 658 3658 670 3661
rect 850 3658 878 3661
rect 942 3658 950 3661
rect 954 3658 977 3661
rect 1002 3658 1046 3661
rect 1050 3658 1206 3661
rect 1238 3661 1241 3668
rect 1422 3662 1425 3668
rect 1798 3662 1801 3668
rect 1218 3658 1241 3661
rect 1306 3658 1334 3661
rect 1434 3658 1518 3661
rect 1522 3658 1566 3661
rect 1586 3658 1654 3661
rect 1738 3658 1742 3661
rect 1850 3658 1862 3661
rect 1866 3658 1934 3661
rect 1962 3658 1998 3661
rect 2106 3658 2118 3661
rect 2122 3658 2142 3661
rect 2274 3658 2294 3661
rect 2306 3658 2318 3661
rect 2322 3658 2398 3661
rect 2402 3658 2462 3661
rect 2514 3658 2518 3661
rect 2522 3658 2542 3661
rect 2650 3658 2742 3661
rect 2838 3658 2870 3661
rect 2914 3658 3094 3661
rect 3114 3658 3150 3661
rect 3370 3658 3374 3661
rect 3658 3658 3694 3661
rect 3850 3658 4086 3661
rect 4178 3658 4241 3661
rect 4330 3658 4366 3661
rect 4434 3658 4446 3661
rect 4534 3661 4537 3668
rect 4894 3662 4897 3668
rect 4514 3658 4537 3661
rect 4770 3658 4782 3661
rect 4986 3658 5097 3661
rect 5178 3658 5254 3661
rect 310 3651 313 3658
rect 258 3648 313 3651
rect 634 3648 654 3651
rect 658 3648 758 3651
rect 798 3651 801 3658
rect 778 3648 801 3651
rect 822 3651 825 3658
rect 974 3652 977 3658
rect 2838 3652 2841 3658
rect 4086 3652 4089 3658
rect 4238 3652 4241 3658
rect 5094 3652 5097 3658
rect 822 3648 945 3651
rect 1034 3648 1142 3651
rect 1146 3648 1150 3651
rect 1162 3648 1230 3651
rect 1402 3648 1430 3651
rect 1438 3648 1502 3651
rect 1522 3648 1529 3651
rect 1554 3648 1606 3651
rect 1610 3648 1614 3651
rect 1626 3648 1630 3651
rect 1634 3648 1646 3651
rect 1730 3648 1822 3651
rect 1842 3648 1854 3651
rect 1858 3648 1902 3651
rect 2134 3648 2174 3651
rect 2242 3648 2342 3651
rect 2362 3648 2390 3651
rect 2426 3648 2446 3651
rect 2498 3648 2534 3651
rect 2538 3648 2558 3651
rect 2906 3648 3118 3651
rect 3122 3648 3326 3651
rect 3562 3648 3750 3651
rect 3826 3648 4006 3651
rect 4114 3648 4182 3651
rect 4362 3648 4398 3651
rect 4578 3648 4598 3651
rect 4722 3648 4902 3651
rect 4906 3648 4990 3651
rect 5018 3648 5030 3651
rect 5242 3648 5246 3651
rect 5282 3648 5310 3651
rect 5342 3651 5346 3652
rect 5314 3648 5346 3651
rect 942 3642 945 3648
rect 178 3638 262 3641
rect 266 3638 286 3641
rect 594 3638 657 3641
rect 794 3638 806 3641
rect 1286 3641 1289 3648
rect 1438 3642 1441 3648
rect 1526 3642 1529 3648
rect 1274 3638 1289 3641
rect 1298 3638 1326 3641
rect 1530 3638 1726 3641
rect 1746 3638 1806 3641
rect 1810 3638 1830 3641
rect 1850 3638 1854 3641
rect 2062 3641 2065 3648
rect 2134 3642 2137 3648
rect 2062 3638 2110 3641
rect 2138 3638 2302 3641
rect 2322 3638 2326 3641
rect 2342 3641 2345 3648
rect 2342 3638 2374 3641
rect 2482 3638 2486 3641
rect 2858 3638 3078 3641
rect 3082 3638 3222 3641
rect 3758 3641 3761 3648
rect 3586 3638 3761 3641
rect 3866 3638 3950 3641
rect 3970 3638 3982 3641
rect 4074 3638 4246 3641
rect 4354 3638 4390 3641
rect 4394 3638 4462 3641
rect 4506 3638 4526 3641
rect 4530 3638 4766 3641
rect 322 3628 350 3631
rect 354 3628 406 3631
rect 410 3628 606 3631
rect 610 3628 622 3631
rect 626 3628 638 3631
rect 654 3631 657 3638
rect 654 3628 822 3631
rect 898 3628 1126 3631
rect 1226 3628 2054 3631
rect 2058 3628 2190 3631
rect 2342 3628 2430 3631
rect 2434 3628 2462 3631
rect 2478 3628 2486 3631
rect 2490 3628 2662 3631
rect 2786 3628 3078 3631
rect 3498 3628 3654 3631
rect 3914 3628 4414 3631
rect 4682 3628 4814 3631
rect 4818 3628 5078 3631
rect 290 3618 342 3621
rect 346 3618 374 3621
rect 646 3621 649 3628
rect 2342 3622 2345 3628
rect 578 3618 649 3621
rect 746 3618 966 3621
rect 1234 3618 1318 3621
rect 2010 3618 2246 3621
rect 2390 3618 2398 3621
rect 2402 3618 2510 3621
rect 2514 3618 2550 3621
rect 2970 3618 3006 3621
rect 3010 3618 3158 3621
rect 3282 3618 3302 3621
rect 3442 3618 3598 3621
rect 3626 3618 3638 3621
rect 3642 3618 3758 3621
rect 4074 3618 4078 3621
rect 4738 3618 4886 3621
rect 4890 3618 5006 3621
rect 5010 3618 5070 3621
rect 5226 3618 5262 3621
rect 226 3608 334 3611
rect 778 3608 830 3611
rect 1274 3608 1278 3611
rect 1282 3608 1334 3611
rect 1338 3608 1358 3611
rect 2522 3608 2670 3611
rect 2682 3608 2862 3611
rect 2994 3608 3398 3611
rect 344 3603 346 3607
rect 350 3603 353 3607
rect 358 3603 360 3607
rect 1368 3603 1370 3607
rect 1374 3603 1377 3607
rect 1382 3603 1384 3607
rect 2392 3603 2394 3607
rect 2398 3603 2401 3607
rect 2406 3603 2408 3607
rect 3416 3603 3418 3607
rect 3422 3603 3425 3607
rect 3430 3603 3432 3607
rect 4440 3603 4442 3607
rect 4446 3603 4449 3607
rect 4454 3603 4456 3607
rect 818 3598 902 3601
rect 1242 3598 1358 3601
rect 1658 3598 1686 3601
rect 2138 3598 2270 3601
rect 2666 3598 2774 3601
rect 2778 3598 2798 3601
rect 326 3588 334 3591
rect 338 3588 542 3591
rect 650 3588 774 3591
rect 830 3588 838 3591
rect 842 3588 878 3591
rect 1194 3588 1446 3591
rect 1450 3588 1510 3591
rect 1650 3588 1742 3591
rect 2162 3588 2238 3591
rect 2242 3588 2302 3591
rect 2562 3588 3022 3591
rect 4394 3588 4438 3591
rect 554 3578 854 3581
rect 1322 3578 1694 3581
rect 2130 3578 2278 3581
rect 2290 3578 2422 3581
rect 2426 3578 2686 3581
rect 2730 3578 3126 3581
rect 4046 3581 4049 3588
rect 4046 3578 4102 3581
rect 4134 3581 4137 3588
rect 4134 3578 4182 3581
rect 4378 3578 4446 3581
rect 4522 3578 4558 3581
rect 4562 3578 4694 3581
rect 178 3568 246 3571
rect 698 3568 742 3571
rect 1306 3568 1326 3571
rect 1346 3568 1374 3571
rect 1378 3568 1414 3571
rect 1518 3568 1526 3571
rect 1530 3568 1550 3571
rect 1578 3568 1622 3571
rect 1626 3568 1686 3571
rect 1810 3568 1902 3571
rect 1906 3568 1934 3571
rect 2178 3568 2209 3571
rect 2370 3568 2534 3571
rect 2594 3568 2622 3571
rect 2658 3568 2662 3571
rect 2746 3568 2950 3571
rect 3194 3568 3198 3571
rect 3810 3568 3910 3571
rect 3914 3568 4310 3571
rect 4338 3568 4350 3571
rect 4354 3568 4374 3571
rect 4466 3568 4518 3571
rect 4522 3568 4590 3571
rect 5066 3568 5214 3571
rect 5306 3568 5358 3571
rect 14 3561 17 3568
rect 14 3558 86 3561
rect 178 3558 214 3561
rect 266 3558 294 3561
rect 298 3558 430 3561
rect 434 3558 446 3561
rect 562 3558 630 3561
rect 650 3558 686 3561
rect 690 3558 742 3561
rect 762 3558 822 3561
rect 826 3558 846 3561
rect 874 3558 918 3561
rect 922 3558 982 3561
rect 1070 3561 1073 3568
rect 986 3558 1073 3561
rect 1098 3558 1126 3561
rect 1130 3558 1137 3561
rect 1146 3558 1150 3561
rect 1282 3558 1326 3561
rect 1330 3558 1342 3561
rect 1506 3558 1662 3561
rect 1750 3561 1753 3568
rect 2206 3562 2209 3568
rect 1730 3558 1753 3561
rect 1770 3558 1894 3561
rect 1898 3558 1958 3561
rect 1962 3558 2014 3561
rect 2150 3558 2182 3561
rect 2210 3558 2246 3561
rect 2282 3558 2318 3561
rect 2418 3558 2446 3561
rect 2494 3558 2510 3561
rect 2550 3561 2553 3568
rect 2550 3558 2606 3561
rect 2610 3558 2630 3561
rect 2674 3558 2782 3561
rect 2966 3558 3038 3561
rect 3042 3558 3062 3561
rect 3122 3558 3198 3561
rect 3202 3558 3350 3561
rect 3354 3558 3638 3561
rect 3890 3558 3982 3561
rect 4178 3558 4222 3561
rect 4314 3558 4342 3561
rect 4410 3558 4470 3561
rect 4530 3558 4582 3561
rect 4586 3558 4614 3561
rect 4674 3558 4702 3561
rect 4722 3558 4734 3561
rect 4766 3561 4769 3568
rect 4766 3558 4846 3561
rect 4850 3558 5022 3561
rect 5298 3558 5310 3561
rect 122 3548 134 3551
rect 202 3548 214 3551
rect 426 3548 438 3551
rect 722 3548 750 3551
rect 906 3548 950 3551
rect 970 3548 998 3551
rect 1002 3548 1041 3551
rect 1098 3548 1118 3551
rect 1122 3548 1166 3551
rect 1298 3548 1318 3551
rect 1362 3548 1382 3551
rect 1406 3551 1409 3558
rect 2150 3552 2153 3558
rect 1386 3548 1409 3551
rect 1474 3548 1478 3551
rect 1482 3548 1486 3551
rect 1554 3548 1574 3551
rect 1578 3548 1598 3551
rect 1618 3548 1718 3551
rect 1722 3548 1785 3551
rect 1794 3548 1846 3551
rect 1858 3548 1862 3551
rect 1914 3548 1926 3551
rect 1930 3548 1950 3551
rect 1954 3548 2030 3551
rect 2194 3548 2230 3551
rect 2266 3548 2334 3551
rect 2338 3548 2358 3551
rect 2362 3548 2398 3551
rect 2402 3548 2438 3551
rect 2446 3551 2449 3558
rect 2494 3552 2497 3558
rect 2966 3552 2969 3558
rect 2446 3548 2486 3551
rect 2586 3548 2670 3551
rect 2722 3548 2822 3551
rect 2826 3548 2854 3551
rect 3330 3548 3446 3551
rect 3626 3548 3630 3551
rect 3650 3548 3822 3551
rect 3846 3548 3886 3551
rect 4094 3551 4097 3558
rect 3906 3548 4110 3551
rect 4170 3548 4214 3551
rect 4218 3548 4238 3551
rect 4242 3548 4350 3551
rect 4386 3548 4398 3551
rect 4490 3548 4494 3551
rect 4498 3548 4630 3551
rect 4642 3548 4662 3551
rect 4786 3548 4806 3551
rect 4890 3548 4918 3551
rect 4994 3548 5078 3551
rect 5082 3548 5086 3551
rect 5158 3551 5161 3558
rect 5130 3548 5161 3551
rect 5194 3548 5246 3551
rect 5282 3548 5286 3551
rect 58 3538 126 3541
rect 454 3541 457 3548
rect 1038 3542 1041 3548
rect 402 3538 457 3541
rect 474 3538 534 3541
rect 562 3538 798 3541
rect 1058 3538 1086 3541
rect 1090 3538 1094 3541
rect 1186 3538 1190 3541
rect 1354 3538 1398 3541
rect 1402 3538 1430 3541
rect 1434 3538 1582 3541
rect 1586 3538 1590 3541
rect 1714 3538 1758 3541
rect 1782 3541 1785 3548
rect 1782 3538 1814 3541
rect 1842 3538 1862 3541
rect 1866 3538 2046 3541
rect 2070 3541 2073 3548
rect 2070 3538 2542 3541
rect 2546 3538 2558 3541
rect 2562 3538 2638 3541
rect 2682 3538 2830 3541
rect 2850 3538 2918 3541
rect 3014 3541 3017 3548
rect 3014 3538 3046 3541
rect 3082 3538 3118 3541
rect 3122 3538 3137 3541
rect 82 3528 86 3531
rect 90 3528 118 3531
rect 122 3528 166 3531
rect 234 3528 262 3531
rect 266 3528 278 3531
rect 306 3528 318 3531
rect 442 3528 478 3531
rect 542 3531 545 3538
rect 542 3528 566 3531
rect 626 3528 646 3531
rect 650 3528 718 3531
rect 914 3528 934 3531
rect 938 3528 942 3531
rect 946 3528 1062 3531
rect 1066 3528 1118 3531
rect 1170 3528 1190 3531
rect 1430 3531 1433 3538
rect 3134 3532 3137 3538
rect 3454 3541 3457 3548
rect 3846 3542 3849 3548
rect 3426 3538 3457 3541
rect 3582 3538 3710 3541
rect 3738 3538 3758 3541
rect 3930 3538 4062 3541
rect 4090 3538 4126 3541
rect 4154 3538 4190 3541
rect 4330 3538 4358 3541
rect 4362 3538 4374 3541
rect 4378 3538 4430 3541
rect 4434 3538 4510 3541
rect 4546 3538 4566 3541
rect 4610 3538 4646 3541
rect 4674 3538 4702 3541
rect 4826 3538 4862 3541
rect 4866 3538 4942 3541
rect 1430 3528 1454 3531
rect 1478 3528 1534 3531
rect 1570 3528 1606 3531
rect 1746 3528 1814 3531
rect 1818 3528 1822 3531
rect 1826 3528 1862 3531
rect 1922 3528 1942 3531
rect 1946 3528 2006 3531
rect 2162 3528 2190 3531
rect 2238 3528 2270 3531
rect 2298 3528 2302 3531
rect 2346 3528 2350 3531
rect 2402 3528 2422 3531
rect 2426 3528 2454 3531
rect 2538 3528 2590 3531
rect 2634 3528 2654 3531
rect 2698 3528 2766 3531
rect 2826 3528 2958 3531
rect 2962 3528 2990 3531
rect 2994 3528 3006 3531
rect 3142 3531 3145 3538
rect 3582 3532 3585 3538
rect 4302 3532 4305 3538
rect 3142 3528 3182 3531
rect 3618 3528 3662 3531
rect 3670 3528 3726 3531
rect 4566 3531 4569 3538
rect 4450 3528 4662 3531
rect 4682 3528 4710 3531
rect 4842 3528 4886 3531
rect 4890 3528 4894 3531
rect 4922 3528 4926 3531
rect 4930 3528 4982 3531
rect 5210 3528 5262 3531
rect 1478 3522 1481 3528
rect 2238 3522 2241 3528
rect 3670 3522 3673 3528
rect 154 3518 230 3521
rect 250 3518 286 3521
rect 346 3518 390 3521
rect 394 3518 494 3521
rect 506 3518 1318 3521
rect 1762 3518 1966 3521
rect 2146 3518 2166 3521
rect 2242 3518 2310 3521
rect 2514 3518 2598 3521
rect 2666 3518 2734 3521
rect 2738 3518 2750 3521
rect 2890 3518 3094 3521
rect 3570 3518 3630 3521
rect 3682 3518 3718 3521
rect 3890 3518 4742 3521
rect 4746 3518 4750 3521
rect 4858 3518 4950 3521
rect 882 3508 926 3511
rect 930 3508 950 3511
rect 954 3508 1014 3511
rect 1298 3508 1414 3511
rect 1418 3508 1510 3511
rect 1666 3508 1766 3511
rect 2122 3508 2158 3511
rect 2218 3508 2414 3511
rect 2426 3508 2494 3511
rect 2498 3508 2526 3511
rect 2730 3508 2742 3511
rect 2818 3508 2894 3511
rect 3178 3508 3502 3511
rect 3506 3508 3670 3511
rect 3698 3508 3814 3511
rect 3818 3508 3870 3511
rect 3874 3508 3902 3511
rect 4122 3508 4718 3511
rect 856 3503 858 3507
rect 862 3503 865 3507
rect 870 3503 872 3507
rect 1872 3503 1874 3507
rect 1878 3503 1881 3507
rect 1886 3503 1888 3507
rect 2904 3503 2906 3507
rect 2910 3503 2913 3507
rect 2918 3503 2920 3507
rect 3928 3503 3930 3507
rect 3934 3503 3937 3507
rect 3942 3503 3944 3507
rect 4952 3503 4954 3507
rect 4958 3503 4961 3507
rect 4966 3503 4968 3507
rect 202 3498 246 3501
rect 250 3498 294 3501
rect 418 3498 422 3501
rect 426 3498 526 3501
rect 594 3498 782 3501
rect 1010 3498 1158 3501
rect 1162 3498 1302 3501
rect 1654 3498 1790 3501
rect 1794 3498 1830 3501
rect 1994 3498 2046 3501
rect 2066 3498 2350 3501
rect 2354 3498 2470 3501
rect 2474 3498 2622 3501
rect 2770 3498 2878 3501
rect 3114 3498 3190 3501
rect 3346 3498 3478 3501
rect 3482 3498 3534 3501
rect 3610 3498 3702 3501
rect 4498 3498 4550 3501
rect 4770 3498 4830 3501
rect 4834 3498 4854 3501
rect 582 3488 614 3491
rect 826 3488 929 3491
rect 1154 3488 1174 3491
rect 1178 3488 1222 3491
rect 1654 3491 1657 3498
rect 1282 3488 1657 3491
rect 1690 3488 1838 3491
rect 1858 3488 1966 3491
rect 1970 3488 2022 3491
rect 2202 3488 2214 3491
rect 2258 3488 2574 3491
rect 2578 3488 2646 3491
rect 2706 3488 2910 3491
rect 2954 3488 2966 3491
rect 2994 3488 3086 3491
rect 3114 3488 3126 3491
rect 3362 3488 3366 3491
rect 4194 3488 4278 3491
rect 4474 3488 4486 3491
rect 4530 3488 4542 3491
rect 4802 3488 4902 3491
rect 5002 3488 5094 3491
rect 582 3482 585 3488
rect 926 3482 929 3488
rect 98 3478 110 3481
rect 114 3478 126 3481
rect 274 3478 446 3481
rect 458 3478 542 3481
rect 546 3478 574 3481
rect 610 3478 630 3481
rect 634 3478 654 3481
rect 658 3478 678 3481
rect 842 3478 918 3481
rect 1402 3478 1446 3481
rect 1490 3478 1513 3481
rect 1522 3478 1622 3481
rect 102 3468 182 3471
rect 186 3468 302 3471
rect 330 3468 390 3471
rect 450 3468 518 3471
rect 554 3468 558 3471
rect 562 3468 590 3471
rect 642 3468 686 3471
rect 842 3468 902 3471
rect 1034 3468 1054 3471
rect 1126 3471 1129 3478
rect 1058 3468 1129 3471
rect 1330 3468 1406 3471
rect 1410 3468 1494 3471
rect 1510 3471 1513 3478
rect 1510 3468 1582 3471
rect 1662 3471 1665 3488
rect 1674 3478 1678 3481
rect 1714 3478 1782 3481
rect 1850 3478 1862 3481
rect 2146 3478 2198 3481
rect 2314 3478 2326 3481
rect 2362 3478 2465 3481
rect 2618 3478 2726 3481
rect 2906 3478 2958 3481
rect 3158 3481 3161 3488
rect 2962 3478 3161 3481
rect 3274 3478 3358 3481
rect 3466 3478 3638 3481
rect 3686 3481 3689 3488
rect 3642 3478 3689 3481
rect 3722 3478 3782 3481
rect 3922 3478 4062 3481
rect 4066 3478 4086 3481
rect 4142 3481 4145 3488
rect 4090 3478 4145 3481
rect 4358 3481 4361 3488
rect 4178 3478 4361 3481
rect 4406 3481 4409 3488
rect 4422 3481 4425 3488
rect 4406 3478 4425 3481
rect 4474 3478 4478 3481
rect 4494 3481 4497 3488
rect 4494 3478 4518 3481
rect 4774 3481 4777 3488
rect 4650 3478 4777 3481
rect 4850 3478 4878 3481
rect 5010 3478 5014 3481
rect 5066 3478 5206 3481
rect 1602 3468 1665 3471
rect 1686 3471 1689 3478
rect 1674 3468 1689 3471
rect 1698 3468 1734 3471
rect 1902 3471 1905 3478
rect 2222 3472 2225 3478
rect 2462 3472 2465 3478
rect 1874 3468 1905 3471
rect 1962 3468 1966 3471
rect 2114 3468 2134 3471
rect 2138 3468 2190 3471
rect 2306 3468 2310 3471
rect 2330 3468 2398 3471
rect 2402 3468 2457 3471
rect 2698 3468 2726 3471
rect 2870 3471 2873 3478
rect 2870 3468 2969 3471
rect 2978 3468 2982 3471
rect 3082 3468 3166 3471
rect 3450 3468 3638 3471
rect 3838 3471 3841 3478
rect 4574 3472 4577 3478
rect 3642 3468 3841 3471
rect 3954 3468 4038 3471
rect 4042 3468 4110 3471
rect 4130 3468 4182 3471
rect 4186 3468 4206 3471
rect 4274 3468 4302 3471
rect 4346 3468 4390 3471
rect 4410 3468 4486 3471
rect 4610 3468 4614 3471
rect 4762 3468 4854 3471
rect 4890 3468 4926 3471
rect 5010 3468 5022 3471
rect 5266 3468 5294 3471
rect 102 3462 105 3468
rect 34 3458 62 3461
rect 154 3458 198 3461
rect 258 3458 262 3461
rect 266 3458 286 3461
rect 310 3461 313 3468
rect 750 3462 753 3468
rect 1198 3462 1201 3468
rect 310 3458 358 3461
rect 362 3458 406 3461
rect 450 3458 454 3461
rect 498 3458 534 3461
rect 570 3458 630 3461
rect 634 3458 670 3461
rect 802 3458 854 3461
rect 1006 3458 1014 3461
rect 1018 3458 1062 3461
rect 1066 3458 1094 3461
rect 1122 3458 1134 3461
rect 1138 3458 1174 3461
rect 1346 3458 1590 3461
rect 1658 3458 1678 3461
rect 1714 3458 1726 3461
rect 1858 3458 1894 3461
rect 2090 3458 2102 3461
rect 2286 3461 2289 3468
rect 2218 3458 2289 3461
rect 2298 3458 2406 3461
rect 2454 3461 2457 3468
rect 2454 3458 2470 3461
rect 2586 3458 2614 3461
rect 2694 3461 2697 3468
rect 2966 3462 2969 3468
rect 2642 3458 2697 3461
rect 2922 3458 2958 3461
rect 2986 3458 2990 3461
rect 3002 3458 3038 3461
rect 3254 3458 3398 3461
rect 3634 3458 3686 3461
rect 3866 3458 4094 3461
rect 4186 3458 4198 3461
rect 4210 3458 4222 3461
rect 4230 3461 4233 3468
rect 4494 3462 4497 3468
rect 4230 3458 4294 3461
rect 4330 3458 4366 3461
rect 4394 3458 4462 3461
rect 4634 3458 4670 3461
rect 4890 3458 4894 3461
rect 4938 3458 4998 3461
rect 5002 3458 5017 3461
rect 5114 3458 5145 3461
rect 118 3451 121 3458
rect 98 3448 121 3451
rect 238 3451 241 3458
rect 138 3448 318 3451
rect 594 3448 614 3451
rect 814 3448 830 3451
rect 942 3451 945 3458
rect 914 3448 945 3451
rect 1042 3448 1065 3451
rect 1330 3448 1350 3451
rect 1422 3448 1430 3451
rect 1434 3448 1606 3451
rect 1750 3451 1753 3458
rect 1682 3448 1753 3451
rect 1786 3448 1814 3451
rect 1818 3448 1942 3451
rect 2114 3448 2126 3451
rect 2226 3448 2230 3451
rect 2258 3448 2278 3451
rect 2294 3451 2297 3458
rect 2294 3448 2318 3451
rect 2354 3448 2382 3451
rect 2386 3448 2494 3451
rect 2546 3448 2750 3451
rect 2898 3448 2926 3451
rect 3018 3448 3118 3451
rect 3142 3451 3145 3458
rect 3130 3448 3145 3451
rect 3254 3452 3257 3458
rect 5014 3452 5017 3458
rect 5142 3452 5145 3458
rect 5270 3452 5273 3458
rect 3578 3448 3590 3451
rect 3706 3448 3710 3451
rect 3714 3448 3950 3451
rect 4194 3448 4254 3451
rect 4286 3448 4294 3451
rect 4298 3448 4334 3451
rect 4366 3448 4374 3451
rect 4378 3448 4622 3451
rect 4786 3448 4798 3451
rect 4818 3448 4830 3451
rect 4878 3448 4886 3451
rect 814 3442 817 3448
rect 1062 3442 1065 3448
rect 226 3438 294 3441
rect 514 3438 526 3441
rect 1370 3438 1390 3441
rect 1438 3438 1446 3441
rect 1450 3438 1534 3441
rect 1554 3438 1702 3441
rect 1714 3438 1718 3441
rect 2134 3441 2137 3448
rect 2134 3438 2334 3441
rect 2522 3438 2558 3441
rect 2794 3438 2830 3441
rect 3058 3438 3150 3441
rect 3778 3438 3782 3441
rect 4154 3438 4214 3441
rect 4250 3438 4270 3441
rect 4342 3441 4345 3448
rect 4878 3442 4881 3448
rect 4274 3438 4398 3441
rect 4466 3438 4478 3441
rect 4722 3438 4726 3441
rect 5266 3438 5270 3441
rect 5278 3432 5281 3438
rect 378 3428 526 3431
rect 650 3428 958 3431
rect 1386 3428 1462 3431
rect 1490 3428 1558 3431
rect 2210 3428 2686 3431
rect 2690 3428 2718 3431
rect 2850 3428 3030 3431
rect 3050 3428 3062 3431
rect 3106 3428 3158 3431
rect 3162 3428 3286 3431
rect 3802 3428 3846 3431
rect 4394 3428 5030 3431
rect 482 3418 494 3421
rect 498 3418 582 3421
rect 762 3418 846 3421
rect 850 3418 950 3421
rect 954 3418 974 3421
rect 1306 3418 1430 3421
rect 1486 3421 1489 3428
rect 1458 3418 1489 3421
rect 2318 3418 2326 3421
rect 2330 3418 2486 3421
rect 2726 3412 2729 3428
rect 3134 3422 3137 3428
rect 4098 3418 4726 3421
rect 4730 3418 4750 3421
rect 402 3408 422 3411
rect 634 3408 670 3411
rect 674 3408 766 3411
rect 1394 3408 1462 3411
rect 2514 3408 2630 3411
rect 3186 3408 3318 3411
rect 3538 3408 3542 3411
rect 4594 3408 4798 3411
rect 344 3403 346 3407
rect 350 3403 353 3407
rect 358 3403 360 3407
rect 1368 3403 1370 3407
rect 1374 3403 1377 3407
rect 1382 3403 1384 3407
rect 2392 3403 2394 3407
rect 2398 3403 2401 3407
rect 2406 3403 2408 3407
rect 3416 3403 3418 3407
rect 3422 3403 3425 3407
rect 3430 3403 3432 3407
rect 4440 3403 4442 3407
rect 4446 3403 4449 3407
rect 4454 3403 4456 3407
rect 666 3398 686 3401
rect 1146 3398 1302 3401
rect 1498 3398 1598 3401
rect 2018 3398 2030 3401
rect 2482 3398 2622 3401
rect 2626 3398 2726 3401
rect 2962 3398 3342 3401
rect 3730 3398 3766 3401
rect 3954 3398 4238 3401
rect 4650 3398 4654 3401
rect 2094 3392 2097 3398
rect 58 3388 62 3391
rect 122 3388 126 3391
rect 130 3388 286 3391
rect 610 3388 686 3391
rect 1322 3388 1446 3391
rect 1450 3388 1486 3391
rect 2530 3388 2678 3391
rect 2986 3388 3206 3391
rect 3338 3388 3566 3391
rect 3954 3388 4118 3391
rect 5018 3388 5238 3391
rect 274 3378 310 3381
rect 314 3378 398 3381
rect 446 3381 449 3388
rect 410 3378 449 3381
rect 490 3378 494 3381
rect 538 3378 566 3381
rect 1182 3381 1185 3388
rect 1146 3378 1185 3381
rect 1518 3381 1521 3388
rect 1338 3378 1521 3381
rect 1666 3378 1782 3381
rect 1962 3378 2206 3381
rect 2318 3381 2321 3388
rect 2282 3378 2321 3381
rect 2538 3378 2585 3381
rect 2594 3378 2598 3381
rect 2658 3378 2662 3381
rect 2770 3378 3046 3381
rect 3066 3378 3214 3381
rect 3218 3378 3270 3381
rect 4018 3378 4174 3381
rect 4698 3378 5110 3381
rect 146 3368 158 3371
rect 194 3368 358 3371
rect 386 3368 414 3371
rect 466 3368 478 3371
rect 530 3368 534 3371
rect 554 3368 574 3371
rect 630 3371 633 3378
rect 2582 3372 2585 3378
rect 594 3368 633 3371
rect 706 3368 710 3371
rect 722 3368 782 3371
rect 802 3368 814 3371
rect 1010 3368 1062 3371
rect 1098 3368 1110 3371
rect 1170 3368 1182 3371
rect 1194 3368 1718 3371
rect 1738 3368 1838 3371
rect 2010 3368 2070 3371
rect 2146 3368 2150 3371
rect 2338 3368 2350 3371
rect 2386 3368 2574 3371
rect 2586 3368 2718 3371
rect 2722 3368 2742 3371
rect 2850 3368 2862 3371
rect 3034 3368 3198 3371
rect 3546 3368 3630 3371
rect 3890 3368 3958 3371
rect 4082 3368 4086 3371
rect 4090 3368 4110 3371
rect 4818 3368 4841 3371
rect 4858 3368 4910 3371
rect 4986 3368 5078 3371
rect 5082 3368 5102 3371
rect 5130 3368 5142 3371
rect 5258 3368 5270 3371
rect 54 3361 57 3368
rect 54 3358 78 3361
rect 282 3358 846 3361
rect 954 3358 1022 3361
rect 1030 3358 1038 3361
rect 1042 3358 1070 3361
rect 1082 3358 1214 3361
rect 1458 3358 1534 3361
rect 1570 3358 1574 3361
rect 1578 3358 1585 3361
rect 1778 3358 1822 3361
rect 1866 3358 1902 3361
rect 2074 3358 2150 3361
rect 2322 3358 2342 3361
rect 2362 3358 2486 3361
rect 2490 3358 2606 3361
rect 2626 3358 2638 3361
rect 2694 3358 2702 3361
rect 2706 3358 2758 3361
rect 2818 3358 2862 3361
rect 2866 3358 2886 3361
rect 2898 3358 2950 3361
rect 2954 3358 2990 3361
rect 3178 3358 3198 3361
rect 3234 3358 3246 3361
rect 3850 3358 3854 3361
rect 4058 3358 4089 3361
rect 4106 3358 4110 3361
rect 4238 3361 4241 3368
rect 4838 3362 4841 3368
rect 4238 3358 4438 3361
rect 4682 3358 4686 3361
rect 4906 3358 4982 3361
rect 5002 3358 5006 3361
rect 5282 3358 5286 3361
rect 5290 3358 5302 3361
rect 1254 3352 1257 3358
rect 18 3348 62 3351
rect 66 3348 150 3351
rect 250 3348 630 3351
rect 634 3348 654 3351
rect 658 3348 1198 3351
rect 1274 3348 1278 3351
rect 1422 3351 1425 3358
rect 1422 3348 1462 3351
rect 1498 3348 1550 3351
rect 1554 3348 1622 3351
rect 1714 3348 1718 3351
rect 1802 3348 1894 3351
rect 2058 3348 2062 3351
rect 2074 3348 2094 3351
rect 2146 3348 2166 3351
rect 2306 3348 2414 3351
rect 2466 3348 2526 3351
rect 2578 3348 2598 3351
rect 2658 3348 2702 3351
rect 2834 3348 2838 3351
rect 3050 3348 3078 3351
rect 3186 3348 3190 3351
rect 3722 3348 3766 3351
rect 3814 3351 3817 3358
rect 4086 3352 4089 3358
rect 3770 3348 3854 3351
rect 3930 3348 4022 3351
rect 4354 3348 4390 3351
rect 4546 3348 4598 3351
rect 4890 3348 4926 3351
rect 4990 3351 4993 3358
rect 5022 3352 5025 3358
rect 5182 3352 5185 3358
rect 4930 3348 4993 3351
rect 5010 3348 5014 3351
rect 5098 3348 5102 3351
rect 98 3338 158 3341
rect 162 3338 230 3341
rect 262 3338 302 3341
rect 394 3338 406 3341
rect 410 3338 414 3341
rect 458 3338 550 3341
rect 578 3338 598 3341
rect 610 3338 630 3341
rect 690 3338 694 3341
rect 706 3340 734 3341
rect 706 3338 737 3340
rect 762 3338 774 3341
rect 786 3338 878 3341
rect 1010 3338 1030 3341
rect 1050 3338 1110 3341
rect 1246 3341 1249 3348
rect 1218 3338 1249 3341
rect 1354 3338 1358 3341
rect 1370 3338 1374 3341
rect 1478 3341 1481 3348
rect 1434 3338 1481 3341
rect 1546 3338 1558 3341
rect 1562 3338 1630 3341
rect 1738 3338 1742 3341
rect 1770 3338 1774 3341
rect 1818 3338 1862 3341
rect 2054 3338 2078 3341
rect 2114 3338 2158 3341
rect 2162 3338 2190 3341
rect 2298 3338 2390 3341
rect 2430 3341 2433 3348
rect 4278 3342 4281 3348
rect 4734 3342 4737 3348
rect 2430 3338 2502 3341
rect 2522 3338 2550 3341
rect 2570 3338 2646 3341
rect 2690 3338 2721 3341
rect 2730 3338 2774 3341
rect 2778 3338 2838 3341
rect 2890 3338 2894 3341
rect 2978 3338 2982 3341
rect 3098 3338 3126 3341
rect 3266 3338 3302 3341
rect 3442 3338 3478 3341
rect 3842 3338 3902 3341
rect 4358 3338 4462 3341
rect 4466 3338 4486 3341
rect 4546 3338 4614 3341
rect 4618 3338 4646 3341
rect 4794 3338 4878 3341
rect 4882 3338 4886 3341
rect 4906 3338 4910 3341
rect 4914 3338 4934 3341
rect 4966 3338 5006 3341
rect 5050 3338 5086 3341
rect 5106 3338 5134 3341
rect 5218 3338 5246 3341
rect 54 3331 57 3338
rect 262 3332 265 3338
rect 646 3332 649 3338
rect 966 3332 969 3338
rect 54 3328 126 3331
rect 298 3328 310 3331
rect 434 3328 481 3331
rect 490 3328 494 3331
rect 710 3328 718 3331
rect 722 3328 798 3331
rect 818 3328 918 3331
rect 994 3328 1110 3331
rect 1114 3328 1166 3331
rect 1198 3331 1201 3338
rect 1702 3332 1705 3338
rect 2054 3332 2057 3338
rect 1170 3328 1201 3331
rect 1242 3328 1262 3331
rect 1274 3328 1454 3331
rect 1474 3328 1510 3331
rect 1514 3328 1518 3331
rect 1610 3328 1670 3331
rect 1714 3328 1814 3331
rect 1818 3328 1838 3331
rect 2130 3328 2174 3331
rect 2186 3328 2302 3331
rect 2322 3328 2358 3331
rect 2482 3328 2486 3331
rect 2506 3328 2590 3331
rect 2594 3328 2606 3331
rect 2650 3328 2678 3331
rect 2718 3331 2721 3338
rect 2718 3328 2782 3331
rect 3006 3331 3009 3338
rect 2834 3328 3009 3331
rect 3066 3328 3110 3331
rect 3130 3328 3166 3331
rect 3190 3331 3193 3338
rect 4358 3332 4361 3338
rect 4966 3332 4969 3338
rect 3190 3328 3222 3331
rect 3434 3328 3454 3331
rect 3658 3328 3798 3331
rect 3802 3328 3894 3331
rect 3922 3328 3974 3331
rect 4038 3328 4078 3331
rect 4106 3328 4326 3331
rect 4442 3328 4614 3331
rect 4634 3328 4670 3331
rect 4842 3328 4870 3331
rect 5150 3328 5190 3331
rect 294 3321 297 3328
rect 478 3322 481 3328
rect 1734 3322 1737 3328
rect 2094 3322 2097 3328
rect 4038 3322 4041 3328
rect 4246 3322 4249 3328
rect 5150 3322 5153 3328
rect 266 3318 297 3321
rect 410 3318 462 3321
rect 490 3318 510 3321
rect 650 3318 1014 3321
rect 1018 3318 1046 3321
rect 1074 3318 1094 3321
rect 1106 3318 1182 3321
rect 1194 3318 1230 3321
rect 1330 3318 1406 3321
rect 1426 3318 1470 3321
rect 1474 3318 1534 3321
rect 1538 3318 1654 3321
rect 1862 3318 2006 3321
rect 2266 3318 2318 3321
rect 2778 3318 2966 3321
rect 2970 3318 3014 3321
rect 3450 3318 3510 3321
rect 3786 3318 3926 3321
rect 4554 3318 4558 3321
rect 4610 3318 4710 3321
rect 4826 3318 4854 3321
rect 210 3308 278 3311
rect 618 3308 622 3311
rect 962 3308 974 3311
rect 1050 3308 1134 3311
rect 1138 3308 1158 3311
rect 1862 3311 1865 3318
rect 1690 3308 1865 3311
rect 2314 3308 2358 3311
rect 3370 3308 3718 3311
rect 3722 3308 3742 3311
rect 3770 3308 3918 3311
rect 4002 3308 4030 3311
rect 4042 3308 4094 3311
rect 4394 3308 4502 3311
rect 4506 3308 4534 3311
rect 4586 3308 4606 3311
rect 4802 3308 4894 3311
rect 856 3303 858 3307
rect 862 3303 865 3307
rect 870 3303 872 3307
rect 942 3302 945 3308
rect 170 3298 222 3301
rect 234 3298 358 3301
rect 362 3298 382 3301
rect 426 3298 486 3301
rect 574 3298 782 3301
rect 906 3298 910 3301
rect 950 3301 953 3308
rect 1872 3303 1874 3307
rect 1878 3303 1881 3307
rect 1886 3303 1888 3307
rect 2038 3302 2041 3308
rect 2904 3303 2906 3307
rect 2910 3303 2913 3307
rect 2918 3303 2920 3307
rect 3928 3303 3930 3307
rect 3934 3303 3937 3307
rect 3942 3303 3944 3307
rect 4952 3303 4954 3307
rect 4958 3303 4961 3307
rect 4966 3303 4968 3307
rect 950 3298 966 3301
rect 986 3298 990 3301
rect 1138 3298 1190 3301
rect 1354 3298 1710 3301
rect 1714 3298 1830 3301
rect 2242 3298 2358 3301
rect 3090 3298 3094 3301
rect 3354 3298 3358 3301
rect 3426 3298 3542 3301
rect 3610 3298 3822 3301
rect 4234 3298 4414 3301
rect 4474 3298 4494 3301
rect 4730 3298 4774 3301
rect 4818 3298 4838 3301
rect 4874 3298 4905 3301
rect 574 3292 577 3298
rect 3846 3292 3849 3298
rect 4902 3292 4905 3298
rect 54 3288 126 3291
rect 130 3288 254 3291
rect 330 3288 574 3291
rect 714 3288 718 3291
rect 722 3288 750 3291
rect 798 3288 806 3291
rect 822 3288 830 3291
rect 834 3288 1006 3291
rect 1034 3288 1062 3291
rect 1082 3288 1249 3291
rect 1258 3288 1262 3291
rect 1290 3288 1390 3291
rect 1454 3288 1926 3291
rect 1930 3288 1990 3291
rect 1994 3288 2014 3291
rect 2018 3288 2022 3291
rect 2034 3288 2182 3291
rect 2190 3288 2198 3291
rect 2202 3288 2222 3291
rect 2230 3288 2238 3291
rect 2242 3288 2270 3291
rect 2274 3288 2302 3291
rect 2874 3288 2974 3291
rect 3026 3288 3038 3291
rect 3074 3288 3102 3291
rect 3106 3288 3158 3291
rect 3298 3288 3310 3291
rect 3330 3288 3550 3291
rect 4058 3288 4126 3291
rect 4362 3288 4550 3291
rect 4666 3288 4670 3291
rect 4866 3288 4870 3291
rect 4906 3288 4934 3291
rect 5250 3288 5262 3291
rect 54 3282 57 3288
rect 798 3282 801 3288
rect 1246 3282 1249 3288
rect 1454 3282 1457 3288
rect 74 3278 86 3281
rect 90 3278 102 3281
rect 114 3278 137 3281
rect 146 3278 206 3281
rect 394 3278 502 3281
rect 618 3278 670 3281
rect 810 3278 830 3281
rect 874 3278 910 3281
rect 962 3278 998 3281
rect 1018 3278 1118 3281
rect 1354 3278 1438 3281
rect 1650 3278 1678 3281
rect 1690 3278 1694 3281
rect 1746 3278 1838 3281
rect 1986 3278 2374 3281
rect 2378 3278 2446 3281
rect 2462 3281 2465 3288
rect 2726 3282 2729 3288
rect 2462 3278 2534 3281
rect 2626 3278 2686 3281
rect 3002 3278 3022 3281
rect 3062 3281 3065 3288
rect 3062 3278 3110 3281
rect 3114 3278 3206 3281
rect 3290 3278 3358 3281
rect 4218 3278 4382 3281
rect 4386 3278 4406 3281
rect 4490 3278 4513 3281
rect 4570 3278 4654 3281
rect 4690 3278 4694 3281
rect 4758 3281 4761 3288
rect 4950 3282 4953 3288
rect 4746 3278 4761 3281
rect 4858 3278 4886 3281
rect 4890 3278 4894 3281
rect 4922 3278 4942 3281
rect 4962 3278 4998 3281
rect 5026 3278 5062 3281
rect 5114 3278 5142 3281
rect 134 3272 137 3278
rect 58 3268 78 3271
rect 122 3268 126 3271
rect 138 3268 150 3271
rect 314 3268 326 3271
rect 562 3268 782 3271
rect 794 3268 1486 3271
rect 1490 3268 1542 3271
rect 1570 3268 1574 3271
rect 1674 3268 1678 3271
rect 1690 3268 2078 3271
rect 2082 3268 2118 3271
rect 2122 3268 2254 3271
rect 2258 3268 2558 3271
rect 2594 3268 2614 3271
rect 2634 3268 2670 3271
rect 2722 3268 2790 3271
rect 2794 3268 2814 3271
rect 2850 3268 2854 3271
rect 2898 3268 2934 3271
rect 2950 3271 2953 3278
rect 4510 3272 4513 3278
rect 2950 3268 2966 3271
rect 3026 3268 3070 3271
rect 3090 3268 3142 3271
rect 3146 3268 3294 3271
rect 3402 3268 3406 3271
rect 3466 3268 3494 3271
rect 3498 3268 3510 3271
rect 3514 3268 3566 3271
rect 4330 3268 4390 3271
rect 4722 3268 4734 3271
rect 4898 3268 4910 3271
rect 4914 3268 4918 3271
rect 4938 3268 4958 3271
rect 4962 3268 5046 3271
rect 5050 3268 5134 3271
rect 5206 3271 5209 3278
rect 5138 3268 5209 3271
rect 5342 3271 5346 3272
rect 5218 3268 5346 3271
rect 422 3262 425 3268
rect 18 3258 22 3261
rect 250 3258 262 3261
rect 338 3258 401 3261
rect 450 3258 470 3261
rect 554 3258 582 3261
rect 610 3258 726 3261
rect 730 3258 790 3261
rect 842 3258 878 3261
rect 914 3258 1022 3261
rect 1042 3258 1046 3261
rect 1074 3258 1102 3261
rect 1106 3258 1158 3261
rect 1278 3258 1318 3261
rect 1450 3258 1638 3261
rect 1698 3258 1718 3261
rect 1722 3258 1734 3261
rect 1774 3258 1782 3261
rect 1802 3258 1806 3261
rect 1838 3258 1886 3261
rect 2026 3258 2054 3261
rect 2066 3258 2110 3261
rect 2218 3258 2230 3261
rect 2282 3258 2329 3261
rect 2410 3258 2478 3261
rect 2482 3258 2510 3261
rect 2514 3258 2518 3261
rect 2570 3258 2646 3261
rect 2658 3258 2766 3261
rect 2770 3258 2918 3261
rect 2934 3261 2937 3268
rect 2934 3258 2998 3261
rect 3034 3258 3126 3261
rect 3258 3258 3286 3261
rect 3402 3258 3438 3261
rect 3574 3261 3577 3268
rect 4742 3262 4745 3268
rect 3506 3258 3545 3261
rect 3574 3258 3654 3261
rect 4154 3258 4169 3261
rect 42 3248 62 3251
rect 190 3251 193 3258
rect 106 3248 193 3251
rect 398 3252 401 3258
rect 902 3252 905 3258
rect 1278 3252 1281 3258
rect 1838 3252 1841 3258
rect 1966 3252 1969 3258
rect 566 3248 574 3251
rect 578 3248 673 3251
rect 682 3248 798 3251
rect 802 3248 814 3251
rect 986 3248 1190 3251
rect 1258 3248 1262 3251
rect 1298 3248 1390 3251
rect 1466 3248 1494 3251
rect 1514 3248 1558 3251
rect 1586 3248 1654 3251
rect 1722 3248 1774 3251
rect 1874 3248 1934 3251
rect 1986 3248 2001 3251
rect 2042 3248 2046 3251
rect 2106 3248 2142 3251
rect 2214 3251 2217 3258
rect 2326 3252 2329 3258
rect 2186 3248 2217 3251
rect 2282 3248 2286 3251
rect 2290 3248 2318 3251
rect 2434 3248 2494 3251
rect 2498 3248 2518 3251
rect 2714 3248 2742 3251
rect 2794 3248 2822 3251
rect 2938 3248 2958 3251
rect 3058 3248 3062 3251
rect 3066 3248 3166 3251
rect 3170 3248 3190 3251
rect 3198 3251 3201 3258
rect 3542 3252 3545 3258
rect 4110 3252 4113 3258
rect 4166 3252 4169 3258
rect 4474 3258 4550 3261
rect 4578 3258 4617 3261
rect 4634 3258 4670 3261
rect 4834 3258 4998 3261
rect 5002 3258 5081 3261
rect 5090 3258 5110 3261
rect 5170 3258 5214 3261
rect 5270 3258 5286 3261
rect 5290 3258 5294 3261
rect 4270 3252 4273 3258
rect 4614 3252 4617 3258
rect 3198 3248 3270 3251
rect 3478 3248 3497 3251
rect 3706 3248 3758 3251
rect 3986 3248 4038 3251
rect 4730 3248 4806 3251
rect 4810 3248 4982 3251
rect 5078 3251 5081 3258
rect 5270 3252 5273 3258
rect 5014 3248 5073 3251
rect 5078 3248 5198 3251
rect 5342 3248 5346 3252
rect 34 3238 94 3241
rect 178 3238 182 3241
rect 370 3238 478 3241
rect 482 3238 486 3241
rect 498 3238 502 3241
rect 506 3238 598 3241
rect 670 3241 673 3248
rect 1998 3242 2001 3248
rect 670 3238 686 3241
rect 858 3238 886 3241
rect 890 3238 926 3241
rect 970 3238 990 3241
rect 1010 3238 1142 3241
rect 1210 3238 1286 3241
rect 1290 3238 1526 3241
rect 1618 3238 1758 3241
rect 2086 3241 2089 3248
rect 2086 3238 2174 3241
rect 2350 3241 2353 3248
rect 3478 3242 3481 3248
rect 3494 3242 3497 3248
rect 5014 3242 5017 3248
rect 5070 3242 5073 3248
rect 2350 3238 2390 3241
rect 2554 3238 2838 3241
rect 3042 3238 3078 3241
rect 3090 3238 3094 3241
rect 3186 3238 3198 3241
rect 3218 3238 3246 3241
rect 3618 3238 3638 3241
rect 3714 3238 3718 3241
rect 4418 3238 4462 3241
rect 4474 3238 4734 3241
rect 5074 3238 5094 3241
rect 5198 3241 5201 3248
rect 5342 3241 5345 3248
rect 5198 3238 5345 3241
rect 274 3228 710 3231
rect 1202 3228 1294 3231
rect 1530 3228 1558 3231
rect 1562 3228 1566 3231
rect 2346 3228 2454 3231
rect 2618 3228 2678 3231
rect 2682 3228 2766 3231
rect 2906 3228 3430 3231
rect 3490 3228 3558 3231
rect 4402 3228 4558 3231
rect 5002 3228 5062 3231
rect 5066 3228 5118 3231
rect 5282 3228 5286 3231
rect 290 3218 350 3221
rect 354 3218 438 3221
rect 666 3218 734 3221
rect 1042 3218 1134 3221
rect 1138 3218 1150 3221
rect 1274 3218 1470 3221
rect 2154 3218 2478 3221
rect 2482 3218 2894 3221
rect 3158 3218 3166 3221
rect 3170 3218 3286 3221
rect 3290 3218 3382 3221
rect 4914 3218 5182 3221
rect 474 3208 534 3211
rect 2674 3208 2702 3211
rect 2722 3208 3102 3211
rect 3154 3208 3174 3211
rect 3178 3208 3222 3211
rect 3346 3208 3382 3211
rect 4202 3208 4214 3211
rect 4218 3208 4246 3211
rect 4250 3208 4334 3211
rect 344 3203 346 3207
rect 350 3203 353 3207
rect 358 3203 360 3207
rect 1368 3203 1370 3207
rect 1374 3203 1377 3207
rect 1382 3203 1384 3207
rect 2392 3203 2394 3207
rect 2398 3203 2401 3207
rect 2406 3203 2408 3207
rect 2702 3202 2705 3208
rect 3416 3203 3418 3207
rect 3422 3203 3425 3207
rect 3430 3203 3432 3207
rect 4440 3203 4442 3207
rect 4446 3203 4449 3207
rect 4454 3203 4456 3207
rect 570 3198 894 3201
rect 898 3198 918 3201
rect 2818 3198 2822 3201
rect 426 3188 798 3191
rect 834 3188 854 3191
rect 1234 3188 1310 3191
rect 1314 3188 1430 3191
rect 2274 3188 2446 3191
rect 2554 3188 2710 3191
rect 2814 3188 2822 3191
rect 2826 3188 2838 3191
rect 3194 3188 3278 3191
rect 3938 3188 3950 3191
rect 4866 3188 4910 3191
rect 5274 3188 5294 3191
rect 42 3178 110 3181
rect 170 3178 366 3181
rect 370 3178 398 3181
rect 1226 3178 1238 3181
rect 1650 3178 1790 3181
rect 1794 3178 1870 3181
rect 1930 3178 2350 3181
rect 2354 3178 2374 3181
rect 2378 3178 2654 3181
rect 3010 3178 3254 3181
rect 3258 3178 3342 3181
rect 4426 3178 4870 3181
rect 4986 3178 5094 3181
rect 5282 3178 5294 3181
rect 6 3171 9 3178
rect 6 3168 22 3171
rect 138 3168 270 3171
rect 306 3168 318 3171
rect 322 3168 329 3171
rect 470 3171 473 3178
rect 442 3168 473 3171
rect 482 3168 526 3171
rect 946 3168 950 3171
rect 1002 3168 1182 3171
rect 1202 3168 1206 3171
rect 1282 3168 1286 3171
rect 1922 3168 1966 3171
rect 2178 3168 2425 3171
rect 2490 3168 2798 3171
rect 2802 3168 2806 3171
rect 2842 3168 2854 3171
rect 2890 3168 2966 3171
rect 3202 3168 3406 3171
rect 3410 3168 3462 3171
rect 3514 3168 3534 3171
rect 3538 3168 3574 3171
rect 4162 3168 4302 3171
rect 4306 3168 4550 3171
rect 4838 3168 4846 3171
rect 4850 3168 5030 3171
rect 5034 3168 5070 3171
rect 5246 3171 5249 3178
rect 5342 3171 5346 3172
rect 5246 3168 5346 3171
rect 58 3158 78 3161
rect 94 3161 97 3168
rect 94 3158 206 3161
rect 322 3158 374 3161
rect 458 3158 470 3161
rect 490 3158 542 3161
rect 546 3158 550 3161
rect 714 3158 966 3161
rect 970 3158 1062 3161
rect 1146 3158 1190 3161
rect 1218 3158 1246 3161
rect 1594 3158 1662 3161
rect 1718 3161 1721 3168
rect 1666 3158 1721 3161
rect 1866 3158 1926 3161
rect 1946 3158 2158 3161
rect 2210 3158 2326 3161
rect 2346 3158 2390 3161
rect 2422 3161 2425 3168
rect 2422 3158 2550 3161
rect 2690 3158 2766 3161
rect 2946 3158 3030 3161
rect 3138 3158 3174 3161
rect 3178 3158 3230 3161
rect 3234 3158 3294 3161
rect 3434 3158 3494 3161
rect 3570 3158 3598 3161
rect 4762 3158 4862 3161
rect 4874 3158 4878 3161
rect 4922 3158 5078 3161
rect 5082 3158 5198 3161
rect 5258 3158 5286 3161
rect 58 3148 94 3151
rect 98 3148 118 3151
rect 238 3151 241 3158
rect 238 3148 582 3151
rect 786 3148 1006 3151
rect 1250 3148 1270 3151
rect 1422 3151 1425 3158
rect 1410 3148 1425 3151
rect 1458 3148 1486 3151
rect 1514 3148 1534 3151
rect 1586 3148 1630 3151
rect 1714 3148 1742 3151
rect 1754 3148 1782 3151
rect 1834 3148 1958 3151
rect 1962 3148 2014 3151
rect 2194 3148 2262 3151
rect 2266 3148 2318 3151
rect 2506 3148 2526 3151
rect 2670 3151 2673 3158
rect 2670 3148 2758 3151
rect 2762 3148 2774 3151
rect 2986 3148 3014 3151
rect 3090 3148 3094 3151
rect 3338 3148 3358 3151
rect 3410 3148 3438 3151
rect 3458 3148 3558 3151
rect 3694 3151 3697 3158
rect 3666 3148 3697 3151
rect 3726 3148 3774 3151
rect 3894 3148 3950 3151
rect 4018 3148 4158 3151
rect 4186 3148 4270 3151
rect 4286 3151 4289 3158
rect 4350 3151 4353 3158
rect 4286 3148 4353 3151
rect 4662 3151 4665 3158
rect 4634 3148 4665 3151
rect 4794 3148 4934 3151
rect 5342 3151 5346 3152
rect 5218 3148 5346 3151
rect 34 3138 54 3141
rect 118 3138 126 3141
rect 142 3141 145 3148
rect 630 3142 633 3148
rect 130 3138 145 3141
rect 418 3138 422 3141
rect 482 3138 494 3141
rect 530 3138 558 3141
rect 690 3138 750 3141
rect 754 3138 774 3141
rect 882 3138 926 3141
rect 930 3138 966 3141
rect 994 3138 1166 3141
rect 1210 3138 1222 3141
rect 1226 3138 1262 3141
rect 1306 3138 1350 3141
rect 1434 3138 1518 3141
rect 1522 3138 1574 3141
rect 1618 3138 1694 3141
rect 1730 3140 1766 3141
rect 1726 3138 1766 3140
rect 1810 3138 1902 3141
rect 2382 3141 2385 3148
rect 2306 3138 2385 3141
rect 2390 3141 2393 3148
rect 2390 3138 2494 3141
rect 2626 3138 2678 3141
rect 2706 3138 2734 3141
rect 2818 3138 2822 3141
rect 3058 3138 3158 3141
rect 3190 3141 3193 3148
rect 3726 3142 3729 3148
rect 3870 3142 3873 3148
rect 3894 3142 3897 3148
rect 3162 3138 3262 3141
rect 3282 3138 3326 3141
rect 3370 3138 3430 3141
rect 3490 3138 3510 3141
rect 3994 3138 4006 3141
rect 4074 3138 4137 3141
rect 4226 3138 4230 3141
rect 4254 3138 4321 3141
rect 4774 3141 4777 3148
rect 4698 3138 4777 3141
rect 4922 3138 4942 3141
rect 5130 3138 5246 3141
rect 5250 3138 5262 3141
rect 574 3132 577 3138
rect 638 3132 641 3138
rect 686 3132 689 3138
rect 42 3128 70 3131
rect 290 3128 302 3131
rect 354 3128 374 3131
rect 378 3128 422 3131
rect 426 3128 438 3131
rect 474 3128 510 3131
rect 794 3128 902 3131
rect 1010 3128 1158 3131
rect 1162 3128 1182 3131
rect 1302 3131 1305 3138
rect 4134 3132 4137 3138
rect 4254 3132 4257 3138
rect 4318 3132 4321 3138
rect 1274 3128 1305 3131
rect 1338 3128 1350 3131
rect 1394 3128 1449 3131
rect 1514 3128 1518 3131
rect 1530 3128 1534 3131
rect 1538 3128 1670 3131
rect 2074 3128 2166 3131
rect 2298 3128 2358 3131
rect 2562 3128 2638 3131
rect 2642 3128 2718 3131
rect 2746 3128 3374 3131
rect 3442 3128 3590 3131
rect 3594 3128 3646 3131
rect 3778 3128 3830 3131
rect 3834 3128 3990 3131
rect 4146 3128 4254 3131
rect 4954 3128 5022 3131
rect 1446 3122 1449 3128
rect 4270 3122 4273 3128
rect 66 3118 86 3121
rect 154 3118 182 3121
rect 418 3118 422 3121
rect 538 3118 646 3121
rect 650 3118 670 3121
rect 826 3118 918 3121
rect 922 3118 974 3121
rect 986 3118 1078 3121
rect 1138 3118 1214 3121
rect 1298 3118 1374 3121
rect 1378 3118 1414 3121
rect 1514 3118 1550 3121
rect 1554 3118 1622 3121
rect 2210 3118 2510 3121
rect 2666 3118 2710 3121
rect 2722 3118 2830 3121
rect 2834 3118 3382 3121
rect 3450 3118 3582 3121
rect 3586 3118 3630 3121
rect 4514 3118 4622 3121
rect 4750 3121 4753 3128
rect 4750 3118 4942 3121
rect 4946 3118 4974 3121
rect 4978 3118 5038 3121
rect 5042 3118 5118 3121
rect 5122 3118 5142 3121
rect 178 3108 454 3111
rect 466 3108 574 3111
rect 578 3108 606 3111
rect 618 3108 670 3111
rect 1218 3108 1342 3111
rect 1346 3108 1366 3111
rect 1370 3108 1470 3111
rect 1482 3108 1582 3111
rect 1634 3108 1750 3111
rect 1754 3108 1782 3111
rect 2234 3108 2238 3111
rect 2250 3108 2302 3111
rect 2314 3108 2398 3111
rect 2450 3108 2550 3111
rect 2706 3108 2718 3111
rect 2930 3108 3038 3111
rect 3042 3108 3318 3111
rect 3322 3108 3390 3111
rect 3394 3108 3502 3111
rect 4090 3108 4262 3111
rect 4266 3108 4462 3111
rect 856 3103 858 3107
rect 862 3103 865 3107
rect 870 3103 872 3107
rect 1872 3103 1874 3107
rect 1878 3103 1881 3107
rect 1886 3103 1888 3107
rect 2904 3103 2906 3107
rect 2910 3103 2913 3107
rect 2918 3103 2920 3107
rect 3928 3103 3930 3107
rect 3934 3103 3937 3107
rect 3942 3103 3944 3107
rect 4952 3103 4954 3107
rect 4958 3103 4961 3107
rect 4966 3103 4968 3107
rect 18 3098 54 3101
rect 410 3098 478 3101
rect 834 3098 838 3101
rect 914 3098 942 3101
rect 946 3098 958 3101
rect 962 3098 990 3101
rect 1042 3098 1190 3101
rect 1194 3098 1238 3101
rect 1242 3098 1270 3101
rect 1410 3098 1438 3101
rect 1610 3098 1830 3101
rect 2082 3098 2094 3101
rect 2098 3098 2753 3101
rect 2954 3098 2982 3101
rect 3266 3098 3358 3101
rect 3882 3098 3910 3101
rect 2750 3092 2753 3098
rect 258 3088 286 3091
rect 618 3088 926 3091
rect 930 3088 950 3091
rect 954 3088 974 3091
rect 1042 3088 1550 3091
rect 1618 3088 1654 3091
rect 1722 3088 1750 3091
rect 1986 3088 1990 3091
rect 2002 3088 2334 3091
rect 2338 3088 2358 3091
rect 2754 3088 2798 3091
rect 2802 3088 3046 3091
rect 3242 3088 3246 3091
rect 3250 3088 3366 3091
rect 3818 3088 4014 3091
rect 4170 3088 4230 3091
rect 4234 3088 4438 3091
rect 4466 3088 4534 3091
rect 4554 3088 4638 3091
rect 4642 3088 4654 3091
rect 4686 3091 4689 3098
rect 4686 3088 4942 3091
rect 4946 3088 4958 3091
rect 5010 3088 5142 3091
rect 5146 3088 5254 3091
rect 82 3078 206 3081
rect 210 3078 254 3081
rect 410 3078 446 3081
rect 458 3078 614 3081
rect 802 3078 841 3081
rect 294 3071 297 3078
rect 838 3072 841 3078
rect 922 3078 1030 3081
rect 1098 3078 1150 3081
rect 1370 3078 1422 3081
rect 1426 3078 1526 3081
rect 1530 3078 1542 3081
rect 1954 3078 1990 3081
rect 1994 3078 2062 3081
rect 2066 3078 2126 3081
rect 2186 3078 2222 3081
rect 2330 3078 2366 3081
rect 2418 3078 2518 3081
rect 2954 3078 2974 3081
rect 2978 3078 2982 3081
rect 2994 3078 3054 3081
rect 3122 3078 3126 3081
rect 3146 3078 3310 3081
rect 3322 3078 3358 3081
rect 3398 3078 3430 3081
rect 3450 3078 3518 3081
rect 3546 3078 3550 3081
rect 3594 3078 3614 3081
rect 3618 3078 3638 3081
rect 4346 3078 4358 3081
rect 4442 3078 4590 3081
rect 4954 3078 5086 3081
rect 5250 3078 5262 3081
rect 918 3072 921 3078
rect 3398 3072 3401 3078
rect 294 3068 390 3071
rect 394 3068 422 3071
rect 674 3068 678 3071
rect 690 3068 750 3071
rect 786 3068 806 3071
rect 922 3068 958 3071
rect 994 3068 1094 3071
rect 1098 3068 1110 3071
rect 1218 3068 1414 3071
rect 1418 3068 1438 3071
rect 1466 3070 1489 3071
rect 1466 3068 1486 3070
rect 90 3058 102 3061
rect 106 3058 118 3061
rect 138 3058 238 3061
rect 354 3058 398 3061
rect 434 3058 446 3061
rect 494 3061 497 3068
rect 1538 3068 1654 3071
rect 1658 3068 1742 3071
rect 2010 3068 2086 3071
rect 2346 3068 2446 3071
rect 2626 3068 2662 3071
rect 2666 3068 2678 3071
rect 2714 3068 2718 3071
rect 2850 3068 2862 3071
rect 2970 3068 3006 3071
rect 3026 3068 3030 3071
rect 3126 3068 3326 3071
rect 3330 3068 3350 3071
rect 3378 3068 3398 3071
rect 3410 3068 3446 3071
rect 3450 3068 3462 3071
rect 3522 3068 3558 3071
rect 3602 3068 3622 3071
rect 3686 3068 3694 3071
rect 3782 3071 3785 3078
rect 3698 3068 3785 3071
rect 3850 3068 3905 3071
rect 3950 3071 3953 3078
rect 3914 3068 3953 3071
rect 4034 3068 4094 3071
rect 4306 3068 4366 3071
rect 4370 3068 4406 3071
rect 4498 3068 4510 3071
rect 4526 3068 4622 3071
rect 4722 3068 4846 3071
rect 4986 3068 5030 3071
rect 5270 3071 5273 3078
rect 5270 3068 5310 3071
rect 494 3058 550 3061
rect 674 3058 742 3061
rect 746 3058 774 3061
rect 778 3058 806 3061
rect 962 3058 1006 3061
rect 1042 3058 1054 3061
rect 1178 3058 1222 3061
rect 1234 3058 1254 3061
rect 1258 3058 1302 3061
rect 1314 3058 1382 3061
rect 1858 3058 1921 3061
rect 2026 3058 2054 3061
rect 2090 3058 2158 3061
rect 2202 3058 2246 3061
rect 2354 3058 2366 3061
rect 2370 3058 2382 3061
rect 2570 3058 2598 3061
rect 2658 3058 2694 3061
rect 2810 3058 2902 3061
rect 2978 3058 2982 3061
rect 3126 3061 3129 3068
rect 3106 3058 3129 3061
rect 3138 3058 3206 3061
rect 3210 3058 3214 3061
rect 3226 3058 3262 3061
rect 3350 3061 3353 3068
rect 3902 3062 3905 3068
rect 4526 3062 4529 3068
rect 3350 3058 3486 3061
rect 3538 3058 3662 3061
rect 3666 3058 3686 3061
rect 3762 3058 3838 3061
rect 3930 3058 4006 3061
rect 4010 3058 4038 3061
rect 4042 3058 4054 3061
rect 4074 3058 4086 3061
rect 4162 3058 4166 3061
rect 4338 3058 4398 3061
rect 4402 3058 4417 3061
rect 4594 3058 4734 3061
rect 4866 3058 4942 3061
rect 5026 3058 5089 3061
rect 5282 3058 5302 3061
rect 574 3052 577 3058
rect 58 3048 78 3051
rect 114 3048 126 3051
rect 162 3048 198 3051
rect 202 3048 222 3051
rect 234 3048 278 3051
rect 426 3048 438 3051
rect 482 3048 502 3051
rect 506 3048 510 3051
rect 842 3048 846 3051
rect 850 3048 910 3051
rect 1002 3048 1006 3051
rect 1194 3048 1214 3051
rect 1234 3048 1241 3051
rect 1290 3048 1318 3051
rect 1330 3048 1390 3051
rect 1446 3051 1449 3058
rect 1718 3052 1721 3058
rect 1918 3052 1921 3058
rect 1446 3048 1470 3051
rect 1730 3048 1790 3051
rect 1794 3048 1902 3051
rect 1986 3048 2038 3051
rect 2050 3048 2110 3051
rect 2234 3048 2254 3051
rect 2366 3048 2422 3051
rect 2582 3048 2646 3051
rect 2866 3048 2878 3051
rect 2998 3051 3001 3058
rect 3870 3052 3873 3058
rect 4414 3052 4417 3058
rect 5086 3052 5089 3058
rect 2998 3048 3030 3051
rect 3186 3048 3222 3051
rect 3274 3048 3342 3051
rect 3354 3048 3398 3051
rect 3494 3048 3606 3051
rect 3610 3048 3622 3051
rect 3674 3048 3702 3051
rect 3706 3048 3846 3051
rect 3978 3048 3982 3051
rect 4050 3048 4110 3051
rect 4330 3048 4342 3051
rect 4434 3048 4542 3051
rect 4754 3048 4822 3051
rect 4826 3048 4830 3051
rect 4938 3048 5030 3051
rect 5234 3048 5270 3051
rect 5342 3051 5346 3052
rect 5314 3048 5346 3051
rect 1238 3042 1241 3048
rect 1326 3042 1329 3048
rect 2366 3042 2369 3048
rect 2582 3042 2585 3048
rect 3494 3042 3497 3048
rect 4278 3042 4281 3048
rect 74 3038 94 3041
rect 178 3038 238 3041
rect 250 3038 270 3041
rect 274 3038 406 3041
rect 674 3038 702 3041
rect 754 3038 886 3041
rect 1018 3038 1046 3041
rect 1066 3038 1078 3041
rect 1082 3038 1118 3041
rect 1242 3038 1294 3041
rect 1470 3038 1518 3041
rect 1826 3038 1830 3041
rect 1842 3038 1870 3041
rect 1874 3038 1902 3041
rect 1906 3038 2118 3041
rect 2978 3038 3198 3041
rect 3242 3038 3262 3041
rect 3370 3038 3398 3041
rect 3402 3038 3438 3041
rect 3458 3038 3462 3041
rect 3722 3038 3838 3041
rect 3842 3038 3894 3041
rect 4082 3038 4110 3041
rect 4114 3038 4158 3041
rect 4386 3038 4478 3041
rect 4482 3038 4494 3041
rect 1470 3032 1473 3038
rect 206 3028 222 3031
rect 234 3028 254 3031
rect 402 3028 558 3031
rect 1106 3028 1118 3031
rect 1122 3028 1134 3031
rect 1998 3028 2038 3031
rect 2378 3028 2774 3031
rect 3074 3028 3262 3031
rect 3266 3028 3310 3031
rect 3314 3028 3390 3031
rect 3398 3028 3598 3031
rect 3618 3028 3790 3031
rect 4162 3028 4190 3031
rect 4194 3028 4246 3031
rect 4250 3028 4318 3031
rect 5058 3028 5286 3031
rect 206 3022 209 3028
rect 1998 3022 2001 3028
rect 234 3018 902 3021
rect 978 3018 1230 3021
rect 2050 3018 2414 3021
rect 2610 3018 2982 3021
rect 3022 3021 3025 3028
rect 3398 3022 3401 3028
rect 4110 3022 4113 3028
rect 3022 3018 3382 3021
rect 5266 3018 5294 3021
rect 50 3008 62 3011
rect 2762 3008 2838 3011
rect 2842 3008 2854 3011
rect 2938 3008 3046 3011
rect 3058 3008 3398 3011
rect 344 3003 346 3007
rect 350 3003 353 3007
rect 358 3003 360 3007
rect 1368 3003 1370 3007
rect 1374 3003 1377 3007
rect 1382 3003 1384 3007
rect 2392 3003 2394 3007
rect 2398 3003 2401 3007
rect 2406 3003 2408 3007
rect 3416 3003 3418 3007
rect 3422 3003 3425 3007
rect 3430 3003 3432 3007
rect 4440 3003 4442 3007
rect 4446 3003 4449 3007
rect 4454 3003 4456 3007
rect 2026 2998 2070 3001
rect 2074 2998 2150 3001
rect 3034 2998 3134 3001
rect 3210 2998 3406 3001
rect 4306 2998 4318 3001
rect 482 2988 590 2991
rect 770 2988 782 2991
rect 1014 2991 1017 2998
rect 850 2988 1017 2991
rect 1478 2992 1481 2998
rect 1522 2988 1574 2991
rect 2066 2988 2078 2991
rect 2394 2988 2958 2991
rect 3118 2988 3126 2991
rect 3130 2988 3366 2991
rect 3386 2988 3486 2991
rect 3634 2988 3678 2991
rect 4858 2988 4998 2991
rect 5034 2988 5134 2991
rect 742 2981 745 2988
rect 714 2978 745 2981
rect 2118 2981 2121 2988
rect 2118 2978 2166 2981
rect 2234 2978 2286 2981
rect 2642 2978 3078 2981
rect 3282 2978 3313 2981
rect 3330 2978 3374 2981
rect 3378 2978 3494 2981
rect 3502 2978 3510 2981
rect 3514 2978 3518 2981
rect 3530 2978 3734 2981
rect 3738 2978 3750 2981
rect 66 2968 158 2971
rect 270 2971 273 2978
rect 258 2968 273 2971
rect 766 2971 769 2978
rect 690 2968 769 2971
rect 1434 2968 1454 2971
rect 1850 2968 1862 2971
rect 1978 2968 2030 2971
rect 2086 2971 2089 2978
rect 3310 2972 3313 2978
rect 2086 2968 2262 2971
rect 2266 2968 2310 2971
rect 2562 2968 2694 2971
rect 2698 2968 2726 2971
rect 2898 2968 3254 2971
rect 3258 2968 3294 2971
rect 3346 2968 3350 2971
rect 3426 2968 3534 2971
rect 3766 2971 3769 2978
rect 3766 2968 3798 2971
rect 4514 2968 4542 2971
rect 5054 2971 5057 2978
rect 5054 2968 5310 2971
rect 50 2958 86 2961
rect 158 2961 161 2968
rect 138 2958 161 2961
rect 190 2961 193 2968
rect 190 2958 222 2961
rect 274 2958 294 2961
rect 382 2961 385 2968
rect 298 2958 385 2961
rect 410 2958 446 2961
rect 562 2958 582 2961
rect 586 2958 878 2961
rect 1146 2958 1166 2961
rect 1170 2958 1222 2961
rect 1226 2958 1342 2961
rect 1410 2958 1566 2961
rect 1814 2961 1817 2968
rect 1794 2958 1817 2961
rect 1962 2958 2006 2961
rect 2042 2958 2062 2961
rect 2114 2958 2126 2961
rect 2162 2958 2198 2961
rect 2202 2958 2214 2961
rect 2290 2958 2294 2961
rect 2466 2958 2513 2961
rect 2530 2958 2582 2961
rect 2586 2958 2614 2961
rect 2690 2958 2734 2961
rect 3042 2958 3070 2961
rect 3074 2958 3118 2961
rect 3122 2958 3126 2961
rect 3138 2958 3174 2961
rect 3178 2958 3222 2961
rect 3294 2961 3297 2968
rect 3582 2962 3585 2968
rect 3294 2958 3382 2961
rect 3386 2958 3406 2961
rect 3418 2958 3470 2961
rect 3618 2958 3622 2961
rect 3674 2958 3702 2961
rect 3706 2958 3806 2961
rect 4090 2958 4134 2961
rect 4450 2958 4518 2961
rect 4522 2958 4574 2961
rect 74 2948 86 2951
rect 154 2948 198 2951
rect 202 2948 230 2951
rect 250 2948 334 2951
rect 370 2948 382 2951
rect 482 2948 526 2951
rect 530 2948 566 2951
rect 698 2948 726 2951
rect 738 2948 758 2951
rect 854 2948 862 2951
rect 966 2951 969 2958
rect 966 2948 1006 2951
rect 1130 2948 1142 2951
rect 1162 2948 1198 2951
rect 1554 2948 1617 2951
rect 662 2942 665 2948
rect 854 2942 857 2948
rect 122 2938 142 2941
rect 162 2938 294 2941
rect 318 2938 422 2941
rect 426 2938 550 2941
rect 722 2938 766 2941
rect 770 2938 782 2941
rect 870 2941 873 2948
rect 1078 2942 1081 2948
rect 1294 2942 1297 2948
rect 1614 2942 1617 2948
rect 1646 2948 1654 2951
rect 1810 2948 1846 2951
rect 2006 2951 2009 2958
rect 2510 2952 2513 2958
rect 1986 2948 2009 2951
rect 2034 2948 2038 2951
rect 2050 2948 2086 2951
rect 2090 2948 2110 2951
rect 2118 2948 2150 2951
rect 2154 2948 2182 2951
rect 2226 2948 2238 2951
rect 2622 2951 2625 2958
rect 3222 2952 3225 2958
rect 2622 2948 2686 2951
rect 2690 2948 2702 2951
rect 2734 2948 2742 2951
rect 2810 2948 2870 2951
rect 2946 2948 2958 2951
rect 3050 2948 3086 2951
rect 3090 2948 3142 2951
rect 3306 2948 3326 2951
rect 3362 2948 3430 2951
rect 3442 2948 3486 2951
rect 3490 2948 3518 2951
rect 3522 2948 3550 2951
rect 3574 2951 3577 2958
rect 3562 2948 3630 2951
rect 3650 2948 3686 2951
rect 3722 2948 3734 2951
rect 3842 2948 3910 2951
rect 4006 2951 4009 2958
rect 4006 2948 4214 2951
rect 4218 2948 4246 2951
rect 4474 2948 4494 2951
rect 4782 2951 4785 2958
rect 4746 2948 4785 2951
rect 4986 2948 5054 2951
rect 5082 2948 5102 2951
rect 5106 2948 5142 2951
rect 5198 2951 5201 2958
rect 5170 2948 5201 2951
rect 5242 2948 5286 2951
rect 5342 2951 5346 2952
rect 5314 2948 5346 2951
rect 1646 2942 1649 2948
rect 1710 2942 1713 2948
rect 870 2938 934 2941
rect 1002 2938 1070 2941
rect 1202 2938 1206 2941
rect 1778 2938 1854 2941
rect 2118 2941 2121 2948
rect 1954 2938 2121 2941
rect 2138 2938 2158 2941
rect 2238 2938 2246 2941
rect 2250 2938 2278 2941
rect 2426 2938 2518 2941
rect 2586 2938 2590 2941
rect 2618 2938 2630 2941
rect 2718 2941 2721 2948
rect 2718 2938 2782 2941
rect 2802 2938 2886 2941
rect 3074 2938 3150 2941
rect 3194 2938 3198 2941
rect 3202 2938 3262 2941
rect 3322 2938 3334 2941
rect 3338 2938 3406 2941
rect 3410 2938 3470 2941
rect 3498 2938 3558 2941
rect 3618 2938 3662 2941
rect 3714 2938 3718 2941
rect 3738 2938 3846 2941
rect 4050 2938 4078 2941
rect 4350 2941 4353 2948
rect 4330 2938 4353 2941
rect 4466 2938 4526 2941
rect 4530 2938 4558 2941
rect 4702 2941 4705 2948
rect 4702 2938 4769 2941
rect 4962 2938 5006 2941
rect 5274 2938 5294 2941
rect 198 2932 201 2938
rect 318 2932 321 2938
rect 82 2928 198 2931
rect 282 2928 318 2931
rect 386 2928 390 2931
rect 450 2928 489 2931
rect 546 2928 550 2931
rect 762 2928 782 2931
rect 786 2928 937 2931
rect 998 2931 1001 2938
rect 946 2928 1001 2931
rect 1438 2931 1441 2938
rect 4766 2932 4769 2938
rect 1010 2928 1441 2931
rect 1794 2928 1918 2931
rect 1946 2928 1993 2931
rect 2162 2928 2318 2931
rect 2594 2928 2654 2931
rect 2674 2928 2766 2931
rect 2770 2928 2798 2931
rect 2802 2928 2878 2931
rect 2890 2928 3086 2931
rect 3234 2928 3238 2931
rect 3306 2928 3438 2931
rect 3450 2928 3470 2931
rect 3634 2928 3758 2931
rect 3906 2928 4070 2931
rect 4418 2928 4470 2931
rect 4474 2928 4558 2931
rect 4770 2928 5110 2931
rect 5114 2928 5182 2931
rect 5226 2928 5262 2931
rect 486 2922 489 2928
rect 58 2918 150 2921
rect 154 2918 206 2921
rect 346 2918 366 2921
rect 610 2918 686 2921
rect 698 2918 822 2921
rect 934 2921 937 2928
rect 1990 2922 1993 2928
rect 934 2918 1398 2921
rect 1810 2918 1926 2921
rect 2650 2918 2702 2921
rect 2706 2918 2822 2921
rect 2826 2918 2838 2921
rect 2850 2918 3142 2921
rect 3278 2921 3281 2928
rect 3278 2918 3366 2921
rect 3386 2918 3430 2921
rect 3434 2918 3454 2921
rect 3466 2918 3494 2921
rect 3562 2918 3638 2921
rect 3658 2918 3694 2921
rect 3698 2918 3798 2921
rect 3826 2918 3846 2921
rect 3850 2918 3950 2921
rect 3978 2918 4078 2921
rect 4210 2918 4214 2921
rect 4442 2918 4502 2921
rect 4506 2918 4606 2921
rect 4610 2918 4638 2921
rect 4950 2918 4958 2921
rect 4962 2918 5118 2921
rect 5130 2918 5254 2921
rect 5258 2918 5270 2921
rect 18 2908 22 2911
rect 206 2911 209 2918
rect 206 2908 398 2911
rect 402 2908 422 2911
rect 442 2908 494 2911
rect 506 2908 510 2911
rect 986 2908 1038 2911
rect 2298 2908 2342 2911
rect 2346 2908 2350 2911
rect 2618 2908 2894 2911
rect 3042 2908 3182 2911
rect 3218 2908 3278 2911
rect 3282 2908 3422 2911
rect 3466 2908 3598 2911
rect 3602 2908 3622 2911
rect 3638 2911 3641 2918
rect 3638 2908 3830 2911
rect 4042 2908 4054 2911
rect 4058 2908 4142 2911
rect 5234 2908 5286 2911
rect 856 2903 858 2907
rect 862 2903 865 2907
rect 870 2903 872 2907
rect 1872 2903 1874 2907
rect 1878 2903 1881 2907
rect 1886 2903 1888 2907
rect 2904 2903 2906 2907
rect 2910 2903 2913 2907
rect 2918 2903 2920 2907
rect 3928 2903 3930 2907
rect 3934 2903 3937 2907
rect 3942 2903 3944 2907
rect 4952 2903 4954 2907
rect 4958 2903 4961 2907
rect 4966 2903 4968 2907
rect 258 2898 310 2901
rect 746 2898 838 2901
rect 914 2898 934 2901
rect 1910 2898 2070 2901
rect 2130 2898 2142 2901
rect 2306 2898 2638 2901
rect 3106 2898 3246 2901
rect 3250 2898 3302 2901
rect 3442 2898 3638 2901
rect 3718 2898 3734 2901
rect 3746 2898 3921 2901
rect 106 2888 166 2891
rect 170 2888 190 2891
rect 282 2888 590 2891
rect 594 2888 630 2891
rect 738 2888 766 2891
rect 1074 2888 1094 2891
rect 1234 2888 1238 2891
rect 1410 2888 1414 2891
rect 1578 2888 1582 2891
rect 1650 2888 1678 2891
rect 1682 2888 1798 2891
rect 1862 2888 1870 2891
rect 1910 2891 1913 2898
rect 1874 2888 1913 2891
rect 1922 2888 1950 2891
rect 2034 2888 2038 2891
rect 2042 2888 2054 2891
rect 2058 2888 2102 2891
rect 2106 2888 2262 2891
rect 2562 2888 2566 2891
rect 2946 2888 2998 2891
rect 3002 2888 3134 2891
rect 3154 2888 3470 2891
rect 3718 2891 3721 2898
rect 3570 2888 3721 2891
rect 3730 2888 3846 2891
rect 3918 2891 3921 2898
rect 5306 2898 5358 2901
rect 3918 2888 4046 2891
rect 4122 2888 4230 2891
rect 4546 2888 4670 2891
rect 4674 2888 4750 2891
rect 5078 2891 5081 2898
rect 5042 2888 5081 2891
rect 90 2878 150 2881
rect 154 2878 158 2881
rect 426 2878 742 2881
rect 922 2878 1014 2881
rect 1018 2878 1078 2881
rect 1082 2878 1182 2881
rect 1658 2878 1694 2881
rect 1698 2878 1894 2881
rect 1898 2878 2062 2881
rect 2066 2878 2142 2881
rect 2146 2878 2166 2881
rect 2178 2878 2302 2881
rect 2338 2878 2422 2881
rect 2426 2878 2638 2881
rect 3130 2878 3209 2881
rect 3282 2878 3294 2881
rect 3314 2878 3438 2881
rect 3586 2878 3654 2881
rect 3714 2878 3782 2881
rect 3970 2878 4014 2881
rect 4086 2881 4089 2888
rect 4018 2878 4089 2881
rect 4094 2881 4097 2888
rect 4094 2878 4142 2881
rect 4498 2878 4598 2881
rect 4602 2878 4614 2881
rect 4858 2878 4886 2881
rect 4914 2878 4942 2881
rect 4946 2878 4990 2881
rect 4994 2878 5014 2881
rect 294 2871 297 2878
rect 294 2868 454 2871
rect 666 2868 806 2871
rect 1182 2871 1185 2878
rect 1182 2868 1254 2871
rect 1378 2868 1438 2871
rect 1594 2868 1638 2871
rect 1642 2868 1662 2871
rect 1714 2868 1806 2871
rect 1834 2868 1846 2871
rect 1934 2868 1977 2871
rect 1986 2868 2078 2871
rect 2082 2868 2110 2871
rect 2162 2868 2174 2871
rect 2286 2868 2334 2871
rect 2562 2868 2566 2871
rect 2650 2868 2678 2871
rect 2682 2868 2686 2871
rect 2734 2868 2742 2871
rect 2746 2868 2774 2871
rect 2794 2868 2862 2871
rect 3006 2871 3009 2878
rect 3206 2872 3209 2878
rect 2922 2868 3022 2871
rect 3258 2868 3366 2871
rect 3698 2868 3806 2871
rect 3810 2868 3814 2871
rect 3874 2868 3894 2871
rect 3994 2868 4110 2871
rect 4154 2868 4214 2871
rect 4218 2868 4278 2871
rect 4594 2868 4694 2871
rect 4698 2868 4726 2871
rect 4730 2868 4790 2871
rect 4834 2868 4918 2871
rect 4922 2868 4982 2871
rect 4986 2868 5038 2871
rect 5042 2868 5174 2871
rect 5342 2871 5346 2872
rect 5226 2868 5346 2871
rect 58 2858 102 2861
rect 170 2858 278 2861
rect 346 2858 398 2861
rect 434 2858 438 2861
rect 634 2858 654 2861
rect 998 2858 1006 2861
rect 1218 2858 1230 2861
rect 1306 2858 1326 2861
rect 1330 2858 1390 2861
rect 1450 2858 1502 2861
rect 1570 2858 1606 2861
rect 1610 2858 1614 2861
rect 1666 2858 1718 2861
rect 1762 2858 1766 2861
rect 1934 2861 1937 2868
rect 1974 2862 1977 2868
rect 2246 2862 2249 2868
rect 2286 2862 2289 2868
rect 1802 2858 1937 2861
rect 1946 2858 1966 2861
rect 1978 2858 2022 2861
rect 2050 2858 2094 2861
rect 2130 2858 2198 2861
rect 2382 2861 2385 2868
rect 2362 2858 2385 2861
rect 2586 2858 2598 2861
rect 2630 2861 2633 2868
rect 2630 2858 2662 2861
rect 2666 2858 2734 2861
rect 2818 2858 2894 2861
rect 2898 2858 2926 2861
rect 2986 2858 3078 2861
rect 3114 2858 3134 2861
rect 3138 2858 3142 2861
rect 3202 2858 3238 2861
rect 3266 2858 3326 2861
rect 3458 2858 3470 2861
rect 3474 2858 3510 2861
rect 3674 2858 3678 2861
rect 3738 2858 3958 2861
rect 3978 2858 4038 2861
rect 4138 2858 4174 2861
rect 4362 2858 4374 2861
rect 4642 2858 4686 2861
rect 4690 2858 4718 2861
rect 4722 2858 4774 2861
rect 4874 2858 4902 2861
rect 4906 2858 4934 2861
rect 4938 2858 5062 2861
rect 138 2848 174 2851
rect 178 2848 254 2851
rect 798 2851 801 2858
rect 778 2848 801 2851
rect 902 2852 905 2858
rect 998 2852 1001 2858
rect 1170 2848 1390 2851
rect 1634 2848 1678 2851
rect 1738 2848 1774 2851
rect 1850 2848 1862 2851
rect 2126 2851 2129 2858
rect 1906 2848 2129 2851
rect 2322 2848 2334 2851
rect 2366 2848 2454 2851
rect 2682 2848 2686 2851
rect 2778 2848 2878 2851
rect 2882 2848 2918 2851
rect 2970 2848 2990 2851
rect 3018 2848 3022 2851
rect 3050 2848 3126 2851
rect 3194 2848 3198 2851
rect 3210 2848 3257 2851
rect 3386 2848 3542 2851
rect 3642 2848 3646 2851
rect 3650 2848 3670 2851
rect 3866 2848 4110 2851
rect 4170 2848 4198 2851
rect 4202 2848 4286 2851
rect 4578 2848 4622 2851
rect 4818 2848 4942 2851
rect 4954 2848 4998 2851
rect 5002 2848 5022 2851
rect 5026 2848 5049 2851
rect 5342 2851 5346 2852
rect 5290 2848 5346 2851
rect 682 2838 686 2841
rect 690 2838 918 2841
rect 1098 2838 1318 2841
rect 1558 2841 1561 2848
rect 2366 2842 2369 2848
rect 1558 2838 1766 2841
rect 1770 2838 1814 2841
rect 1858 2838 1998 2841
rect 2010 2838 2038 2841
rect 2058 2838 2062 2841
rect 2154 2838 2190 2841
rect 2194 2838 2342 2841
rect 2630 2841 2633 2848
rect 2670 2841 2673 2848
rect 2630 2838 2673 2841
rect 2686 2838 2758 2841
rect 2802 2838 2806 2841
rect 2826 2838 2830 2841
rect 2834 2838 2846 2841
rect 2866 2838 2886 2841
rect 2942 2841 2945 2848
rect 3254 2842 3257 2848
rect 2942 2838 3086 2841
rect 3618 2838 3686 2841
rect 3770 2838 3918 2841
rect 3922 2838 3942 2841
rect 3946 2838 3974 2841
rect 4002 2838 4022 2841
rect 4142 2841 4145 2848
rect 4050 2838 4145 2841
rect 4574 2841 4577 2848
rect 5046 2842 5049 2848
rect 4574 2838 4582 2841
rect 4602 2838 4646 2841
rect 4650 2838 4742 2841
rect 2686 2832 2689 2838
rect 106 2828 414 2831
rect 418 2828 606 2831
rect 674 2828 1286 2831
rect 1298 2828 1654 2831
rect 1746 2828 1926 2831
rect 2098 2828 2366 2831
rect 2874 2828 2894 2831
rect 2898 2828 2950 2831
rect 2954 2828 2974 2831
rect 3226 2828 3270 2831
rect 3698 2828 3878 2831
rect 3882 2828 3990 2831
rect 4018 2828 4030 2831
rect 4074 2828 4494 2831
rect 4570 2828 4710 2831
rect 4714 2828 4758 2831
rect 4890 2828 5222 2831
rect 194 2818 374 2821
rect 378 2818 470 2821
rect 578 2818 1174 2821
rect 1474 2818 1790 2821
rect 2026 2818 2182 2821
rect 2234 2818 2622 2821
rect 2626 2818 2654 2821
rect 2658 2818 2750 2821
rect 2754 2818 3534 2821
rect 3538 2818 3614 2821
rect 3786 2818 3998 2821
rect 4018 2818 4190 2821
rect 4194 2818 4270 2821
rect 2514 2808 2518 2811
rect 2706 2808 2726 2811
rect 3154 2808 3230 2811
rect 3234 2808 3334 2811
rect 3474 2808 3494 2811
rect 3954 2808 4030 2811
rect 4042 2808 4078 2811
rect 4082 2808 4310 2811
rect 344 2803 346 2807
rect 350 2803 353 2807
rect 358 2803 360 2807
rect 1368 2803 1370 2807
rect 1374 2803 1377 2807
rect 1382 2803 1384 2807
rect 2392 2803 2394 2807
rect 2398 2803 2401 2807
rect 2406 2803 2408 2807
rect 3022 2802 3025 2808
rect 3416 2803 3418 2807
rect 3422 2803 3425 2807
rect 3430 2803 3432 2807
rect 4440 2803 4442 2807
rect 4446 2803 4449 2807
rect 4454 2803 4456 2807
rect 450 2798 910 2801
rect 1650 2798 1782 2801
rect 1786 2798 1878 2801
rect 1882 2798 1934 2801
rect 2058 2798 2374 2801
rect 2378 2798 2385 2801
rect 2602 2798 2614 2801
rect 2786 2798 2926 2801
rect 3170 2798 3222 2801
rect 3754 2798 4358 2801
rect 170 2788 638 2791
rect 1338 2788 1350 2791
rect 1770 2788 1838 2791
rect 1842 2788 1902 2791
rect 2058 2788 2118 2791
rect 2258 2788 2302 2791
rect 2382 2791 2385 2798
rect 2382 2788 3118 2791
rect 3122 2788 3454 2791
rect 3458 2788 3710 2791
rect 4086 2788 4094 2791
rect 4098 2788 4430 2791
rect 4434 2788 4518 2791
rect 1650 2778 1654 2781
rect 1826 2778 1838 2781
rect 1922 2778 1974 2781
rect 2226 2778 2470 2781
rect 2482 2778 2630 2781
rect 3154 2778 3174 2781
rect 3178 2778 3198 2781
rect 3218 2778 3310 2781
rect 3886 2778 4046 2781
rect 4050 2778 4134 2781
rect 4698 2778 4718 2781
rect 90 2768 94 2771
rect 262 2771 265 2778
rect 302 2771 305 2778
rect 262 2768 350 2771
rect 354 2768 414 2771
rect 490 2768 534 2771
rect 738 2768 1134 2771
rect 1546 2768 1702 2771
rect 1834 2768 1958 2771
rect 2002 2768 2022 2771
rect 2346 2768 2374 2771
rect 2434 2768 2518 2771
rect 2834 2768 2854 2771
rect 2914 2768 2926 2771
rect 2958 2771 2961 2778
rect 2958 2768 2990 2771
rect 2994 2768 3030 2771
rect 3130 2768 3254 2771
rect 3738 2768 3766 2771
rect 3774 2771 3777 2778
rect 3770 2768 3777 2771
rect 3798 2771 3801 2778
rect 3886 2772 3889 2778
rect 3798 2768 3886 2771
rect 3978 2768 4022 2771
rect 4390 2771 4393 2778
rect 4390 2768 4398 2771
rect 4418 2768 4598 2771
rect 4602 2768 4630 2771
rect 4634 2768 4678 2771
rect 4882 2768 4990 2771
rect 5138 2768 5278 2771
rect 54 2761 57 2768
rect 54 2758 142 2761
rect 146 2758 174 2761
rect 238 2761 241 2768
rect 238 2758 278 2761
rect 802 2758 846 2761
rect 1186 2758 1206 2761
rect 1458 2758 1494 2761
rect 1586 2758 1670 2761
rect 1758 2761 1761 2768
rect 1758 2758 1830 2761
rect 1842 2758 1950 2761
rect 1954 2758 1998 2761
rect 2010 2758 2142 2761
rect 2314 2758 2326 2761
rect 2346 2758 2374 2761
rect 2378 2758 2398 2761
rect 2474 2758 2734 2761
rect 2802 2758 2822 2761
rect 2850 2758 2870 2761
rect 2874 2758 2918 2761
rect 3410 2758 3486 2761
rect 3602 2758 3606 2761
rect 3642 2758 3662 2761
rect 3682 2758 3694 2761
rect 3714 2758 3782 2761
rect 3858 2758 3966 2761
rect 3970 2758 3998 2761
rect 4062 2761 4065 2768
rect 4062 2758 4094 2761
rect 4362 2758 4430 2761
rect 4458 2758 4502 2761
rect 4506 2758 4526 2761
rect 4710 2761 4713 2768
rect 4710 2758 4726 2761
rect 4746 2758 4862 2761
rect 4898 2758 5086 2761
rect 5218 2758 5270 2761
rect 34 2748 62 2751
rect 86 2748 110 2751
rect 114 2748 262 2751
rect 346 2748 366 2751
rect 370 2748 430 2751
rect 494 2751 497 2758
rect 434 2748 497 2751
rect 678 2751 681 2758
rect 594 2748 681 2751
rect 754 2748 766 2751
rect 786 2748 902 2751
rect 906 2748 950 2751
rect 978 2748 982 2751
rect 1118 2751 1121 2758
rect 1090 2748 1222 2751
rect 1250 2748 1262 2751
rect 1522 2748 1542 2751
rect 1610 2748 1726 2751
rect 1778 2748 1910 2751
rect 1946 2748 2070 2751
rect 2178 2748 2182 2751
rect 86 2742 89 2748
rect 50 2738 70 2741
rect 106 2738 174 2741
rect 178 2738 214 2741
rect 218 2738 246 2741
rect 250 2738 486 2741
rect 710 2742 713 2748
rect 522 2740 550 2741
rect 518 2738 550 2740
rect 554 2738 654 2741
rect 742 2738 806 2741
rect 830 2738 886 2741
rect 1162 2738 1182 2741
rect 1210 2738 1246 2741
rect 1438 2741 1441 2748
rect 1454 2741 1457 2748
rect 1250 2738 1257 2741
rect 1438 2738 1550 2741
rect 1566 2741 1569 2748
rect 1554 2738 1569 2741
rect 1714 2738 1782 2741
rect 1786 2738 1814 2741
rect 1938 2738 2046 2741
rect 2246 2741 2249 2758
rect 2354 2748 2366 2751
rect 2418 2748 2462 2751
rect 2514 2748 2553 2751
rect 2794 2748 2806 2751
rect 2810 2748 2838 2751
rect 2842 2748 2862 2751
rect 2882 2748 2950 2751
rect 2954 2748 2966 2751
rect 3138 2748 3169 2751
rect 3282 2748 3294 2751
rect 3394 2748 3406 2751
rect 3610 2748 3622 2751
rect 3626 2748 3702 2751
rect 3706 2748 3742 2751
rect 3754 2748 3814 2751
rect 3818 2748 3841 2751
rect 3850 2748 3870 2751
rect 3970 2748 3982 2751
rect 4050 2748 4094 2751
rect 4298 2748 4302 2751
rect 2130 2738 2249 2741
rect 2550 2742 2553 2748
rect 3166 2742 3169 2748
rect 3342 2742 3345 2748
rect 2634 2738 2638 2741
rect 2698 2738 2718 2741
rect 2834 2738 2990 2741
rect 2994 2738 3038 2741
rect 3178 2738 3206 2741
rect 3542 2741 3545 2748
rect 3490 2738 3545 2741
rect 3562 2738 3798 2741
rect 3802 2738 3822 2741
rect 3838 2741 3841 2748
rect 3894 2742 3897 2748
rect 3838 2738 3846 2741
rect 3858 2738 3873 2741
rect 3946 2738 4054 2741
rect 4106 2738 4134 2741
rect 4278 2741 4281 2748
rect 4506 2748 4510 2751
rect 4666 2748 4694 2751
rect 4738 2748 4798 2751
rect 4802 2748 4846 2751
rect 4930 2748 5006 2751
rect 5010 2748 5022 2751
rect 5098 2748 5102 2751
rect 5342 2751 5346 2752
rect 5106 2748 5346 2751
rect 4234 2738 4281 2741
rect 4386 2738 4462 2741
rect 4534 2741 4537 2748
rect 4498 2738 4537 2741
rect 4554 2738 4574 2741
rect 4578 2738 4622 2741
rect 4810 2738 4822 2741
rect 4898 2738 4902 2741
rect 4906 2738 4926 2741
rect 4970 2738 5070 2741
rect 5258 2738 5302 2741
rect 66 2728 78 2731
rect 154 2728 182 2731
rect 306 2728 326 2731
rect 346 2728 390 2731
rect 394 2728 422 2731
rect 426 2728 518 2731
rect 530 2728 606 2731
rect 742 2731 745 2738
rect 830 2732 833 2738
rect 1118 2732 1121 2738
rect 722 2728 745 2731
rect 810 2728 814 2731
rect 906 2728 966 2731
rect 970 2728 1094 2731
rect 1146 2728 1166 2731
rect 1274 2728 1318 2731
rect 1322 2728 1446 2731
rect 1450 2728 1518 2731
rect 1674 2728 1726 2731
rect 1730 2728 1798 2731
rect 1914 2728 1934 2731
rect 2058 2728 2062 2731
rect 2066 2728 2118 2731
rect 2138 2728 2678 2731
rect 2682 2728 2702 2731
rect 2858 2728 2966 2731
rect 2970 2728 3030 2731
rect 3054 2731 3057 2738
rect 3870 2732 3873 2738
rect 3042 2728 3057 2731
rect 3178 2728 3190 2731
rect 3194 2728 3286 2731
rect 3602 2728 3630 2731
rect 3690 2728 3718 2731
rect 3722 2728 3750 2731
rect 3782 2728 3814 2731
rect 4490 2728 4542 2731
rect 4618 2728 4638 2731
rect 4798 2731 4801 2738
rect 4754 2728 4801 2731
rect 4826 2728 4873 2731
rect 4898 2728 4942 2731
rect 4946 2728 5006 2731
rect 5010 2728 5022 2731
rect 742 2722 745 2728
rect 314 2718 358 2721
rect 362 2718 462 2721
rect 466 2718 638 2721
rect 794 2718 846 2721
rect 874 2718 926 2721
rect 930 2718 974 2721
rect 978 2718 982 2721
rect 1714 2718 1742 2721
rect 1802 2718 1830 2721
rect 1958 2721 1961 2728
rect 3782 2722 3785 2728
rect 4870 2722 4873 2728
rect 1958 2718 2126 2721
rect 2658 2718 2662 2721
rect 2986 2718 3062 2721
rect 3066 2718 3126 2721
rect 3130 2718 3158 2721
rect 3514 2718 3558 2721
rect 3570 2718 3638 2721
rect 3642 2718 3654 2721
rect 4274 2718 4374 2721
rect 4650 2718 4686 2721
rect 4762 2718 4790 2721
rect 4794 2718 4814 2721
rect 4918 2718 4926 2721
rect 4930 2718 4974 2721
rect 4978 2718 5030 2721
rect 3726 2712 3729 2718
rect 226 2708 254 2711
rect 258 2708 390 2711
rect 402 2708 766 2711
rect 890 2708 934 2711
rect 978 2708 1182 2711
rect 1266 2708 1454 2711
rect 1722 2708 1782 2711
rect 1938 2708 1966 2711
rect 2042 2708 2078 2711
rect 2346 2708 2806 2711
rect 2810 2708 2854 2711
rect 3162 2708 3246 2711
rect 3330 2708 3462 2711
rect 3466 2708 3582 2711
rect 3666 2708 3678 2711
rect 4714 2708 4822 2711
rect 856 2703 858 2707
rect 862 2703 865 2707
rect 870 2703 872 2707
rect 1872 2703 1874 2707
rect 1878 2703 1881 2707
rect 1886 2703 1888 2707
rect 2904 2703 2906 2707
rect 2910 2703 2913 2707
rect 2918 2703 2920 2707
rect 3928 2703 3930 2707
rect 3934 2703 3937 2707
rect 3942 2703 3944 2707
rect 4952 2703 4954 2707
rect 4958 2703 4961 2707
rect 4966 2703 4968 2707
rect 474 2698 558 2701
rect 898 2698 1006 2701
rect 1178 2698 1590 2701
rect 1802 2698 1814 2701
rect 1898 2698 1902 2701
rect 2106 2698 2638 2701
rect 2642 2698 2897 2701
rect 122 2688 150 2691
rect 330 2688 414 2691
rect 458 2688 582 2691
rect 786 2688 894 2691
rect 954 2688 1046 2691
rect 1122 2688 1126 2691
rect 1202 2688 1302 2691
rect 1530 2688 1734 2691
rect 1762 2688 1934 2691
rect 1938 2688 2070 2691
rect 2306 2688 2750 2691
rect 2894 2691 2897 2698
rect 3106 2698 3190 2701
rect 3226 2698 3230 2701
rect 3234 2698 3310 2701
rect 3378 2698 3806 2701
rect 3810 2698 3878 2701
rect 4674 2698 4678 2701
rect 4738 2698 4750 2701
rect 4786 2698 4846 2701
rect 5010 2698 5134 2701
rect 5274 2698 5278 2701
rect 3038 2691 3041 2698
rect 2894 2688 3033 2691
rect 3038 2688 3054 2691
rect 3450 2688 3454 2691
rect 3466 2688 3470 2691
rect 3594 2688 4206 2691
rect 4626 2688 4790 2691
rect 4794 2688 4814 2691
rect 5010 2688 5038 2691
rect 5050 2688 5142 2691
rect 5266 2688 5302 2691
rect 378 2678 414 2681
rect 434 2678 478 2681
rect 650 2678 654 2681
rect 658 2678 678 2681
rect 738 2678 982 2681
rect 1002 2678 1006 2681
rect 1058 2678 1062 2681
rect 1114 2678 1254 2681
rect 1258 2678 1326 2681
rect 1634 2678 1718 2681
rect 1722 2678 1814 2681
rect 2050 2678 2214 2681
rect 2266 2678 2278 2681
rect 2282 2678 2334 2681
rect 2426 2678 2526 2681
rect 2586 2678 2590 2681
rect 2634 2678 2654 2681
rect 2902 2678 3006 2681
rect 3030 2681 3033 2688
rect 3030 2678 3094 2681
rect 3098 2678 3118 2681
rect 3122 2678 3382 2681
rect 3786 2678 4086 2681
rect 4090 2678 4190 2681
rect 4194 2678 4230 2681
rect 4242 2678 4286 2681
rect 4602 2678 4638 2681
rect 4730 2678 4822 2681
rect 4858 2678 4878 2681
rect 5042 2678 5070 2681
rect 5298 2678 5302 2681
rect 70 2671 73 2678
rect 110 2671 113 2678
rect 166 2672 169 2678
rect 70 2668 113 2671
rect 122 2668 134 2671
rect 306 2668 342 2671
rect 386 2668 446 2671
rect 578 2668 582 2671
rect 666 2668 721 2671
rect 826 2668 838 2671
rect 922 2668 1022 2671
rect 1042 2668 1054 2671
rect 1090 2668 1094 2671
rect 1114 2668 1158 2671
rect 1170 2668 1214 2671
rect 1218 2668 1230 2671
rect 1238 2668 1246 2671
rect 1250 2668 1265 2671
rect 1346 2668 1366 2671
rect 1602 2668 1830 2671
rect 1926 2671 1929 2678
rect 1926 2668 1982 2671
rect 1986 2670 2017 2671
rect 1986 2668 2014 2670
rect 50 2658 78 2661
rect 98 2658 153 2661
rect 162 2658 198 2661
rect 202 2658 294 2661
rect 298 2658 310 2661
rect 410 2658 438 2661
rect 442 2658 470 2661
rect 534 2661 537 2668
rect 718 2662 721 2668
rect 1262 2662 1265 2668
rect 2066 2668 2070 2671
rect 2098 2668 2166 2671
rect 2254 2671 2257 2678
rect 2254 2668 2278 2671
rect 2282 2668 2286 2671
rect 2330 2668 2374 2671
rect 2406 2671 2409 2678
rect 2386 2668 2409 2671
rect 2902 2672 2905 2678
rect 3614 2672 3617 2678
rect 3178 2668 3214 2671
rect 3234 2668 3238 2671
rect 3258 2668 3294 2671
rect 3646 2671 3649 2678
rect 3634 2668 3649 2671
rect 3706 2668 3822 2671
rect 3826 2668 3830 2671
rect 4094 2668 4142 2671
rect 4162 2668 4262 2671
rect 4334 2668 4350 2671
rect 4382 2671 4385 2678
rect 4382 2668 4590 2671
rect 4594 2668 4622 2671
rect 4626 2668 4646 2671
rect 4722 2668 4734 2671
rect 4882 2668 4910 2671
rect 4994 2668 5046 2671
rect 5050 2668 5054 2671
rect 5058 2668 5182 2671
rect 5290 2668 5294 2671
rect 4094 2662 4097 2668
rect 4334 2662 4337 2668
rect 534 2658 550 2661
rect 674 2658 694 2661
rect 898 2658 942 2661
rect 962 2658 990 2661
rect 1050 2658 1078 2661
rect 1130 2658 1134 2661
rect 1218 2658 1254 2661
rect 1658 2658 1918 2661
rect 1922 2658 1934 2661
rect 1962 2658 1982 2661
rect 1986 2658 1990 2661
rect 2038 2658 2086 2661
rect 2130 2658 2174 2661
rect 2266 2658 2310 2661
rect 2386 2658 2550 2661
rect 2698 2658 2702 2661
rect 2794 2658 2878 2661
rect 2882 2658 2934 2661
rect 3194 2658 3310 2661
rect 3414 2658 3502 2661
rect 3522 2658 3526 2661
rect 3698 2658 3721 2661
rect 150 2651 153 2658
rect 806 2652 809 2658
rect 58 2648 129 2651
rect 150 2648 166 2651
rect 194 2648 262 2651
rect 282 2648 302 2651
rect 402 2648 422 2651
rect 426 2648 446 2651
rect 458 2648 502 2651
rect 546 2648 558 2651
rect 830 2651 833 2658
rect 810 2648 833 2651
rect 942 2651 945 2658
rect 2038 2652 2041 2658
rect 942 2648 966 2651
rect 1066 2648 1142 2651
rect 1210 2648 1286 2651
rect 1314 2648 1366 2651
rect 1674 2648 1702 2651
rect 1994 2648 1998 2651
rect 2138 2648 2206 2651
rect 2238 2651 2241 2658
rect 2210 2648 2241 2651
rect 2262 2651 2265 2658
rect 2366 2652 2369 2658
rect 2974 2652 2977 2658
rect 3414 2652 3417 2658
rect 3718 2652 3721 2658
rect 3866 2658 3918 2661
rect 4130 2658 4166 2661
rect 4170 2658 4302 2661
rect 4514 2658 4542 2661
rect 4690 2658 5150 2661
rect 5154 2658 5190 2661
rect 5298 2658 5302 2661
rect 2262 2648 2294 2651
rect 2306 2648 2350 2651
rect 2374 2648 2414 2651
rect 2450 2648 2454 2651
rect 3218 2648 3262 2651
rect 3282 2648 3305 2651
rect 3330 2648 3414 2651
rect 3650 2648 3654 2651
rect 3658 2648 3678 2651
rect 3862 2651 3865 2658
rect 3842 2648 3865 2651
rect 3902 2648 3926 2651
rect 4074 2648 4118 2651
rect 4226 2648 4238 2651
rect 4266 2648 4278 2651
rect 4282 2648 4326 2651
rect 4330 2648 4358 2651
rect 4578 2648 4606 2651
rect 4610 2648 4702 2651
rect 4898 2648 4910 2651
rect 5002 2648 5025 2651
rect 5074 2648 5126 2651
rect 5130 2648 5193 2651
rect 126 2642 129 2648
rect 146 2638 150 2641
rect 482 2638 1350 2641
rect 2374 2641 2377 2648
rect 3302 2642 3305 2648
rect 3902 2642 3905 2648
rect 1706 2638 2377 2641
rect 2386 2638 3174 2641
rect 3310 2638 3342 2641
rect 3858 2638 3902 2641
rect 4018 2638 4174 2641
rect 4218 2638 4254 2641
rect 4258 2638 4342 2641
rect 4646 2638 4710 2641
rect 4738 2638 4742 2641
rect 4862 2641 4865 2648
rect 5022 2642 5025 2648
rect 5190 2642 5193 2648
rect 5270 2642 5273 2648
rect 4862 2638 4894 2641
rect 5034 2638 5054 2641
rect 5106 2638 5110 2641
rect 5142 2638 5161 2641
rect 166 2632 169 2638
rect 258 2628 526 2631
rect 546 2628 646 2631
rect 890 2628 950 2631
rect 954 2628 961 2631
rect 970 2628 1118 2631
rect 1122 2628 1270 2631
rect 1274 2628 1302 2631
rect 1698 2628 1990 2631
rect 1998 2628 2054 2631
rect 2114 2628 2246 2631
rect 2250 2628 2334 2631
rect 2338 2628 2422 2631
rect 2426 2628 2438 2631
rect 2586 2628 2598 2631
rect 2602 2628 2742 2631
rect 2746 2628 2838 2631
rect 2842 2628 2910 2631
rect 2914 2628 2958 2631
rect 3066 2628 3150 2631
rect 3226 2628 3294 2631
rect 3310 2631 3313 2638
rect 4646 2632 4649 2638
rect 3298 2628 3313 2631
rect 3330 2628 3982 2631
rect 3986 2628 3998 2631
rect 4202 2628 4534 2631
rect 4682 2628 4990 2631
rect 5134 2631 5137 2638
rect 4994 2628 5137 2631
rect 5142 2632 5145 2638
rect 5158 2632 5161 2638
rect 5234 2628 5294 2631
rect 1998 2622 2001 2628
rect 122 2618 1214 2621
rect 1282 2618 1310 2621
rect 1434 2618 1974 2621
rect 2018 2618 2406 2621
rect 2746 2618 2790 2621
rect 2946 2618 2982 2621
rect 2986 2618 3054 2621
rect 3266 2618 3630 2621
rect 4338 2618 4414 2621
rect 4418 2618 4462 2621
rect 4642 2618 4902 2621
rect 10 2608 14 2611
rect 98 2608 206 2611
rect 626 2608 1006 2611
rect 1082 2608 1110 2611
rect 1130 2608 1134 2611
rect 1394 2608 2206 2611
rect 2658 2608 3382 2611
rect 4538 2608 4886 2611
rect 5242 2608 5270 2611
rect 344 2603 346 2607
rect 350 2603 353 2607
rect 358 2603 360 2607
rect 1368 2603 1370 2607
rect 1374 2603 1377 2607
rect 1382 2603 1384 2607
rect 2392 2603 2394 2607
rect 2398 2603 2401 2607
rect 2406 2603 2408 2607
rect 3416 2603 3418 2607
rect 3422 2603 3425 2607
rect 3430 2603 3432 2607
rect 4440 2603 4442 2607
rect 4446 2603 4449 2607
rect 4454 2603 4456 2607
rect 722 2598 742 2601
rect 802 2598 846 2601
rect 1466 2598 1734 2601
rect 3018 2598 3030 2601
rect 3114 2598 3126 2601
rect 3610 2598 4070 2601
rect 4802 2598 4846 2601
rect 4850 2598 4982 2601
rect 1750 2592 1753 2598
rect 1950 2592 1953 2598
rect 2142 2592 2145 2598
rect 346 2588 366 2591
rect 790 2588 998 2591
rect 1002 2588 1022 2591
rect 1202 2588 1246 2591
rect 1506 2588 1606 2591
rect 2518 2591 2521 2598
rect 2466 2588 2521 2591
rect 2662 2592 2665 2598
rect 2802 2588 3590 2591
rect 3706 2588 3710 2591
rect 3962 2588 4182 2591
rect 4658 2588 4758 2591
rect 486 2581 489 2588
rect 790 2582 793 2588
rect 274 2578 489 2581
rect 734 2578 742 2581
rect 746 2578 758 2581
rect 954 2578 1078 2581
rect 1114 2578 1118 2581
rect 1198 2581 1201 2588
rect 1122 2578 1201 2581
rect 1658 2578 1798 2581
rect 1954 2578 1958 2581
rect 1970 2578 2262 2581
rect 2270 2581 2273 2588
rect 2270 2578 2502 2581
rect 3842 2578 3982 2581
rect 4482 2578 4662 2581
rect 4682 2578 5102 2581
rect 34 2568 118 2571
rect 282 2568 310 2571
rect 714 2568 798 2571
rect 906 2568 1662 2571
rect 1818 2568 2614 2571
rect 3150 2571 3153 2578
rect 3130 2568 3153 2571
rect 3874 2568 4102 2571
rect 4394 2568 4422 2571
rect 4426 2568 4462 2571
rect 4506 2568 4622 2571
rect 4674 2568 4886 2571
rect 4946 2568 4982 2571
rect 4986 2568 4998 2571
rect 5138 2568 5198 2571
rect 66 2558 270 2561
rect 562 2558 582 2561
rect 586 2558 630 2561
rect 642 2558 742 2561
rect 786 2558 806 2561
rect 858 2558 862 2561
rect 986 2558 1102 2561
rect 1662 2561 1665 2568
rect 1662 2558 2206 2561
rect 2210 2558 2486 2561
rect 3082 2558 3102 2561
rect 3578 2558 3670 2561
rect 3682 2558 3862 2561
rect 3866 2558 3942 2561
rect 3946 2558 3982 2561
rect 3994 2558 4014 2561
rect 4026 2558 4030 2561
rect 4050 2558 4422 2561
rect 4426 2558 4494 2561
rect 4498 2558 4558 2561
rect 4582 2558 4590 2561
rect 4594 2558 4670 2561
rect 4714 2558 4718 2561
rect 4866 2558 4894 2561
rect 4938 2558 4966 2561
rect 4970 2558 5022 2561
rect 5026 2558 5094 2561
rect 5290 2558 5294 2561
rect 414 2552 417 2558
rect 670 2552 673 2558
rect 18 2548 22 2551
rect 26 2548 46 2551
rect 122 2548 158 2551
rect 306 2548 318 2551
rect 418 2548 518 2551
rect 554 2548 566 2551
rect 626 2548 662 2551
rect 778 2548 814 2551
rect 866 2548 902 2551
rect 1074 2548 1078 2551
rect 1298 2548 1390 2551
rect 1518 2551 1521 2558
rect 3198 2552 3201 2558
rect 3542 2552 3545 2558
rect 1518 2548 1822 2551
rect 1834 2548 1889 2551
rect 154 2538 166 2541
rect 202 2538 206 2541
rect 266 2538 310 2541
rect 506 2538 510 2541
rect 598 2538 686 2541
rect 746 2538 782 2541
rect 842 2538 910 2541
rect 990 2541 993 2548
rect 1886 2542 1889 2548
rect 2042 2548 2081 2551
rect 2022 2542 2025 2548
rect 2078 2542 2081 2548
rect 2238 2548 2294 2551
rect 2306 2548 2310 2551
rect 2238 2542 2241 2548
rect 2726 2548 2761 2551
rect 2850 2548 2870 2551
rect 2890 2548 2969 2551
rect 3066 2548 3086 2551
rect 3122 2548 3150 2551
rect 3670 2551 3673 2558
rect 3642 2548 3646 2551
rect 2726 2542 2729 2548
rect 2758 2542 2761 2548
rect 2966 2542 2969 2548
rect 3670 2548 3726 2551
rect 3890 2548 3910 2551
rect 4018 2548 4054 2551
rect 4130 2548 4134 2551
rect 4370 2548 4406 2551
rect 4410 2548 4526 2551
rect 4570 2548 4574 2551
rect 4690 2548 4830 2551
rect 4842 2548 4846 2551
rect 4874 2548 4990 2551
rect 5098 2548 5182 2551
rect 5258 2548 5289 2551
rect 4526 2542 4529 2548
rect 5286 2542 5289 2548
rect 914 2538 993 2541
rect 1082 2538 1094 2541
rect 1618 2538 1646 2541
rect 1682 2538 1686 2541
rect 2162 2538 2214 2541
rect 2410 2538 2478 2541
rect 2778 2538 2782 2541
rect 2818 2538 2838 2541
rect 2866 2538 2894 2541
rect 3042 2538 3070 2541
rect 3074 2538 3110 2541
rect 3666 2538 4198 2541
rect 4354 2538 4382 2541
rect 4402 2538 4422 2541
rect 4426 2538 4478 2541
rect 4626 2538 4678 2541
rect 4794 2538 4814 2541
rect 4826 2538 4838 2541
rect 4842 2538 4934 2541
rect 5018 2538 5161 2541
rect 5170 2538 5249 2541
rect 5306 2538 5310 2541
rect 134 2532 137 2538
rect 150 2532 153 2538
rect 598 2532 601 2538
rect 58 2528 118 2531
rect 194 2528 206 2531
rect 498 2528 502 2531
rect 618 2528 678 2531
rect 682 2528 790 2531
rect 810 2528 910 2531
rect 1058 2528 1254 2531
rect 1326 2531 1329 2538
rect 2254 2532 2257 2538
rect 2494 2532 2497 2538
rect 2790 2532 2793 2538
rect 1314 2528 1329 2531
rect 1338 2528 1678 2531
rect 1682 2528 1702 2531
rect 1754 2528 2150 2531
rect 3374 2531 3377 2538
rect 4246 2532 4249 2538
rect 5158 2532 5161 2538
rect 5246 2532 5249 2538
rect 3374 2528 3454 2531
rect 3706 2528 3742 2531
rect 3882 2528 3910 2531
rect 3914 2528 3950 2531
rect 3978 2528 4190 2531
rect 4514 2528 4590 2531
rect 4646 2528 4702 2531
rect 4706 2528 4734 2531
rect 4746 2528 4870 2531
rect 4918 2528 5014 2531
rect 5018 2528 5022 2531
rect 5266 2528 5302 2531
rect 114 2518 118 2521
rect 458 2518 518 2521
rect 682 2518 966 2521
rect 1002 2518 1022 2521
rect 1026 2518 1038 2521
rect 1194 2518 1318 2521
rect 1546 2518 1646 2521
rect 1650 2518 2246 2521
rect 2250 2518 2262 2521
rect 2362 2518 2558 2521
rect 2642 2518 2782 2521
rect 2814 2521 2817 2528
rect 2786 2518 2817 2521
rect 3154 2518 3750 2521
rect 3786 2518 3822 2521
rect 3826 2518 3958 2521
rect 3986 2518 4030 2521
rect 4034 2518 4038 2521
rect 4066 2518 4086 2521
rect 4162 2518 4246 2521
rect 4646 2521 4649 2528
rect 4434 2518 4649 2521
rect 4918 2521 4921 2528
rect 4770 2518 4921 2521
rect 4930 2518 4982 2521
rect 5106 2518 5270 2521
rect 5294 2512 5297 2518
rect 434 2508 454 2511
rect 706 2508 766 2511
rect 1090 2508 1102 2511
rect 1106 2508 1174 2511
rect 1282 2508 1334 2511
rect 1674 2508 1718 2511
rect 1898 2508 2246 2511
rect 2250 2508 2630 2511
rect 2634 2508 2750 2511
rect 2778 2508 2806 2511
rect 3346 2508 3470 2511
rect 3954 2508 3982 2511
rect 4394 2508 4534 2511
rect 4538 2508 4558 2511
rect 4562 2508 4614 2511
rect 4618 2508 4630 2511
rect 4738 2508 4878 2511
rect 4986 2508 5022 2511
rect 5026 2508 5102 2511
rect 5178 2508 5206 2511
rect 5210 2508 5262 2511
rect 5274 2508 5278 2511
rect 856 2503 858 2507
rect 862 2503 865 2507
rect 870 2503 872 2507
rect 1526 2502 1529 2508
rect 1872 2503 1874 2507
rect 1878 2503 1881 2507
rect 1886 2503 1888 2507
rect 2904 2503 2906 2507
rect 2910 2503 2913 2507
rect 2918 2503 2920 2507
rect 3246 2502 3249 2508
rect 3928 2503 3930 2507
rect 3934 2503 3937 2507
rect 3942 2503 3944 2507
rect 4190 2502 4193 2508
rect 4952 2503 4954 2507
rect 4958 2503 4961 2507
rect 4966 2503 4968 2507
rect 658 2498 670 2501
rect 1162 2498 1318 2501
rect 1802 2498 1822 2501
rect 2138 2498 2142 2501
rect 2162 2498 2182 2501
rect 2242 2498 2254 2501
rect 2498 2498 2582 2501
rect 2626 2498 2830 2501
rect 3042 2498 3054 2501
rect 3410 2498 3462 2501
rect 3466 2498 3478 2501
rect 3994 2498 4022 2501
rect 4026 2498 4062 2501
rect 4706 2498 4790 2501
rect 4794 2498 4806 2501
rect 5098 2498 5214 2501
rect 298 2488 374 2491
rect 514 2488 630 2491
rect 818 2488 830 2491
rect 834 2488 857 2491
rect 1098 2488 1134 2491
rect 1210 2488 1246 2491
rect 1250 2488 1305 2491
rect 1442 2488 3286 2491
rect 3290 2488 3294 2491
rect 3906 2488 3998 2491
rect 4018 2488 4238 2491
rect 4546 2488 4641 2491
rect 4770 2488 4814 2491
rect 4854 2488 5110 2491
rect 854 2482 857 2488
rect 1302 2482 1305 2488
rect 4638 2482 4641 2488
rect 4854 2482 4857 2488
rect 34 2478 86 2481
rect 114 2478 150 2481
rect 314 2478 358 2481
rect 738 2478 814 2481
rect 938 2478 950 2481
rect 954 2478 1126 2481
rect 1146 2478 1198 2481
rect 1202 2478 1294 2481
rect 1450 2478 1606 2481
rect 2106 2478 2158 2481
rect 2522 2478 2678 2481
rect 2794 2478 2846 2481
rect 2850 2478 2974 2481
rect 3014 2478 3086 2481
rect 3354 2478 3406 2481
rect 3410 2478 3446 2481
rect 3602 2478 3630 2481
rect 3634 2478 3686 2481
rect 3738 2478 3822 2481
rect 3882 2478 4014 2481
rect 4234 2478 4270 2481
rect 4490 2478 4582 2481
rect 4586 2478 4598 2481
rect 4666 2478 4726 2481
rect 4782 2478 4817 2481
rect 4898 2478 4934 2481
rect 4938 2478 5038 2481
rect 5082 2478 5086 2481
rect 5186 2478 5214 2481
rect 5218 2478 5302 2481
rect 82 2468 166 2471
rect 214 2471 217 2478
rect 1446 2472 1449 2478
rect 214 2468 246 2471
rect 282 2468 318 2471
rect 410 2468 497 2471
rect 682 2468 769 2471
rect 778 2468 798 2471
rect 842 2468 894 2471
rect 1490 2468 1518 2471
rect 1670 2468 1678 2471
rect 1682 2468 1718 2471
rect 1722 2468 1806 2471
rect 1810 2468 1854 2471
rect 1998 2471 2001 2478
rect 1954 2468 2001 2471
rect 2018 2468 2038 2471
rect 2146 2468 2150 2471
rect 2286 2471 2289 2478
rect 3014 2471 3017 2478
rect 4782 2472 4785 2478
rect 4814 2472 4817 2478
rect 2286 2468 3017 2471
rect 3026 2468 3169 2471
rect 3250 2468 3281 2471
rect 494 2462 497 2468
rect 66 2458 78 2461
rect 146 2458 190 2461
rect 194 2458 310 2461
rect 530 2458 574 2461
rect 706 2458 710 2461
rect 766 2461 769 2468
rect 766 2458 1046 2461
rect 1074 2458 1110 2461
rect 1122 2458 1158 2461
rect 1162 2458 1206 2461
rect 1250 2458 1262 2461
rect 1298 2458 1678 2461
rect 1738 2459 1758 2461
rect 1734 2458 1758 2459
rect 1802 2458 1806 2461
rect 3070 2462 3073 2468
rect 3166 2462 3169 2468
rect 3278 2462 3281 2468
rect 3490 2468 3534 2471
rect 3570 2468 3670 2471
rect 3802 2468 3974 2471
rect 3986 2468 4046 2471
rect 4194 2468 4222 2471
rect 4226 2468 4238 2471
rect 4250 2468 4313 2471
rect 4410 2468 4462 2471
rect 4506 2468 4510 2471
rect 4514 2468 4534 2471
rect 4594 2468 4614 2471
rect 4618 2468 4670 2471
rect 4682 2468 4777 2471
rect 4890 2468 4918 2471
rect 4922 2468 4958 2471
rect 5042 2468 5094 2471
rect 5158 2471 5161 2478
rect 5130 2468 5161 2471
rect 1882 2459 1886 2461
rect 1878 2458 1886 2459
rect 1970 2458 2022 2461
rect 2074 2458 3038 2461
rect 3366 2461 3369 2468
rect 3346 2458 3369 2461
rect 3530 2458 3534 2461
rect 3566 2461 3569 2468
rect 4310 2462 4313 2468
rect 3566 2458 3606 2461
rect 3634 2458 3646 2461
rect 3762 2458 3854 2461
rect 3874 2458 3894 2461
rect 3922 2458 3934 2461
rect 3954 2458 4030 2461
rect 4034 2458 4046 2461
rect 4098 2458 4214 2461
rect 4218 2458 4262 2461
rect 4514 2458 4566 2461
rect 4602 2458 4638 2461
rect 4642 2458 4694 2461
rect 4762 2458 4766 2461
rect 4774 2461 4777 2468
rect 5286 2462 5289 2468
rect 4774 2458 4830 2461
rect 5034 2458 5054 2461
rect 5058 2458 5086 2461
rect 5106 2458 5150 2461
rect 5154 2458 5190 2461
rect 486 2452 489 2458
rect 122 2448 158 2451
rect 274 2448 278 2451
rect 282 2448 334 2451
rect 722 2448 734 2451
rect 754 2448 774 2451
rect 898 2448 942 2451
rect 1210 2448 1230 2451
rect 1298 2448 1310 2451
rect 1322 2448 1790 2451
rect 1794 2448 2006 2451
rect 2018 2448 2070 2451
rect 2122 2448 2198 2451
rect 2226 2448 2302 2451
rect 2314 2448 2318 2451
rect 2354 2448 2414 2451
rect 2502 2448 2518 2451
rect 2674 2448 2678 2451
rect 2826 2448 3182 2451
rect 3314 2448 3342 2451
rect 3538 2448 3542 2451
rect 3546 2448 3582 2451
rect 3586 2448 3638 2451
rect 3722 2448 3806 2451
rect 3810 2448 3886 2451
rect 3890 2448 3910 2451
rect 4002 2448 4086 2451
rect 4090 2448 4118 2451
rect 4178 2448 4206 2451
rect 4210 2448 4222 2451
rect 4270 2448 4278 2451
rect 4282 2448 4358 2451
rect 4394 2448 4398 2451
rect 4402 2448 4422 2451
rect 4466 2448 4478 2451
rect 4482 2448 4518 2451
rect 4634 2448 4726 2451
rect 4730 2448 4750 2451
rect 5082 2448 5126 2451
rect 5130 2448 5142 2451
rect 5146 2448 5150 2451
rect 42 2438 62 2441
rect 138 2438 166 2441
rect 170 2438 294 2441
rect 314 2438 414 2441
rect 642 2438 686 2441
rect 690 2438 726 2441
rect 822 2441 825 2448
rect 810 2438 825 2441
rect 898 2438 918 2441
rect 1018 2438 1038 2441
rect 1178 2438 1278 2441
rect 1522 2438 1550 2441
rect 1554 2438 1574 2441
rect 1594 2438 1798 2441
rect 1802 2438 1822 2441
rect 2502 2441 2505 2448
rect 2622 2442 2625 2448
rect 2194 2438 2505 2441
rect 2514 2438 2518 2441
rect 2834 2438 2854 2441
rect 2986 2438 2990 2441
rect 3390 2441 3393 2448
rect 3386 2438 3393 2441
rect 3494 2441 3497 2448
rect 3494 2438 3502 2441
rect 3530 2438 3558 2441
rect 3630 2438 3726 2441
rect 3946 2438 4006 2441
rect 4074 2438 4209 2441
rect 4538 2438 4558 2441
rect 5066 2438 5078 2441
rect 5082 2438 5086 2441
rect 5098 2438 5110 2441
rect 682 2428 758 2431
rect 762 2428 790 2431
rect 818 2428 958 2431
rect 1382 2431 1385 2438
rect 1354 2428 1385 2431
rect 1570 2428 1598 2431
rect 1618 2428 1766 2431
rect 1778 2428 3326 2431
rect 3630 2431 3633 2438
rect 4206 2432 4209 2438
rect 3410 2428 3633 2431
rect 3642 2428 3742 2431
rect 3746 2428 3806 2431
rect 4146 2428 4190 2431
rect 202 2418 302 2421
rect 330 2418 342 2421
rect 382 2421 385 2428
rect 382 2418 502 2421
rect 850 2418 926 2421
rect 1330 2418 1926 2421
rect 2010 2418 2126 2421
rect 2170 2418 2526 2421
rect 2530 2418 2550 2421
rect 2850 2418 3526 2421
rect 4154 2418 4166 2421
rect 4402 2418 5054 2421
rect 18 2408 22 2411
rect 202 2408 222 2411
rect 386 2408 398 2411
rect 1426 2408 1710 2411
rect 1714 2408 2142 2411
rect 2154 2408 2158 2411
rect 2162 2408 2182 2411
rect 2482 2408 2782 2411
rect 2786 2408 2894 2411
rect 3730 2408 3934 2411
rect 3978 2408 4014 2411
rect 4018 2408 4174 2411
rect 5198 2411 5201 2418
rect 5198 2408 5206 2411
rect 344 2403 346 2407
rect 350 2403 353 2407
rect 358 2403 360 2407
rect 1368 2403 1370 2407
rect 1374 2403 1377 2407
rect 1382 2403 1384 2407
rect 2392 2403 2394 2407
rect 2398 2403 2401 2407
rect 2406 2403 2408 2407
rect 3416 2403 3418 2407
rect 3422 2403 3425 2407
rect 3430 2403 3432 2407
rect 4440 2403 4442 2407
rect 4446 2403 4449 2407
rect 4454 2403 4456 2407
rect 1042 2398 1126 2401
rect 1762 2398 1918 2401
rect 1930 2398 1966 2401
rect 1986 2398 2118 2401
rect 2130 2398 2190 2401
rect 2346 2398 2374 2401
rect 2786 2398 2798 2401
rect 2834 2398 2870 2401
rect 3458 2398 4350 2401
rect 5050 2398 5134 2401
rect 5138 2398 5182 2401
rect 354 2388 390 2391
rect 482 2388 486 2391
rect 490 2388 497 2391
rect 674 2388 766 2391
rect 770 2388 777 2391
rect 1034 2388 1486 2391
rect 390 2381 393 2388
rect 1710 2382 1713 2398
rect 1826 2388 2590 2391
rect 2610 2388 2614 2391
rect 3178 2388 3214 2391
rect 3218 2388 3342 2391
rect 3586 2388 3734 2391
rect 3802 2388 3830 2391
rect 4134 2388 4158 2391
rect 4322 2388 4326 2391
rect 4690 2388 4822 2391
rect 390 2378 798 2381
rect 802 2378 934 2381
rect 1058 2378 1062 2381
rect 1094 2378 1102 2381
rect 1106 2378 1118 2381
rect 1322 2378 1566 2381
rect 1730 2378 1750 2381
rect 1814 2381 1817 2388
rect 1814 2378 1830 2381
rect 1918 2378 1942 2381
rect 1994 2378 2006 2381
rect 2130 2378 2382 2381
rect 2674 2378 2710 2381
rect 2714 2378 2766 2381
rect 2770 2378 2950 2381
rect 2990 2381 2993 2388
rect 4134 2382 4137 2388
rect 2990 2378 3014 2381
rect 3018 2378 3054 2381
rect 3266 2378 3358 2381
rect 3698 2378 3766 2381
rect 3834 2378 3942 2381
rect 3954 2378 4054 2381
rect 4074 2378 4134 2381
rect 4674 2378 4758 2381
rect 4770 2378 4910 2381
rect 5214 2381 5217 2388
rect 5106 2378 5217 2381
rect 30 2371 33 2378
rect 1918 2372 1921 2378
rect 18 2368 118 2371
rect 426 2368 486 2371
rect 602 2368 622 2371
rect 682 2368 718 2371
rect 794 2368 862 2371
rect 986 2368 1014 2371
rect 1018 2368 1022 2371
rect 1074 2368 1182 2371
rect 1394 2368 1398 2371
rect 1610 2368 1694 2371
rect 1810 2368 1846 2371
rect 1850 2368 1886 2371
rect 1926 2368 2078 2371
rect 2082 2368 2374 2371
rect 2626 2368 2806 2371
rect 2914 2368 3198 2371
rect 3202 2368 3230 2371
rect 3482 2368 3518 2371
rect 3522 2368 3758 2371
rect 3970 2368 3982 2371
rect 4010 2368 4030 2371
rect 4034 2368 4062 2371
rect 4066 2368 4110 2371
rect 4130 2368 4270 2371
rect 4338 2368 4369 2371
rect 4498 2368 4534 2371
rect 4542 2371 4545 2378
rect 5062 2372 5065 2378
rect 4538 2368 4545 2371
rect 4738 2368 4750 2371
rect 4754 2368 4918 2371
rect 4962 2368 5022 2371
rect 5082 2368 5126 2371
rect 42 2358 118 2361
rect 198 2361 201 2368
rect 170 2358 201 2361
rect 258 2358 278 2361
rect 282 2358 646 2361
rect 698 2358 742 2361
rect 766 2361 769 2368
rect 754 2358 769 2361
rect 1010 2358 1014 2361
rect 1062 2358 1078 2361
rect 1482 2358 1662 2361
rect 1670 2358 1726 2361
rect 1742 2361 1745 2368
rect 1742 2358 1766 2361
rect 1926 2361 1929 2368
rect 1770 2358 1929 2361
rect 1946 2358 1950 2361
rect 1978 2358 1990 2361
rect 1994 2358 1998 2361
rect 2026 2358 2694 2361
rect 2698 2358 2734 2361
rect 2802 2358 2878 2361
rect 2882 2358 2950 2361
rect 2970 2358 3038 2361
rect 3042 2358 3062 2361
rect 3138 2358 3142 2361
rect 3154 2358 3206 2361
rect 3254 2361 3257 2368
rect 3210 2358 3257 2361
rect 3278 2361 3281 2368
rect 3274 2358 3281 2361
rect 3326 2361 3329 2368
rect 4366 2362 4369 2368
rect 3322 2358 3329 2361
rect 3346 2358 3350 2361
rect 3370 2358 3382 2361
rect 3498 2358 3622 2361
rect 3754 2358 3774 2361
rect 3786 2358 3822 2361
rect 3922 2358 3926 2361
rect 4098 2358 4118 2361
rect 4250 2358 4254 2361
rect 4282 2358 4302 2361
rect 4306 2358 4350 2361
rect 4370 2358 4398 2361
rect 4578 2358 4582 2361
rect 4738 2358 4766 2361
rect 4794 2358 4822 2361
rect 4834 2358 4865 2361
rect 5010 2358 5014 2361
rect 5066 2358 5150 2361
rect 5154 2358 5190 2361
rect 90 2348 150 2351
rect 210 2348 230 2351
rect 322 2348 374 2351
rect 418 2348 430 2351
rect 506 2348 518 2351
rect 618 2348 630 2351
rect 650 2348 726 2351
rect 786 2348 814 2351
rect 910 2351 913 2358
rect 1062 2352 1065 2358
rect 1462 2352 1465 2358
rect 1670 2352 1673 2358
rect 4862 2352 4865 2358
rect 910 2348 942 2351
rect 970 2348 998 2351
rect 1082 2348 1174 2351
rect 1498 2348 1502 2351
rect 1722 2348 1758 2351
rect 1818 2348 1822 2351
rect 1842 2348 1846 2351
rect 1858 2348 1894 2351
rect 1906 2348 1910 2351
rect 1938 2348 1942 2351
rect 2218 2348 2222 2351
rect 2250 2348 2281 2351
rect 2370 2348 2398 2351
rect 2506 2348 2510 2351
rect 2822 2348 2830 2351
rect 2890 2348 2926 2351
rect 2946 2348 3166 2351
rect 3170 2348 3270 2351
rect 3274 2348 3318 2351
rect 3370 2348 3398 2351
rect 3498 2348 3526 2351
rect 3594 2348 3614 2351
rect 3618 2348 3625 2351
rect 3650 2348 3678 2351
rect 3682 2348 3870 2351
rect 3978 2348 3985 2351
rect 86 2342 89 2348
rect 18 2338 86 2341
rect 114 2338 118 2341
rect 178 2338 222 2341
rect 226 2338 270 2341
rect 306 2338 326 2341
rect 370 2338 422 2341
rect 506 2338 510 2341
rect 642 2338 654 2341
rect 682 2338 742 2341
rect 746 2338 894 2341
rect 978 2338 1006 2341
rect 1010 2338 1054 2341
rect 1130 2338 1166 2341
rect 1270 2341 1273 2348
rect 1202 2338 1350 2341
rect 1582 2341 1585 2348
rect 2278 2342 2281 2348
rect 2822 2342 2825 2348
rect 1554 2338 1585 2341
rect 1634 2338 1638 2341
rect 1722 2338 1774 2341
rect 1810 2338 2030 2341
rect 2194 2338 2198 2341
rect 2218 2338 2225 2341
rect 2354 2338 2430 2341
rect 2858 2338 2862 2341
rect 2866 2340 2982 2341
rect 2986 2340 2998 2341
rect 2866 2338 2998 2340
rect 3034 2338 3078 2341
rect 3106 2338 3190 2341
rect 3194 2338 3278 2341
rect 3282 2338 3310 2341
rect 3362 2338 3374 2341
rect 3378 2338 3414 2341
rect 3522 2338 3526 2341
rect 3530 2338 3662 2341
rect 3666 2338 3710 2341
rect 3762 2338 3790 2341
rect 3794 2338 3854 2341
rect 3982 2342 3985 2348
rect 3998 2348 4046 2351
rect 4050 2348 4070 2351
rect 4074 2348 4078 2351
rect 4166 2348 4182 2351
rect 4266 2348 4809 2351
rect 4826 2348 4846 2351
rect 4890 2348 4894 2351
rect 5050 2348 5070 2351
rect 5082 2348 5086 2351
rect 5106 2348 5121 2351
rect 5218 2348 5286 2351
rect 3998 2342 4001 2348
rect 4166 2342 4169 2348
rect 3906 2340 3942 2341
rect 3902 2338 3942 2340
rect 4018 2338 4142 2341
rect 4210 2338 4278 2341
rect 4306 2338 4422 2341
rect 4426 2338 4470 2341
rect 4474 2338 4566 2341
rect 4570 2338 4590 2341
rect 4658 2338 4710 2341
rect 4722 2338 4798 2341
rect 4806 2341 4809 2348
rect 5118 2342 5121 2348
rect 4806 2338 4814 2341
rect 4834 2338 4838 2341
rect 4850 2338 4902 2341
rect 4986 2338 5006 2341
rect 5010 2338 5022 2341
rect 5026 2338 5094 2341
rect 5186 2338 5214 2341
rect 5282 2338 5294 2341
rect 162 2328 534 2331
rect 634 2328 718 2331
rect 738 2328 758 2331
rect 762 2328 902 2331
rect 954 2328 958 2331
rect 1010 2328 1102 2331
rect 1106 2328 1182 2331
rect 1194 2328 1742 2331
rect 1874 2328 1878 2331
rect 1890 2328 1894 2331
rect 1906 2328 2006 2331
rect 2050 2328 2182 2331
rect 2194 2328 2214 2331
rect 2222 2331 2225 2338
rect 2222 2328 2366 2331
rect 2402 2328 2646 2331
rect 2874 2328 2918 2331
rect 3058 2328 3150 2331
rect 3162 2328 3182 2331
rect 3250 2328 3294 2331
rect 3314 2328 3382 2331
rect 3386 2328 3470 2331
rect 3682 2328 3761 2331
rect 3882 2328 3886 2331
rect 4058 2328 4078 2331
rect 4082 2328 4126 2331
rect 4274 2328 4470 2331
rect 4474 2328 4510 2331
rect 4554 2328 4574 2331
rect 4682 2328 4697 2331
rect 4746 2328 4790 2331
rect 4794 2328 4934 2331
rect 4938 2328 4942 2331
rect 5194 2328 5222 2331
rect 5226 2328 5302 2331
rect 146 2318 369 2321
rect 378 2318 406 2321
rect 458 2318 510 2321
rect 514 2318 518 2321
rect 530 2318 614 2321
rect 618 2318 678 2321
rect 930 2318 1046 2321
rect 1394 2318 1518 2321
rect 1562 2318 1798 2321
rect 1862 2321 1865 2328
rect 2030 2322 2033 2328
rect 3758 2322 3761 2328
rect 1862 2318 1902 2321
rect 1930 2318 1942 2321
rect 2042 2318 2062 2321
rect 2218 2318 2254 2321
rect 3074 2318 3118 2321
rect 3122 2318 3206 2321
rect 3218 2318 3382 2321
rect 3386 2318 3510 2321
rect 3602 2318 3614 2321
rect 3766 2318 3774 2321
rect 3778 2318 3958 2321
rect 4466 2318 4502 2321
rect 4506 2318 4518 2321
rect 4530 2318 4686 2321
rect 4694 2321 4697 2328
rect 4694 2318 4838 2321
rect 5162 2318 5166 2321
rect 58 2308 174 2311
rect 178 2308 190 2311
rect 210 2308 254 2311
rect 366 2311 369 2318
rect 366 2308 590 2311
rect 594 2308 694 2311
rect 718 2308 806 2311
rect 810 2308 846 2311
rect 994 2308 1030 2311
rect 1034 2308 1150 2311
rect 1282 2308 1526 2311
rect 1578 2308 1630 2311
rect 1714 2308 1734 2311
rect 1906 2308 1934 2311
rect 1938 2308 1966 2311
rect 2018 2308 2214 2311
rect 2242 2308 2534 2311
rect 2538 2308 2894 2311
rect 3010 2308 3142 2311
rect 3530 2308 3678 2311
rect 3730 2308 3750 2311
rect 3778 2308 3910 2311
rect 4042 2308 4198 2311
rect 4546 2308 4614 2311
rect 5066 2308 5134 2311
rect 5138 2308 5174 2311
rect 186 2298 214 2301
rect 234 2298 246 2301
rect 718 2301 721 2308
rect 856 2303 858 2307
rect 862 2303 865 2307
rect 870 2303 872 2307
rect 1872 2303 1874 2307
rect 1878 2303 1881 2307
rect 1886 2303 1888 2307
rect 2904 2303 2906 2307
rect 2910 2303 2913 2307
rect 2918 2303 2920 2307
rect 3928 2303 3930 2307
rect 3934 2303 3937 2307
rect 3942 2303 3944 2307
rect 4952 2303 4954 2307
rect 4958 2303 4961 2307
rect 4966 2303 4968 2307
rect 274 2298 721 2301
rect 786 2298 790 2301
rect 1346 2298 1390 2301
rect 1482 2298 1494 2301
rect 1506 2298 1518 2301
rect 1626 2298 1726 2301
rect 1738 2298 1742 2301
rect 1954 2298 1966 2301
rect 2378 2298 2758 2301
rect 3082 2298 3550 2301
rect 3642 2298 3878 2301
rect 4594 2298 4894 2301
rect 4994 2298 5086 2301
rect 5130 2298 5166 2301
rect 66 2288 110 2291
rect 114 2288 118 2291
rect 214 2291 217 2298
rect 2846 2292 2849 2298
rect 214 2288 262 2291
rect 266 2288 286 2291
rect 290 2288 526 2291
rect 666 2288 806 2291
rect 1034 2288 1038 2291
rect 1130 2288 1134 2291
rect 1258 2288 1598 2291
rect 1610 2288 1854 2291
rect 1866 2288 1878 2291
rect 1882 2288 1958 2291
rect 2058 2288 2174 2291
rect 2178 2288 2198 2291
rect 2202 2288 2454 2291
rect 2890 2288 3006 2291
rect 3090 2288 3142 2291
rect 3146 2288 3222 2291
rect 3226 2288 3366 2291
rect 3538 2288 3558 2291
rect 3746 2288 3766 2291
rect 3770 2288 3774 2291
rect 3858 2288 3878 2291
rect 3882 2288 3889 2291
rect 3930 2288 3966 2291
rect 3970 2288 4022 2291
rect 4314 2288 4334 2291
rect 4354 2288 4366 2291
rect 4370 2288 4526 2291
rect 4566 2288 4574 2291
rect 4578 2288 4630 2291
rect 4642 2288 4694 2291
rect 4778 2288 5025 2291
rect 5050 2288 5110 2291
rect 186 2278 190 2281
rect 218 2278 270 2281
rect 274 2278 310 2281
rect 386 2278 398 2281
rect 1138 2278 1246 2281
rect 1594 2278 1598 2281
rect 1834 2278 1894 2281
rect 2098 2278 2110 2281
rect 2250 2278 2366 2281
rect 2370 2278 2374 2281
rect 2466 2278 2686 2281
rect 2886 2281 2889 2288
rect 5022 2282 5025 2288
rect 5150 2282 5153 2288
rect 2886 2278 2918 2281
rect 2978 2278 3070 2281
rect 3170 2278 3422 2281
rect 3426 2278 3478 2281
rect 3594 2278 3670 2281
rect 3674 2278 3734 2281
rect 3762 2278 3886 2281
rect 3890 2278 3894 2281
rect 3898 2278 3918 2281
rect 3946 2278 3990 2281
rect 4082 2278 4134 2281
rect 4330 2278 4342 2281
rect 4402 2278 4470 2281
rect 4474 2278 4550 2281
rect 4554 2278 4654 2281
rect 4682 2278 4686 2281
rect 4738 2278 4742 2281
rect 4762 2278 4854 2281
rect 4858 2278 4910 2281
rect 4914 2278 4982 2281
rect 5206 2281 5209 2288
rect 5154 2278 5246 2281
rect 5250 2278 5278 2281
rect 5306 2278 5310 2281
rect 106 2268 158 2271
rect 382 2271 385 2278
rect 346 2268 385 2271
rect 410 2268 422 2271
rect 474 2268 478 2271
rect 546 2268 558 2271
rect 654 2271 657 2278
rect 602 2268 657 2271
rect 926 2271 929 2278
rect 802 2268 929 2271
rect 1118 2271 1121 2278
rect 1118 2268 1166 2271
rect 1286 2271 1289 2278
rect 1286 2268 1350 2271
rect 1530 2268 1542 2271
rect 1546 2268 1558 2271
rect 1570 2268 1598 2271
rect 1718 2271 1721 2278
rect 3582 2272 3585 2278
rect 1718 2268 1750 2271
rect 1874 2268 1878 2271
rect 2066 2268 2094 2271
rect 2098 2268 2102 2271
rect 2282 2268 2286 2271
rect 2290 2268 2350 2271
rect 2354 2268 2358 2271
rect 2370 2268 2494 2271
rect 2498 2268 2510 2271
rect 2698 2268 2790 2271
rect 2906 2268 3062 2271
rect 3106 2268 3134 2271
rect 3282 2268 3294 2271
rect 3378 2268 3390 2271
rect 3662 2268 3790 2271
rect 3906 2268 3934 2271
rect 3986 2268 4014 2271
rect 4018 2268 4025 2271
rect 4034 2268 4102 2271
rect 4114 2268 4158 2271
rect 4166 2271 4169 2278
rect 4166 2268 4321 2271
rect 4338 2268 4374 2271
rect 4386 2268 4430 2271
rect 4490 2268 4534 2271
rect 4674 2268 4734 2271
rect 4738 2268 4766 2271
rect 4902 2268 4942 2271
rect 4970 2268 5062 2271
rect 5138 2268 5153 2271
rect 5178 2268 5222 2271
rect 54 2262 57 2268
rect 238 2262 241 2268
rect 1510 2262 1513 2268
rect 322 2258 406 2261
rect 426 2258 430 2261
rect 458 2258 550 2261
rect 594 2258 710 2261
rect 714 2258 958 2261
rect 1290 2258 1342 2261
rect 1346 2258 1382 2261
rect 1402 2258 1430 2261
rect 1566 2261 1569 2268
rect 1942 2262 1945 2268
rect 2638 2262 2641 2268
rect 3662 2262 3665 2268
rect 1554 2258 1569 2261
rect 1702 2258 1710 2261
rect 1794 2258 1878 2261
rect 1978 2258 1990 2261
rect 2074 2258 2102 2261
rect 2194 2258 2222 2261
rect 2226 2258 2233 2261
rect 2250 2258 2254 2261
rect 2298 2258 2302 2261
rect 2802 2258 2806 2261
rect 2962 2258 2966 2261
rect 2986 2258 3102 2261
rect 3138 2258 3142 2261
rect 3482 2258 3502 2261
rect 3718 2258 3766 2261
rect 3850 2258 3854 2261
rect 4022 2261 4025 2268
rect 4110 2262 4113 2268
rect 4022 2258 4054 2261
rect 4098 2258 4102 2261
rect 4138 2258 4150 2261
rect 4226 2258 4302 2261
rect 4306 2258 4310 2261
rect 4318 2261 4321 2268
rect 4798 2262 4801 2268
rect 4902 2262 4905 2268
rect 5150 2262 5153 2268
rect 4318 2258 4406 2261
rect 4426 2258 4502 2261
rect 4506 2258 4566 2261
rect 4578 2258 4638 2261
rect 4722 2258 4726 2261
rect 4850 2258 4889 2261
rect 4914 2258 4926 2261
rect 4930 2258 4937 2261
rect 5002 2258 5006 2261
rect 5154 2258 5214 2261
rect 5218 2258 5278 2261
rect 110 2252 113 2258
rect 174 2252 177 2258
rect 190 2251 193 2258
rect 1102 2252 1105 2258
rect 1198 2252 1201 2258
rect 190 2248 206 2251
rect 410 2248 422 2251
rect 650 2248 758 2251
rect 1034 2248 1038 2251
rect 1590 2251 1593 2258
rect 1702 2252 1705 2258
rect 3718 2252 3721 2258
rect 4014 2252 4017 2258
rect 4886 2252 4889 2258
rect 1570 2248 1593 2251
rect 1770 2248 2022 2251
rect 2058 2248 2134 2251
rect 2154 2248 2174 2251
rect 2226 2248 2262 2251
rect 2410 2248 2430 2251
rect 2682 2248 2710 2251
rect 2714 2248 2798 2251
rect 3018 2248 3286 2251
rect 3330 2248 3366 2251
rect 3370 2248 3566 2251
rect 3786 2248 3806 2251
rect 3810 2248 3942 2251
rect 4058 2248 4222 2251
rect 4274 2248 4414 2251
rect 4418 2248 4574 2251
rect 4594 2248 4750 2251
rect 5002 2248 5006 2251
rect 5010 2248 5086 2251
rect 5242 2248 5246 2251
rect 1638 2242 1641 2248
rect 370 2238 414 2241
rect 554 2238 678 2241
rect 954 2238 1014 2241
rect 1018 2238 1334 2241
rect 1410 2238 1470 2241
rect 1650 2238 1718 2241
rect 1738 2238 1766 2241
rect 1922 2238 2126 2241
rect 2186 2238 2254 2241
rect 2258 2238 2318 2241
rect 2522 2238 2854 2241
rect 2970 2238 3382 2241
rect 3794 2238 3814 2241
rect 3818 2238 3857 2241
rect 3906 2238 3926 2241
rect 4218 2238 4286 2241
rect 4290 2238 4294 2241
rect 4314 2238 4382 2241
rect 4394 2238 4446 2241
rect 4450 2238 4606 2241
rect 4610 2238 4774 2241
rect 5034 2238 5062 2241
rect 5066 2238 5206 2241
rect 330 2228 534 2231
rect 538 2228 798 2231
rect 858 2228 1638 2231
rect 1954 2228 1974 2231
rect 1978 2228 2358 2231
rect 2750 2228 3334 2231
rect 3338 2228 3622 2231
rect 3698 2228 3846 2231
rect 3854 2231 3857 2238
rect 3854 2228 4022 2231
rect 4066 2228 4278 2231
rect 4294 2228 4390 2231
rect 4402 2228 4526 2231
rect 4530 2228 4558 2231
rect 4602 2228 4622 2231
rect 2750 2222 2753 2228
rect 4294 2222 4297 2228
rect 370 2218 486 2221
rect 490 2218 542 2221
rect 546 2218 990 2221
rect 994 2218 1062 2221
rect 1186 2218 1438 2221
rect 1530 2218 1838 2221
rect 1842 2218 2222 2221
rect 2230 2218 2502 2221
rect 2906 2218 2985 2221
rect 3178 2218 3190 2221
rect 3402 2218 3478 2221
rect 3482 2218 3694 2221
rect 3874 2218 3910 2221
rect 4034 2218 4049 2221
rect 4162 2218 4190 2221
rect 4306 2218 4430 2221
rect 5262 2221 5265 2228
rect 5186 2218 5265 2221
rect 378 2208 566 2211
rect 1402 2208 1542 2211
rect 1546 2208 1630 2211
rect 1642 2208 2078 2211
rect 2130 2208 2134 2211
rect 2146 2208 2174 2211
rect 2230 2211 2233 2218
rect 2194 2208 2233 2211
rect 2578 2208 2974 2211
rect 2982 2211 2985 2218
rect 2982 2208 3246 2211
rect 3498 2208 3742 2211
rect 3746 2208 4038 2211
rect 4046 2211 4049 2218
rect 4046 2208 4270 2211
rect 4994 2208 5222 2211
rect 5266 2208 5278 2211
rect 344 2203 346 2207
rect 350 2203 353 2207
rect 358 2203 360 2207
rect 1368 2203 1370 2207
rect 1374 2203 1377 2207
rect 1382 2203 1384 2207
rect 10 2198 14 2201
rect 1466 2198 1990 2201
rect 2074 2198 2078 2201
rect 2090 2198 2150 2201
rect 2190 2201 2193 2208
rect 2392 2203 2394 2207
rect 2398 2203 2401 2207
rect 2406 2203 2408 2207
rect 3416 2203 3418 2207
rect 3422 2203 3425 2207
rect 3430 2203 3432 2207
rect 4440 2203 4442 2207
rect 4446 2203 4449 2207
rect 4454 2203 4456 2207
rect 2162 2198 2193 2201
rect 2226 2198 2382 2201
rect 2594 2198 2822 2201
rect 2826 2198 2862 2201
rect 2874 2198 2942 2201
rect 3146 2198 3366 2201
rect 3370 2198 3406 2201
rect 3618 2198 3630 2201
rect 3722 2198 3998 2201
rect 4258 2198 4422 2201
rect 4738 2198 4958 2201
rect 5146 2198 5206 2201
rect 1414 2192 1417 2198
rect 778 2188 1182 2191
rect 1426 2188 1569 2191
rect 1634 2188 1830 2191
rect 1850 2188 2142 2191
rect 2274 2188 4062 2191
rect 4154 2188 4294 2191
rect 4642 2188 4726 2191
rect 4866 2188 4934 2191
rect 4938 2188 5150 2191
rect 5158 2188 5281 2191
rect 162 2178 166 2181
rect 486 2181 489 2188
rect 466 2178 534 2181
rect 642 2178 694 2181
rect 766 2181 769 2188
rect 1566 2182 1569 2188
rect 698 2178 769 2181
rect 930 2178 950 2181
rect 1474 2178 1478 2181
rect 1642 2178 1654 2181
rect 1810 2178 1958 2181
rect 2106 2178 2254 2181
rect 2858 2178 2886 2181
rect 3050 2178 3534 2181
rect 3994 2178 4065 2181
rect 4222 2178 4230 2181
rect 4234 2178 4262 2181
rect 4658 2178 4678 2181
rect 4794 2178 4870 2181
rect 5158 2181 5161 2188
rect 5278 2182 5281 2188
rect 5122 2178 5161 2181
rect 5194 2178 5214 2181
rect 130 2168 158 2171
rect 162 2168 166 2171
rect 282 2168 414 2171
rect 418 2168 662 2171
rect 682 2168 686 2171
rect 1542 2171 1545 2178
rect 4062 2172 4065 2178
rect 1542 2168 1614 2171
rect 1658 2168 1670 2171
rect 1674 2168 1702 2171
rect 1866 2168 1934 2171
rect 1938 2168 1958 2171
rect 1994 2168 2118 2171
rect 2146 2168 2478 2171
rect 2482 2168 3438 2171
rect 3570 2168 3670 2171
rect 3850 2168 3990 2171
rect 4066 2168 4094 2171
rect 4098 2168 4238 2171
rect 4278 2171 4281 2178
rect 4258 2168 4310 2171
rect 4346 2168 4502 2171
rect 4506 2168 4550 2171
rect 4554 2168 4598 2171
rect 4634 2168 4665 2171
rect 58 2158 62 2161
rect 158 2158 174 2161
rect 178 2158 214 2161
rect 402 2158 454 2161
rect 482 2158 622 2161
rect 626 2158 662 2161
rect 742 2161 745 2168
rect 4662 2162 4665 2168
rect 4950 2171 4953 2178
rect 4950 2168 4982 2171
rect 5082 2168 5094 2171
rect 5202 2168 5254 2171
rect 666 2158 745 2161
rect 1162 2158 1286 2161
rect 1338 2158 1542 2161
rect 1626 2158 1654 2161
rect 1746 2158 2054 2161
rect 2362 2158 2438 2161
rect 2458 2158 2470 2161
rect 2562 2158 2582 2161
rect 2586 2158 2614 2161
rect 2762 2158 2846 2161
rect 2874 2158 2894 2161
rect 2994 2158 3070 2161
rect 3074 2158 3190 2161
rect 3194 2158 3198 2161
rect 3218 2158 3230 2161
rect 3258 2158 3574 2161
rect 3914 2158 3926 2161
rect 3982 2158 4022 2161
rect 4106 2158 4214 2161
rect 4218 2158 4222 2161
rect 4306 2158 4334 2161
rect 4570 2158 4590 2161
rect 4738 2158 4766 2161
rect 4830 2161 4833 2168
rect 4770 2158 4833 2161
rect 4906 2158 4926 2161
rect 5026 2158 5030 2161
rect 5102 2161 5105 2168
rect 5038 2158 5105 2161
rect 5198 2162 5201 2168
rect 5274 2158 5289 2161
rect 158 2152 161 2158
rect 782 2152 785 2158
rect 114 2148 134 2151
rect 210 2148 390 2151
rect 426 2148 446 2151
rect 522 2148 558 2151
rect 562 2148 606 2151
rect 610 2148 622 2151
rect 650 2148 702 2151
rect 762 2148 774 2151
rect 834 2148 894 2151
rect 898 2148 934 2151
rect 1062 2151 1065 2158
rect 1542 2152 1545 2158
rect 1062 2148 1190 2151
rect 1250 2148 1254 2151
rect 1362 2148 1390 2151
rect 1490 2148 1494 2151
rect 1562 2148 1590 2151
rect 1650 2148 1678 2151
rect 1686 2151 1689 2158
rect 1686 2148 1710 2151
rect 1714 2148 1726 2151
rect 1746 2148 2014 2151
rect 82 2138 102 2141
rect 106 2138 142 2141
rect 242 2138 286 2141
rect 354 2138 382 2141
rect 546 2138 582 2141
rect 586 2138 598 2141
rect 602 2138 806 2141
rect 834 2138 854 2141
rect 858 2138 910 2141
rect 930 2138 942 2141
rect 1078 2138 1150 2141
rect 1154 2138 1222 2141
rect 1422 2141 1425 2148
rect 1502 2142 1505 2148
rect 2082 2148 2121 2151
rect 2130 2148 2150 2151
rect 2182 2151 2185 2158
rect 2154 2148 2185 2151
rect 2190 2148 2270 2151
rect 2326 2151 2329 2158
rect 3982 2152 3985 2158
rect 2306 2148 2329 2151
rect 2418 2148 2462 2151
rect 2490 2148 2646 2151
rect 2698 2148 2718 2151
rect 2722 2148 2814 2151
rect 2818 2148 2822 2151
rect 2834 2148 2894 2151
rect 2930 2148 3030 2151
rect 3050 2148 3062 2151
rect 3082 2148 3134 2151
rect 3146 2148 3214 2151
rect 3234 2148 3262 2151
rect 3274 2148 3278 2151
rect 3282 2148 3302 2151
rect 3322 2148 3326 2151
rect 3394 2148 3406 2151
rect 3602 2148 3606 2151
rect 3682 2148 3798 2151
rect 3834 2148 3902 2151
rect 3914 2148 3982 2151
rect 4250 2148 4278 2151
rect 4282 2148 4294 2151
rect 4418 2148 4438 2151
rect 4442 2148 4526 2151
rect 4554 2148 4582 2151
rect 4602 2148 4718 2151
rect 4762 2148 4790 2151
rect 5038 2151 5041 2158
rect 5286 2152 5289 2158
rect 5302 2152 5305 2158
rect 4970 2148 5041 2151
rect 5066 2148 5198 2151
rect 5202 2148 5230 2151
rect 5250 2148 5254 2151
rect 2118 2142 2121 2148
rect 1362 2138 1502 2141
rect 1618 2138 1638 2141
rect 1642 2138 1654 2141
rect 1706 2138 1718 2141
rect 1898 2138 1942 2141
rect 2190 2141 2193 2148
rect 2146 2138 2193 2141
rect 2286 2141 2289 2148
rect 2646 2142 2649 2148
rect 3118 2142 3121 2148
rect 2210 2138 2414 2141
rect 2434 2138 2446 2141
rect 2450 2138 2630 2141
rect 2778 2138 2934 2141
rect 2938 2138 2977 2141
rect 1078 2132 1081 2138
rect 58 2128 70 2131
rect 82 2128 94 2131
rect 98 2128 105 2131
rect 114 2128 206 2131
rect 210 2128 262 2131
rect 346 2128 366 2131
rect 442 2128 566 2131
rect 666 2128 854 2131
rect 1090 2128 1094 2131
rect 1490 2128 1502 2131
rect 1574 2131 1577 2138
rect 1574 2128 1670 2131
rect 1754 2128 1761 2131
rect 2006 2131 2009 2138
rect 1882 2128 2009 2131
rect 2086 2131 2089 2138
rect 2974 2132 2977 2138
rect 3058 2138 3094 2141
rect 3098 2138 3102 2141
rect 3122 2138 3158 2141
rect 3242 2138 3270 2141
rect 3274 2138 3286 2141
rect 3334 2141 3337 2148
rect 5062 2142 5065 2148
rect 3298 2138 3337 2141
rect 3754 2138 3846 2141
rect 3914 2138 4606 2141
rect 4618 2138 4646 2141
rect 4690 2138 4822 2141
rect 4826 2138 4846 2141
rect 4850 2138 4926 2141
rect 4954 2138 4958 2141
rect 5066 2138 5078 2141
rect 5218 2138 5246 2141
rect 5306 2138 5310 2141
rect 2982 2132 2985 2138
rect 2086 2128 2126 2131
rect 2146 2128 2158 2131
rect 2166 2128 2214 2131
rect 2266 2128 2270 2131
rect 2330 2128 2502 2131
rect 2522 2128 2750 2131
rect 2802 2128 2926 2131
rect 3074 2128 3142 2131
rect 3826 2128 3830 2131
rect 3858 2128 4006 2131
rect 4026 2128 4030 2131
rect 4082 2128 4094 2131
rect 4098 2128 4206 2131
rect 4442 2128 4470 2131
rect 4474 2128 4558 2131
rect 4610 2128 4697 2131
rect 102 2122 105 2128
rect 1758 2122 1761 2128
rect 354 2118 606 2121
rect 626 2118 782 2121
rect 994 2118 998 2121
rect 1090 2118 1334 2121
rect 1490 2118 1662 2121
rect 1666 2118 1694 2121
rect 1862 2118 1998 2121
rect 2166 2121 2169 2128
rect 2066 2118 2169 2121
rect 2178 2118 2270 2121
rect 2290 2118 2294 2121
rect 2402 2118 2718 2121
rect 2730 2118 2814 2121
rect 2818 2118 3454 2121
rect 3838 2121 3841 2128
rect 4694 2122 4697 2128
rect 4702 2128 4742 2131
rect 4906 2128 5014 2131
rect 5106 2128 5158 2131
rect 5186 2128 5230 2131
rect 5234 2128 5246 2131
rect 5298 2128 5302 2131
rect 5314 2128 5358 2131
rect 4702 2122 4705 2128
rect 3466 2118 3841 2121
rect 4042 2118 4054 2121
rect 4354 2118 4414 2121
rect 4418 2118 4542 2121
rect 4546 2118 4622 2121
rect 4754 2118 4902 2121
rect 5034 2118 5078 2121
rect 110 2112 113 2118
rect 26 2108 46 2111
rect 274 2108 318 2111
rect 322 2108 406 2111
rect 418 2108 494 2111
rect 1050 2108 1214 2111
rect 1474 2108 1606 2111
rect 1634 2108 1646 2111
rect 1862 2111 1865 2118
rect 1650 2108 1865 2111
rect 1906 2108 1998 2111
rect 2050 2108 2094 2111
rect 2098 2108 2622 2111
rect 2650 2108 2678 2111
rect 2726 2111 2729 2118
rect 4142 2112 4145 2118
rect 2682 2108 2729 2111
rect 3082 2108 3486 2111
rect 3514 2108 3870 2111
rect 4162 2108 4310 2111
rect 4314 2108 4342 2111
rect 4346 2108 4478 2111
rect 4482 2108 4486 2111
rect 4522 2108 4526 2111
rect 5002 2108 5110 2111
rect 856 2103 858 2107
rect 862 2103 865 2107
rect 870 2103 872 2107
rect 1872 2103 1874 2107
rect 1878 2103 1881 2107
rect 1886 2103 1888 2107
rect 2904 2103 2906 2107
rect 2910 2103 2913 2107
rect 2918 2103 2920 2107
rect 3928 2103 3930 2107
rect 3934 2103 3937 2107
rect 3942 2103 3944 2107
rect 4952 2103 4954 2107
rect 4958 2103 4961 2107
rect 4966 2103 4968 2107
rect 34 2098 134 2101
rect 178 2098 438 2101
rect 1050 2098 1086 2101
rect 1498 2098 1542 2101
rect 1658 2098 1814 2101
rect 2194 2098 2534 2101
rect 2706 2098 2726 2101
rect 3178 2098 3326 2101
rect 3354 2098 3414 2101
rect 3418 2098 3502 2101
rect 4010 2098 4070 2101
rect 4338 2098 4790 2101
rect 5066 2098 5086 2101
rect 234 2088 254 2091
rect 402 2088 422 2091
rect 430 2088 454 2091
rect 478 2091 481 2098
rect 478 2088 486 2091
rect 586 2088 1270 2091
rect 1418 2088 1478 2091
rect 1482 2088 1534 2091
rect 1570 2088 1582 2091
rect 1914 2088 1926 2091
rect 1930 2088 2166 2091
rect 2266 2088 2302 2091
rect 2370 2088 2542 2091
rect 2874 2088 3054 2091
rect 3066 2088 3654 2091
rect 3714 2088 3721 2091
rect 3730 2088 4022 2091
rect 4658 2088 4686 2091
rect 4694 2088 4854 2091
rect 4962 2088 4982 2091
rect 5282 2088 5302 2091
rect 430 2082 433 2088
rect 90 2078 142 2081
rect 178 2078 206 2081
rect 210 2078 246 2081
rect 442 2078 566 2081
rect 586 2078 646 2081
rect 650 2078 806 2081
rect 810 2078 1022 2081
rect 1034 2078 1054 2081
rect 1522 2078 1558 2081
rect 1562 2078 1569 2081
rect 1594 2078 1742 2081
rect 1758 2078 1774 2081
rect 1778 2078 1782 2081
rect 2010 2078 2078 2081
rect 2298 2078 2318 2081
rect 2378 2078 2401 2081
rect 2426 2078 2454 2081
rect 2458 2078 2502 2081
rect 2506 2078 2574 2081
rect 2858 2078 2870 2081
rect 2930 2078 3006 2081
rect 3050 2078 3102 2081
rect 3106 2078 3134 2081
rect 3202 2078 3254 2081
rect 3362 2078 3406 2081
rect 3426 2078 3566 2081
rect 3570 2078 3622 2081
rect 3750 2078 3758 2081
rect 3762 2078 3822 2081
rect 4066 2078 4102 2081
rect 4178 2078 4198 2081
rect 4378 2078 4422 2081
rect 4426 2078 4550 2081
rect 4694 2081 4697 2088
rect 4602 2078 4697 2081
rect 4890 2078 5046 2081
rect 5098 2078 5174 2081
rect 66 2068 158 2071
rect 266 2068 270 2071
rect 314 2068 582 2071
rect 954 2068 1014 2071
rect 1070 2071 1073 2078
rect 1018 2068 1073 2071
rect 1262 2071 1265 2078
rect 1758 2072 1761 2078
rect 1262 2068 1310 2071
rect 1346 2068 1414 2071
rect 1418 2068 1441 2071
rect 1570 2068 1582 2071
rect 1770 2068 1846 2071
rect 1930 2068 1934 2071
rect 2050 2068 2094 2071
rect 2198 2068 2206 2071
rect 2298 2068 2302 2071
rect 2326 2071 2329 2078
rect 2326 2068 2390 2071
rect 2398 2071 2401 2078
rect 3630 2072 3633 2078
rect 2398 2068 2542 2071
rect 2578 2068 2742 2071
rect 2778 2068 2790 2071
rect 3082 2068 3094 2071
rect 3162 2068 3222 2071
rect 3234 2068 3318 2071
rect 3354 2068 3366 2071
rect 3394 2068 3430 2071
rect 3490 2068 3494 2071
rect 3506 2068 3577 2071
rect 3802 2068 3966 2071
rect 3970 2068 3993 2071
rect 4058 2068 4062 2071
rect 4234 2068 4270 2071
rect 4490 2068 4494 2071
rect 4542 2068 4550 2071
rect 4778 2068 4982 2071
rect 4994 2068 4998 2071
rect 5082 2068 5094 2071
rect 1334 2062 1337 2068
rect 1438 2062 1441 2068
rect 2118 2062 2121 2068
rect 2174 2062 2177 2068
rect 2198 2062 2201 2068
rect 154 2058 246 2061
rect 250 2058 270 2061
rect 274 2058 286 2061
rect 306 2058 414 2061
rect 458 2058 518 2061
rect 906 2058 958 2061
rect 962 2058 1022 2061
rect 1466 2058 1470 2061
rect 1562 2058 1566 2061
rect 1586 2058 2022 2061
rect 2026 2058 2070 2061
rect 2074 2058 2086 2061
rect 2338 2058 2446 2061
rect 2450 2058 2478 2061
rect 2566 2061 2569 2068
rect 2822 2062 2825 2068
rect 2830 2062 2833 2068
rect 2498 2058 2569 2061
rect 2666 2058 2678 2061
rect 2682 2058 2686 2061
rect 2690 2058 2702 2061
rect 2770 2058 2798 2061
rect 2982 2061 2985 2068
rect 3574 2062 3577 2068
rect 3990 2062 3993 2068
rect 4542 2062 4545 2068
rect 4718 2062 4721 2068
rect 4766 2062 4769 2068
rect 2978 2058 2985 2061
rect 3074 2058 3078 2061
rect 3106 2058 3134 2061
rect 3194 2058 3214 2061
rect 3290 2058 3294 2061
rect 3362 2058 3374 2061
rect 3442 2058 3550 2061
rect 3590 2058 3982 2061
rect 4122 2058 4142 2061
rect 4146 2058 4166 2061
rect 4242 2058 4246 2061
rect 4338 2058 4342 2061
rect 4770 2058 5246 2061
rect 1246 2052 1249 2058
rect 42 2048 78 2051
rect 218 2048 233 2051
rect 298 2048 318 2051
rect 418 2048 518 2051
rect 522 2048 574 2051
rect 1074 2048 1078 2051
rect 1082 2048 1182 2051
rect 1282 2048 1574 2051
rect 1658 2048 1662 2051
rect 1730 2048 1750 2051
rect 1778 2048 1798 2051
rect 1866 2048 1870 2051
rect 2066 2048 2094 2051
rect 2186 2048 2190 2051
rect 2322 2048 2326 2051
rect 2434 2048 2462 2051
rect 2494 2051 2497 2058
rect 3590 2052 3593 2058
rect 2466 2048 2497 2051
rect 2514 2048 2542 2051
rect 2546 2048 2574 2051
rect 2618 2048 2622 2051
rect 2634 2048 2670 2051
rect 2674 2048 2726 2051
rect 2730 2048 2766 2051
rect 2794 2048 2798 2051
rect 2818 2048 2838 2051
rect 2842 2048 2849 2051
rect 2858 2048 3134 2051
rect 3138 2048 3174 2051
rect 3178 2048 3182 2051
rect 3186 2048 3206 2051
rect 3226 2048 3294 2051
rect 3346 2048 3438 2051
rect 3442 2048 3470 2051
rect 3610 2048 3838 2051
rect 4094 2051 4097 2058
rect 4406 2052 4409 2058
rect 4094 2048 4134 2051
rect 4218 2048 4222 2051
rect 4690 2048 4774 2051
rect 4802 2048 5230 2051
rect 5258 2048 5310 2051
rect 230 2042 233 2048
rect 1726 2042 1729 2048
rect 114 2038 134 2041
rect 138 2038 158 2041
rect 218 2038 222 2041
rect 394 2038 422 2041
rect 746 2038 1118 2041
rect 1122 2038 1166 2041
rect 1482 2038 1622 2041
rect 1674 2038 1686 2041
rect 1822 2041 1825 2048
rect 2782 2042 2785 2048
rect 1818 2038 1825 2041
rect 1994 2038 2246 2041
rect 2250 2038 2478 2041
rect 2490 2038 2510 2041
rect 2650 2038 2686 2041
rect 2690 2038 2694 2041
rect 2846 2041 2849 2048
rect 2846 2038 2894 2041
rect 3110 2038 3182 2041
rect 3198 2038 3206 2041
rect 3210 2038 3214 2041
rect 3226 2038 3254 2041
rect 3298 2038 3366 2041
rect 3558 2041 3561 2048
rect 3558 2038 3734 2041
rect 3986 2038 4102 2041
rect 4258 2038 4278 2041
rect 4282 2038 4574 2041
rect 4826 2038 5198 2041
rect 5234 2038 5238 2041
rect 178 2028 238 2031
rect 470 2031 473 2038
rect 3110 2032 3113 2038
rect 274 2028 473 2031
rect 482 2028 694 2031
rect 698 2028 758 2031
rect 1154 2028 1534 2031
rect 1786 2028 1790 2031
rect 1794 2028 1838 2031
rect 1842 2028 2150 2031
rect 2530 2028 2670 2031
rect 3154 2028 3358 2031
rect 3370 2028 3406 2031
rect 3414 2031 3417 2038
rect 3414 2028 3454 2031
rect 3534 2031 3537 2038
rect 3534 2028 3686 2031
rect 4170 2028 4510 2031
rect 4634 2028 4830 2031
rect 5026 2028 5057 2031
rect 5146 2028 5174 2031
rect 426 2018 454 2021
rect 474 2018 494 2021
rect 1306 2018 1390 2021
rect 1718 2021 1721 2028
rect 1562 2018 1721 2021
rect 1738 2018 1806 2021
rect 2114 2018 2158 2021
rect 2162 2018 2230 2021
rect 2422 2021 2425 2028
rect 2338 2018 2425 2021
rect 2458 2018 2598 2021
rect 2694 2021 2697 2028
rect 2618 2018 2697 2021
rect 2946 2018 2950 2021
rect 3058 2018 3286 2021
rect 3314 2018 3462 2021
rect 3466 2018 3478 2021
rect 3482 2018 3542 2021
rect 3750 2021 3753 2028
rect 5054 2022 5057 2028
rect 3658 2018 3753 2021
rect 4122 2018 4398 2021
rect 5082 2018 5094 2021
rect 5098 2018 5118 2021
rect 5170 2018 5198 2021
rect 410 2008 526 2011
rect 922 2008 926 2011
rect 1570 2008 1734 2011
rect 1818 2008 1846 2011
rect 1898 2008 1918 2011
rect 1930 2008 2142 2011
rect 2562 2008 2630 2011
rect 2930 2008 3246 2011
rect 4802 2008 5014 2011
rect 5042 2008 5070 2011
rect 344 2003 346 2007
rect 350 2003 353 2007
rect 358 2003 360 2007
rect 1368 2003 1370 2007
rect 1374 2003 1377 2007
rect 1382 2003 1384 2007
rect 2392 2003 2394 2007
rect 2398 2003 2401 2007
rect 2406 2003 2408 2007
rect 3416 2003 3418 2007
rect 3422 2003 3425 2007
rect 3430 2003 3432 2007
rect 4440 2003 4442 2007
rect 4446 2003 4449 2007
rect 4454 2003 4456 2007
rect 402 1998 502 2001
rect 506 1998 574 2001
rect 1626 1998 1926 2001
rect 2034 1998 2046 2001
rect 2426 1998 2510 2001
rect 2530 1998 2606 2001
rect 2730 1998 2838 2001
rect 3082 1998 3102 2001
rect 3162 1998 3190 2001
rect 3442 1998 3750 2001
rect 3754 1998 4270 2001
rect 5010 1998 5166 2001
rect 210 1988 462 1991
rect 466 1988 494 1991
rect 506 1988 518 1991
rect 730 1988 1150 1991
rect 1298 1988 1350 1991
rect 1354 1988 1446 1991
rect 1570 1988 3606 1991
rect 3682 1988 4070 1991
rect 4434 1988 4886 1991
rect 4938 1988 4942 1991
rect 5130 1988 5166 1991
rect 90 1978 214 1981
rect 258 1978 294 1981
rect 946 1978 1206 1981
rect 1418 1978 1574 1981
rect 1690 1978 1718 1981
rect 1722 1978 1777 1981
rect 1842 1978 1950 1981
rect 2042 1978 2054 1981
rect 2058 1978 2270 1981
rect 2282 1978 2462 1981
rect 2466 1978 2614 1981
rect 2626 1978 3390 1981
rect 3394 1978 4150 1981
rect 4714 1978 5150 1981
rect 6 1971 9 1978
rect 30 1971 33 1978
rect 1774 1972 1777 1978
rect 6 1968 33 1971
rect 42 1968 134 1971
rect 234 1968 238 1971
rect 274 1968 398 1971
rect 874 1968 902 1971
rect 906 1968 934 1971
rect 994 1968 1054 1971
rect 1082 1968 1118 1971
rect 1122 1968 1150 1971
rect 1266 1968 1502 1971
rect 1706 1968 1742 1971
rect 1838 1968 2014 1971
rect 2018 1968 2134 1971
rect 2138 1968 2166 1971
rect 2234 1968 2254 1971
rect 2282 1968 2302 1971
rect 2314 1968 2358 1971
rect 2378 1968 2454 1971
rect 3322 1968 3534 1971
rect 3578 1968 3894 1971
rect 3898 1968 4022 1971
rect 4026 1968 4070 1971
rect 5250 1968 5262 1971
rect 58 1958 78 1961
rect 146 1958 302 1961
rect 322 1958 390 1961
rect 394 1958 438 1961
rect 446 1961 449 1968
rect 446 1958 470 1961
rect 530 1958 534 1961
rect 582 1961 585 1968
rect 638 1961 641 1968
rect 582 1958 641 1961
rect 826 1958 910 1961
rect 938 1958 942 1961
rect 946 1958 990 1961
rect 994 1958 1110 1961
rect 1290 1958 1318 1961
rect 1602 1958 1614 1961
rect 1618 1958 1630 1961
rect 1838 1961 1841 1968
rect 1666 1958 1841 1961
rect 1850 1958 1862 1961
rect 1866 1958 2062 1961
rect 2066 1958 2110 1961
rect 2138 1958 2142 1961
rect 2274 1958 2430 1961
rect 2450 1958 2470 1961
rect 2482 1958 3238 1961
rect 3258 1958 3310 1961
rect 3362 1958 3406 1961
rect 4010 1958 4038 1961
rect 4042 1958 4054 1961
rect 4078 1961 4081 1968
rect 4078 1958 4118 1961
rect 4838 1961 4841 1968
rect 4838 1958 5038 1961
rect 5042 1958 5054 1961
rect 5194 1958 5214 1961
rect 5218 1958 5238 1961
rect 58 1948 94 1951
rect 266 1948 326 1951
rect 354 1948 366 1951
rect 578 1948 590 1951
rect 786 1948 830 1951
rect 922 1948 1022 1951
rect 1042 1948 1062 1951
rect 1102 1948 1134 1951
rect 1138 1948 1166 1951
rect 1222 1951 1225 1958
rect 1254 1951 1257 1958
rect 1222 1948 1257 1951
rect 1290 1948 1310 1951
rect 1450 1948 1494 1951
rect 1514 1948 1550 1951
rect 1594 1948 1601 1951
rect 1738 1948 1742 1951
rect 1778 1948 1790 1951
rect 1946 1948 1982 1951
rect 2002 1948 2646 1951
rect 2778 1948 2782 1951
rect 2810 1948 2830 1951
rect 2842 1948 2886 1951
rect 2994 1948 2998 1951
rect 3146 1948 3198 1951
rect 3202 1948 3214 1951
rect 3262 1948 3366 1951
rect 3370 1948 3398 1951
rect 3502 1948 3510 1951
rect 3514 1948 3694 1951
rect 3742 1948 3750 1951
rect 3754 1948 3865 1951
rect 3902 1951 3905 1958
rect 3874 1948 3878 1951
rect 38 1942 41 1948
rect 42 1938 62 1941
rect 82 1938 206 1941
rect 290 1938 294 1941
rect 382 1941 385 1948
rect 1102 1942 1105 1948
rect 3022 1942 3025 1948
rect 338 1938 478 1941
rect 522 1938 590 1941
rect 642 1938 646 1941
rect 842 1938 886 1941
rect 890 1938 926 1941
rect 994 1938 1006 1941
rect 1050 1938 1086 1941
rect 1282 1938 1294 1941
rect 1322 1938 1334 1941
rect 1354 1938 1390 1941
rect 1506 1938 1526 1941
rect 1530 1938 1542 1941
rect 1546 1938 1590 1941
rect 1746 1938 1838 1941
rect 1914 1938 1934 1941
rect 2010 1938 2014 1941
rect 2034 1938 2070 1941
rect 2074 1938 2086 1941
rect 2098 1938 2102 1941
rect 2122 1938 2150 1941
rect 2154 1938 2198 1941
rect 2226 1938 2230 1941
rect 2298 1938 2374 1941
rect 2378 1938 2454 1941
rect 2534 1938 2550 1941
rect 2554 1938 2646 1941
rect 2818 1938 2854 1941
rect 2882 1938 3022 1941
rect 3118 1941 3121 1948
rect 3262 1942 3265 1948
rect 3118 1938 3174 1941
rect 3298 1938 3334 1941
rect 3354 1938 3358 1941
rect 3862 1941 3865 1948
rect 3902 1948 3934 1951
rect 3938 1948 3950 1951
rect 3974 1951 3977 1958
rect 3974 1948 4030 1951
rect 4034 1948 4062 1951
rect 4386 1948 4422 1951
rect 4426 1948 4510 1951
rect 4914 1948 5094 1951
rect 5186 1948 5262 1951
rect 4182 1942 4185 1948
rect 3862 1938 3977 1941
rect 4050 1938 4102 1941
rect 4418 1938 4438 1941
rect 4806 1941 4809 1948
rect 4714 1938 4809 1941
rect 5026 1938 5030 1941
rect 5034 1938 5065 1941
rect 5210 1938 5214 1941
rect 1390 1932 1393 1938
rect 1654 1932 1657 1938
rect 34 1928 46 1931
rect 74 1928 78 1931
rect 218 1928 262 1931
rect 430 1928 470 1931
rect 474 1928 510 1931
rect 554 1928 614 1931
rect 978 1928 1014 1931
rect 1162 1928 1286 1931
rect 1538 1928 1646 1931
rect 1826 1928 1902 1931
rect 2066 1928 2078 1931
rect 2138 1928 2174 1931
rect 2178 1928 2185 1931
rect 2238 1931 2241 1938
rect 2534 1932 2537 1938
rect 2854 1932 2857 1938
rect 2210 1928 2241 1931
rect 2258 1928 2278 1931
rect 2290 1928 2302 1931
rect 2322 1928 2462 1931
rect 2802 1928 2822 1931
rect 2946 1928 2998 1931
rect 3214 1931 3217 1938
rect 3534 1932 3537 1938
rect 3742 1932 3745 1938
rect 3974 1932 3977 1938
rect 3146 1928 3193 1931
rect 3214 1928 3278 1931
rect 4350 1931 4353 1938
rect 5062 1932 5065 1938
rect 4350 1928 4390 1931
rect 4738 1928 4742 1931
rect 430 1922 433 1928
rect 210 1918 222 1921
rect 226 1918 310 1921
rect 594 1918 598 1921
rect 602 1918 630 1921
rect 958 1921 961 1928
rect 2934 1922 2937 1928
rect 3086 1922 3089 1928
rect 3190 1922 3193 1928
rect 786 1918 961 1921
rect 1330 1918 1446 1921
rect 1578 1918 1694 1921
rect 1706 1918 1822 1921
rect 1906 1918 1926 1921
rect 2130 1918 2158 1921
rect 2162 1918 2214 1921
rect 2218 1918 2318 1921
rect 2322 1918 2374 1921
rect 2394 1918 2510 1921
rect 2618 1918 2622 1921
rect 2834 1918 2862 1921
rect 2870 1918 2934 1921
rect 2946 1918 2998 1921
rect 3194 1918 3230 1921
rect 3314 1918 3486 1921
rect 3514 1918 3566 1921
rect 3574 1918 3582 1921
rect 3590 1921 3593 1928
rect 3590 1918 3598 1921
rect 3602 1918 3630 1921
rect 3698 1918 3702 1921
rect 3714 1918 4094 1921
rect 4146 1918 4190 1921
rect 4490 1918 4518 1921
rect 4522 1918 4534 1921
rect 4538 1918 4574 1921
rect 4582 1918 4774 1921
rect 4942 1918 5110 1921
rect 2798 1912 2801 1918
rect 162 1908 222 1911
rect 258 1908 342 1911
rect 362 1908 662 1911
rect 914 1908 1430 1911
rect 1450 1908 1454 1911
rect 1602 1908 1710 1911
rect 1922 1908 1958 1911
rect 1962 1908 2158 1911
rect 2170 1908 2190 1911
rect 2194 1908 2342 1911
rect 2346 1908 2438 1911
rect 2642 1908 2734 1911
rect 2870 1911 2873 1918
rect 2810 1908 2873 1911
rect 2930 1908 2958 1911
rect 3218 1908 3398 1911
rect 3490 1908 3542 1911
rect 3746 1908 3790 1911
rect 4582 1911 4585 1918
rect 4242 1908 4585 1911
rect 4690 1908 4694 1911
rect 4942 1911 4945 1918
rect 4706 1908 4945 1911
rect 856 1903 858 1907
rect 862 1903 865 1907
rect 870 1903 872 1907
rect 1872 1903 1874 1907
rect 1878 1903 1881 1907
rect 1886 1903 1888 1907
rect 2904 1903 2906 1907
rect 2910 1903 2913 1907
rect 2918 1903 2920 1907
rect 3928 1903 3930 1907
rect 3934 1903 3937 1907
rect 3942 1903 3944 1907
rect 4952 1903 4954 1907
rect 4958 1903 4961 1907
rect 4966 1903 4968 1907
rect 18 1898 62 1901
rect 170 1898 198 1901
rect 202 1898 238 1901
rect 1106 1898 1294 1901
rect 1386 1898 1606 1901
rect 1618 1898 1718 1901
rect 2002 1898 2014 1901
rect 2018 1898 2086 1901
rect 2226 1898 2238 1901
rect 2242 1898 2270 1901
rect 2282 1898 2350 1901
rect 2370 1898 2470 1901
rect 2634 1898 2662 1901
rect 2666 1898 2694 1901
rect 2706 1898 2718 1901
rect 2730 1898 2766 1901
rect 2818 1898 2846 1901
rect 2962 1898 3294 1901
rect 3954 1898 3982 1901
rect 3986 1898 4142 1901
rect 4146 1898 4254 1901
rect 4346 1898 4422 1901
rect 4426 1898 4470 1901
rect 4602 1898 4630 1901
rect 242 1888 334 1891
rect 826 1888 838 1891
rect 842 1888 870 1891
rect 890 1888 918 1891
rect 986 1888 1270 1891
rect 1554 1888 1582 1891
rect 1618 1888 1622 1891
rect 1770 1888 1838 1891
rect 1842 1888 1934 1891
rect 1938 1888 1974 1891
rect 2090 1888 2102 1891
rect 2182 1891 2185 1898
rect 2182 1888 2190 1891
rect 2298 1888 2302 1891
rect 2434 1888 2438 1891
rect 2626 1888 2638 1891
rect 2642 1888 2758 1891
rect 2762 1888 3078 1891
rect 3110 1888 3118 1891
rect 3122 1888 3158 1891
rect 3330 1888 3350 1891
rect 3394 1888 3406 1891
rect 3410 1888 3478 1891
rect 3678 1888 3774 1891
rect 3850 1888 4190 1891
rect 4274 1888 4302 1891
rect 4362 1888 4366 1891
rect 4778 1888 4806 1891
rect 4922 1888 4974 1891
rect 5050 1888 5166 1891
rect 5170 1888 5238 1891
rect 226 1878 270 1881
rect 330 1878 342 1881
rect 346 1878 366 1881
rect 382 1881 385 1888
rect 382 1878 526 1881
rect 530 1878 558 1881
rect 778 1878 998 1881
rect 1058 1878 1318 1881
rect 1442 1878 1494 1881
rect 1498 1878 1710 1881
rect 2102 1878 2110 1881
rect 2114 1878 2150 1881
rect 2178 1878 2422 1881
rect 2426 1878 2566 1881
rect 2570 1878 2606 1881
rect 2610 1878 2694 1881
rect 2698 1878 2718 1881
rect 2722 1878 3174 1881
rect 3678 1881 3681 1888
rect 3254 1878 3681 1881
rect 3938 1878 4110 1881
rect 4186 1878 4198 1881
rect 4242 1878 4278 1881
rect 4282 1878 4398 1881
rect 4402 1878 4654 1881
rect 5082 1878 5150 1881
rect 5194 1878 5198 1881
rect 694 1872 697 1878
rect 3254 1872 3257 1878
rect 114 1868 118 1871
rect 298 1868 302 1871
rect 306 1868 358 1871
rect 434 1868 441 1871
rect 450 1868 462 1871
rect 654 1868 670 1871
rect 994 1868 1054 1871
rect 1142 1868 1158 1871
rect 1258 1868 1350 1871
rect 1358 1868 1598 1871
rect 1602 1868 1614 1871
rect 1626 1868 1681 1871
rect 1738 1868 1750 1871
rect 1834 1868 1942 1871
rect 1946 1868 1998 1871
rect 2050 1868 2062 1871
rect 2066 1868 2094 1871
rect 2218 1868 2230 1871
rect 2234 1870 2278 1871
rect 2234 1868 2270 1870
rect 90 1858 102 1861
rect 214 1861 217 1868
rect 254 1861 257 1868
rect 438 1862 441 1868
rect 654 1862 657 1868
rect 214 1858 257 1861
rect 266 1858 286 1861
rect 658 1858 726 1861
rect 918 1861 921 1868
rect 1142 1862 1145 1868
rect 890 1858 942 1861
rect 962 1858 1009 1861
rect 1026 1858 1038 1861
rect 1042 1858 1086 1861
rect 1150 1858 1305 1861
rect 1358 1861 1361 1868
rect 1678 1862 1681 1868
rect 2274 1868 2278 1870
rect 2290 1868 2294 1871
rect 2374 1868 2422 1871
rect 2626 1868 2654 1871
rect 2674 1870 2766 1871
rect 2674 1868 2702 1870
rect 2374 1862 2377 1868
rect 2706 1868 2766 1870
rect 2834 1868 2846 1871
rect 2874 1868 2910 1871
rect 2922 1868 2958 1871
rect 2994 1868 3110 1871
rect 3114 1868 3126 1871
rect 3162 1868 3190 1871
rect 3338 1868 3422 1871
rect 3686 1871 3689 1878
rect 4158 1872 4161 1878
rect 4894 1872 4897 1878
rect 5014 1872 5017 1878
rect 5022 1872 5025 1878
rect 3686 1868 3806 1871
rect 4194 1868 4254 1871
rect 4298 1868 4302 1871
rect 4314 1868 4358 1871
rect 4362 1868 4382 1871
rect 4562 1868 4590 1871
rect 4594 1868 4662 1871
rect 4682 1868 4697 1871
rect 4826 1868 4830 1871
rect 4914 1868 4945 1871
rect 5218 1868 5246 1871
rect 5250 1868 5254 1871
rect 5258 1868 5294 1871
rect 1314 1858 1361 1861
rect 1554 1858 1590 1861
rect 1746 1858 1766 1861
rect 1770 1858 1926 1861
rect 1954 1858 2046 1861
rect 2050 1858 2110 1861
rect 2146 1858 2166 1861
rect 2418 1858 2449 1861
rect 2506 1858 2521 1861
rect 2538 1858 2566 1861
rect 2570 1858 2574 1861
rect 2594 1858 2670 1861
rect 2738 1858 2774 1861
rect 2826 1858 2854 1861
rect 2870 1858 2894 1861
rect 2906 1858 2918 1861
rect 2938 1858 2966 1861
rect 3066 1858 3078 1861
rect 3218 1858 3342 1861
rect 3362 1858 3390 1861
rect 3566 1861 3569 1868
rect 3410 1858 3622 1861
rect 3706 1858 3718 1861
rect 3722 1858 3742 1861
rect 3806 1861 3809 1868
rect 4694 1862 4697 1868
rect 4942 1862 4945 1868
rect 5126 1862 5129 1868
rect 3806 1858 3854 1861
rect 4186 1858 4238 1861
rect 4266 1858 4326 1861
rect 4330 1858 4342 1861
rect 4354 1858 4358 1861
rect 4458 1858 4486 1861
rect 4490 1858 4494 1861
rect 4586 1858 4638 1861
rect 4802 1858 4838 1861
rect 5010 1858 5070 1861
rect 5202 1858 5206 1861
rect 5210 1858 5230 1861
rect 5234 1858 5262 1861
rect 66 1848 110 1851
rect 162 1848 209 1851
rect 326 1851 329 1858
rect 638 1852 641 1858
rect 282 1848 329 1851
rect 546 1848 550 1851
rect 954 1848 974 1851
rect 1006 1851 1009 1858
rect 1150 1852 1153 1858
rect 1302 1852 1305 1858
rect 2446 1852 2449 1858
rect 978 1848 1001 1851
rect 1006 1848 1022 1851
rect 1026 1848 1038 1851
rect 1042 1848 1049 1851
rect 1498 1848 1606 1851
rect 1674 1848 1678 1851
rect 1690 1848 1750 1851
rect 1930 1848 1998 1851
rect 2106 1848 2350 1851
rect 2370 1848 2382 1851
rect 2506 1848 2510 1851
rect 2518 1851 2521 1858
rect 2870 1852 2873 1858
rect 4886 1852 4889 1858
rect 2518 1848 2630 1851
rect 2754 1848 2774 1851
rect 2778 1848 2782 1851
rect 3106 1848 3110 1851
rect 3154 1848 3158 1851
rect 3202 1848 3206 1851
rect 3330 1848 3334 1851
rect 3338 1848 3366 1851
rect 3398 1848 3438 1851
rect 4050 1848 4534 1851
rect 4538 1848 4574 1851
rect 4602 1848 4606 1851
rect 4634 1848 4678 1851
rect 4682 1848 4710 1851
rect 4942 1851 4945 1858
rect 4942 1848 5134 1851
rect 5138 1848 5174 1851
rect 38 1842 41 1848
rect 206 1842 209 1848
rect 998 1842 1001 1848
rect 2646 1842 2649 1848
rect 3398 1842 3401 1848
rect 82 1838 94 1841
rect 178 1838 198 1841
rect 250 1838 350 1841
rect 354 1838 582 1841
rect 1274 1838 1310 1841
rect 1362 1838 1526 1841
rect 1586 1838 1670 1841
rect 1930 1838 1942 1841
rect 2002 1838 2014 1841
rect 2130 1838 2294 1841
rect 2298 1838 2302 1841
rect 2530 1838 2558 1841
rect 2570 1838 2646 1841
rect 2690 1838 2830 1841
rect 2834 1838 2878 1841
rect 2882 1838 3014 1841
rect 3722 1838 4054 1841
rect 4058 1838 4182 1841
rect 4218 1838 4230 1841
rect 4498 1838 4505 1841
rect 4578 1838 4606 1841
rect 4610 1838 4694 1841
rect 5182 1841 5185 1848
rect 5182 1838 5222 1841
rect 5262 1841 5265 1848
rect 5226 1838 5265 1841
rect 4502 1832 4505 1838
rect 186 1828 214 1831
rect 802 1828 1454 1831
rect 1474 1828 2638 1831
rect 2722 1828 2854 1831
rect 2858 1828 4014 1831
rect 4018 1828 4406 1831
rect 5162 1828 5206 1831
rect 154 1818 582 1821
rect 746 1818 790 1821
rect 794 1818 814 1821
rect 818 1818 1006 1821
rect 1514 1818 1598 1821
rect 1610 1818 1870 1821
rect 1898 1818 1934 1821
rect 2014 1818 2110 1821
rect 2118 1818 2126 1821
rect 2130 1818 2182 1821
rect 2186 1818 2270 1821
rect 2390 1818 2398 1821
rect 2402 1818 2430 1821
rect 2538 1818 2606 1821
rect 2610 1818 2638 1821
rect 2858 1818 2870 1821
rect 3026 1818 3134 1821
rect 3138 1818 3174 1821
rect 3194 1818 3870 1821
rect 4058 1818 4070 1821
rect 4258 1818 4950 1821
rect 2014 1812 2017 1818
rect 738 1808 798 1811
rect 1762 1808 2014 1811
rect 2026 1808 2094 1811
rect 2098 1808 2326 1811
rect 2474 1808 3270 1811
rect 3274 1808 3406 1811
rect 4066 1808 4246 1811
rect 5050 1808 5142 1811
rect 344 1803 346 1807
rect 350 1803 353 1807
rect 358 1803 360 1807
rect 1368 1803 1370 1807
rect 1374 1803 1377 1807
rect 1382 1803 1384 1807
rect 2392 1803 2394 1807
rect 2398 1803 2401 1807
rect 2406 1803 2408 1807
rect 3416 1803 3418 1807
rect 3422 1803 3425 1807
rect 3430 1803 3432 1807
rect 4440 1803 4442 1807
rect 4446 1803 4449 1807
rect 4454 1803 4456 1807
rect 706 1798 846 1801
rect 882 1798 1318 1801
rect 1658 1798 1686 1801
rect 1706 1798 1950 1801
rect 1954 1798 1966 1801
rect 2122 1798 2134 1801
rect 2146 1798 2198 1801
rect 4218 1798 4238 1801
rect 4242 1798 4278 1801
rect 4282 1798 4334 1801
rect 4338 1798 4382 1801
rect 4642 1798 4710 1801
rect 4722 1798 4910 1801
rect 90 1788 126 1791
rect 162 1788 334 1791
rect 762 1788 918 1791
rect 1722 1788 1814 1791
rect 1842 1788 2038 1791
rect 2042 1788 2494 1791
rect 2498 1788 3982 1791
rect 4106 1788 4198 1791
rect 4202 1788 4214 1791
rect 4218 1788 4742 1791
rect 18 1778 70 1781
rect 74 1778 174 1781
rect 178 1778 574 1781
rect 730 1778 742 1781
rect 746 1778 750 1781
rect 754 1778 894 1781
rect 922 1778 998 1781
rect 1002 1778 1078 1781
rect 1154 1778 1174 1781
rect 1178 1778 1542 1781
rect 1634 1778 1894 1781
rect 2018 1778 2078 1781
rect 2146 1778 3190 1781
rect 4354 1778 4478 1781
rect 4482 1778 4526 1781
rect 4666 1778 4694 1781
rect 4698 1778 4742 1781
rect 4754 1778 4878 1781
rect 5202 1778 5262 1781
rect 6 1771 9 1778
rect 6 1768 22 1771
rect 42 1768 94 1771
rect 98 1768 134 1771
rect 282 1768 294 1771
rect 298 1768 390 1771
rect 418 1768 462 1771
rect 554 1768 910 1771
rect 1146 1768 1150 1771
rect 1234 1768 1654 1771
rect 2034 1768 2158 1771
rect 2194 1768 2222 1771
rect 2234 1768 2321 1771
rect 2394 1768 2414 1771
rect 2434 1768 2438 1771
rect 2450 1768 2462 1771
rect 2466 1768 2537 1771
rect 2554 1768 2558 1771
rect 2994 1768 3030 1771
rect 3186 1768 3710 1771
rect 4190 1768 4262 1771
rect 4370 1768 4414 1771
rect 4418 1768 4486 1771
rect 4546 1768 4582 1771
rect 4770 1768 4862 1771
rect 4898 1768 4926 1771
rect 4930 1768 4942 1771
rect 5202 1768 5214 1771
rect 34 1758 94 1761
rect 290 1758 310 1761
rect 394 1758 398 1761
rect 402 1758 894 1761
rect 926 1761 929 1768
rect 906 1758 929 1761
rect 1038 1761 1041 1768
rect 1010 1758 1041 1761
rect 1242 1758 1430 1761
rect 1694 1761 1697 1768
rect 2318 1762 2321 1768
rect 1694 1758 1718 1761
rect 1746 1758 1774 1761
rect 1866 1758 1990 1761
rect 2154 1758 2166 1761
rect 2202 1758 2294 1761
rect 2298 1758 2310 1761
rect 2354 1758 2366 1761
rect 2370 1758 2518 1761
rect 2522 1758 2526 1761
rect 2534 1761 2537 1768
rect 2534 1758 2553 1761
rect 2582 1761 2585 1768
rect 4190 1762 4193 1768
rect 2570 1758 2585 1761
rect 2642 1758 2646 1761
rect 2650 1758 2654 1761
rect 2898 1758 2934 1761
rect 2938 1758 2942 1761
rect 2962 1758 2982 1761
rect 2986 1758 2990 1761
rect 3170 1758 3462 1761
rect 3762 1758 3790 1761
rect 4354 1758 4358 1761
rect 4370 1758 4438 1761
rect 4622 1761 4625 1768
rect 4546 1758 4625 1761
rect 4634 1758 4638 1761
rect 4702 1761 4705 1768
rect 4690 1758 4705 1761
rect 4754 1758 4814 1761
rect 4834 1758 4854 1761
rect 4858 1758 4894 1761
rect 4898 1758 4958 1761
rect 4962 1758 5014 1761
rect 5066 1758 5070 1761
rect 5274 1758 5294 1761
rect 90 1748 94 1751
rect 130 1748 142 1751
rect 498 1748 686 1751
rect 746 1748 766 1751
rect 778 1748 798 1751
rect 906 1748 950 1751
rect 1086 1751 1089 1758
rect 954 1748 1089 1751
rect 1182 1751 1185 1758
rect 1170 1748 1185 1751
rect 1214 1752 1217 1758
rect 1494 1752 1497 1758
rect 1426 1748 1465 1751
rect 1542 1751 1545 1758
rect 2550 1752 2553 1758
rect 1542 1748 1606 1751
rect 1682 1748 1702 1751
rect 1722 1748 1734 1751
rect 1738 1748 1854 1751
rect 1882 1748 1974 1751
rect 1994 1748 2014 1751
rect 2138 1748 2342 1751
rect 2354 1748 2422 1751
rect 2466 1748 2478 1751
rect 2506 1748 2542 1751
rect 2578 1748 2598 1751
rect 2674 1748 2729 1751
rect 2802 1748 2822 1751
rect 2866 1748 2878 1751
rect 2970 1748 3014 1751
rect 3018 1748 3046 1751
rect 3506 1748 3550 1751
rect 3554 1748 3569 1751
rect 3594 1748 3614 1751
rect 3618 1748 3718 1751
rect 3722 1748 3726 1751
rect 3730 1748 3750 1751
rect 3894 1751 3897 1758
rect 5214 1752 5217 1758
rect 5238 1752 5241 1758
rect 3866 1748 3897 1751
rect 4090 1748 4102 1751
rect 4186 1748 4198 1751
rect 4258 1748 4286 1751
rect 4290 1748 4310 1751
rect 4346 1748 4358 1751
rect 4362 1748 4366 1751
rect 4602 1748 4734 1751
rect 4754 1748 4758 1751
rect 4818 1748 4822 1751
rect 4882 1748 4902 1751
rect 4906 1748 4926 1751
rect 4946 1748 4966 1751
rect 4986 1748 5110 1751
rect 66 1738 134 1741
rect 138 1738 150 1741
rect 182 1738 190 1741
rect 286 1741 289 1748
rect 266 1738 289 1741
rect 334 1741 337 1748
rect 374 1741 377 1748
rect 438 1742 441 1748
rect 1382 1742 1385 1748
rect 1462 1742 1465 1748
rect 334 1738 377 1741
rect 410 1738 422 1741
rect 498 1738 502 1741
rect 690 1738 694 1741
rect 698 1738 782 1741
rect 834 1738 942 1741
rect 978 1738 1022 1741
rect 1026 1738 1102 1741
rect 1306 1738 1310 1741
rect 1602 1738 1694 1741
rect 2114 1738 2118 1741
rect 2206 1738 2230 1741
rect 2266 1738 2297 1741
rect 2322 1738 2430 1741
rect 2442 1738 2470 1741
rect 2514 1738 2542 1741
rect 2546 1738 2582 1741
rect 182 1732 185 1738
rect 614 1732 617 1738
rect 458 1728 486 1731
rect 490 1728 534 1731
rect 674 1728 694 1731
rect 830 1731 833 1738
rect 2206 1732 2209 1738
rect 2294 1732 2297 1738
rect 770 1728 833 1731
rect 994 1728 1070 1731
rect 1074 1728 1142 1731
rect 1426 1728 1566 1731
rect 1682 1728 1702 1731
rect 1802 1728 1806 1731
rect 1842 1728 1846 1731
rect 1858 1728 1982 1731
rect 2274 1728 2278 1731
rect 2298 1728 2342 1731
rect 2486 1731 2489 1738
rect 2386 1728 2489 1731
rect 2506 1728 2534 1731
rect 2606 1731 2609 1748
rect 2646 1742 2649 1748
rect 2726 1742 2729 1748
rect 2858 1738 2870 1741
rect 2874 1738 2894 1741
rect 2934 1741 2937 1748
rect 3094 1742 3097 1748
rect 2934 1738 3006 1741
rect 3010 1738 3038 1741
rect 3254 1741 3257 1748
rect 3334 1742 3337 1748
rect 3566 1742 3569 1748
rect 3254 1738 3302 1741
rect 3498 1738 3510 1741
rect 3522 1738 3534 1741
rect 3538 1738 3558 1741
rect 3722 1738 3758 1741
rect 3782 1741 3785 1748
rect 3782 1738 3806 1741
rect 4126 1738 4230 1741
rect 4298 1738 4366 1741
rect 4410 1738 4446 1741
rect 4450 1738 4510 1741
rect 4578 1738 4590 1741
rect 4610 1738 4614 1741
rect 4674 1738 4726 1741
rect 4730 1738 4766 1741
rect 4850 1738 4886 1741
rect 4890 1738 5014 1741
rect 5018 1738 5094 1741
rect 5170 1738 5238 1741
rect 2926 1732 2929 1738
rect 4126 1732 4129 1738
rect 2562 1728 2609 1731
rect 2618 1728 2662 1731
rect 2666 1728 2694 1731
rect 2706 1728 2734 1731
rect 2930 1728 2942 1731
rect 3242 1728 3462 1731
rect 3490 1728 3550 1731
rect 3554 1728 3862 1731
rect 4382 1731 4385 1738
rect 4306 1728 4385 1731
rect 4434 1728 4486 1731
rect 4530 1728 4542 1731
rect 5162 1728 5286 1731
rect 186 1718 222 1721
rect 1018 1718 1134 1721
rect 1402 1718 1766 1721
rect 1778 1718 1894 1721
rect 1930 1718 2230 1721
rect 2242 1718 2358 1721
rect 2370 1718 2566 1721
rect 2746 1718 2766 1721
rect 2770 1718 2798 1721
rect 2810 1718 2982 1721
rect 3114 1718 3142 1721
rect 3466 1718 3502 1721
rect 3682 1718 3734 1721
rect 4010 1718 4054 1721
rect 4122 1718 4153 1721
rect 4386 1718 4462 1721
rect 4558 1721 4561 1728
rect 4466 1718 4561 1721
rect 4950 1721 4953 1728
rect 4706 1718 4953 1721
rect 5106 1718 5166 1721
rect 5170 1718 5270 1721
rect 5282 1718 5286 1721
rect 542 1712 545 1718
rect 202 1708 254 1711
rect 258 1708 366 1711
rect 930 1708 1046 1711
rect 1050 1708 1166 1711
rect 1170 1708 1214 1711
rect 1218 1708 1790 1711
rect 1810 1708 1862 1711
rect 1898 1708 2046 1711
rect 2162 1708 2302 1711
rect 2306 1708 2462 1711
rect 2482 1708 2774 1711
rect 2850 1708 2870 1711
rect 2938 1708 3078 1711
rect 3346 1708 3390 1711
rect 3698 1708 3798 1711
rect 3962 1708 4142 1711
rect 4150 1711 4153 1718
rect 4150 1708 4462 1711
rect 5010 1708 5038 1711
rect 5178 1708 5238 1711
rect 5250 1708 5262 1711
rect 856 1703 858 1707
rect 862 1703 865 1707
rect 870 1703 872 1707
rect 1872 1703 1874 1707
rect 1878 1703 1881 1707
rect 1886 1703 1888 1707
rect 2904 1703 2906 1707
rect 2910 1703 2913 1707
rect 2918 1703 2920 1707
rect 3928 1703 3930 1707
rect 3934 1703 3937 1707
rect 3942 1703 3944 1707
rect 4952 1703 4954 1707
rect 4958 1703 4961 1707
rect 4966 1703 4968 1707
rect 490 1698 558 1701
rect 650 1698 694 1701
rect 762 1698 822 1701
rect 1146 1698 1222 1701
rect 1458 1698 1502 1701
rect 1618 1698 1649 1701
rect 1786 1698 1814 1701
rect 1914 1698 2062 1701
rect 2066 1698 2110 1701
rect 2186 1698 2310 1701
rect 2442 1698 2446 1701
rect 2458 1698 2574 1701
rect 3058 1698 3078 1701
rect 3426 1698 3526 1701
rect 3610 1698 3710 1701
rect 3714 1698 3830 1701
rect 3970 1698 4086 1701
rect 4338 1698 4470 1701
rect 5154 1698 5190 1701
rect 5250 1698 5294 1701
rect 50 1688 494 1691
rect 698 1688 702 1691
rect 722 1688 726 1691
rect 826 1688 886 1691
rect 906 1688 942 1691
rect 1162 1688 1182 1691
rect 1186 1688 1206 1691
rect 1210 1688 1622 1691
rect 1634 1688 1638 1691
rect 1646 1691 1649 1698
rect 1646 1688 1734 1691
rect 1818 1688 1846 1691
rect 1898 1688 1950 1691
rect 1958 1688 1966 1691
rect 1978 1688 2038 1691
rect 2050 1688 2110 1691
rect 2170 1688 2206 1691
rect 2266 1688 2294 1691
rect 2534 1688 2598 1691
rect 2818 1688 2958 1691
rect 2974 1691 2977 1698
rect 2974 1688 2990 1691
rect 3338 1688 3374 1691
rect 3378 1688 3478 1691
rect 3654 1688 3662 1691
rect 3666 1688 3718 1691
rect 3778 1688 3806 1691
rect 3826 1688 3886 1691
rect 3890 1688 4126 1691
rect 4134 1688 4257 1691
rect 314 1678 318 1681
rect 490 1678 622 1681
rect 626 1678 681 1681
rect 690 1678 694 1681
rect 714 1678 750 1681
rect 814 1681 817 1688
rect 1958 1682 1961 1688
rect 794 1678 817 1681
rect 838 1678 846 1681
rect 850 1678 862 1681
rect 890 1678 934 1681
rect 938 1678 966 1681
rect 1586 1678 1662 1681
rect 1666 1678 1670 1681
rect 1906 1678 1942 1681
rect 2058 1678 2062 1681
rect 2106 1678 2142 1681
rect 2254 1681 2257 1688
rect 2534 1682 2537 1688
rect 2226 1678 2257 1681
rect 2274 1678 2414 1681
rect 2506 1678 2510 1681
rect 2642 1678 2646 1681
rect 3050 1678 3318 1681
rect 3526 1681 3529 1688
rect 3370 1678 3529 1681
rect 3602 1678 3662 1681
rect 4134 1681 4137 1688
rect 4254 1682 4257 1688
rect 4562 1688 4582 1691
rect 4586 1688 4662 1691
rect 4802 1688 4822 1691
rect 4954 1688 5046 1691
rect 5082 1688 5110 1691
rect 5114 1688 5142 1691
rect 5146 1688 5153 1691
rect 5178 1688 5198 1691
rect 5218 1688 5238 1691
rect 4350 1682 4353 1688
rect 4114 1678 4137 1681
rect 4290 1678 4350 1681
rect 4362 1678 4422 1681
rect 4426 1678 4526 1681
rect 4578 1678 4598 1681
rect 4602 1678 4678 1681
rect 4690 1678 4766 1681
rect 4770 1678 4806 1681
rect 4842 1678 4870 1681
rect 4874 1678 5006 1681
rect 5194 1678 5214 1681
rect 5234 1678 5241 1681
rect 110 1671 113 1678
rect 166 1672 169 1678
rect 110 1668 166 1671
rect 302 1671 305 1678
rect 366 1672 369 1678
rect 302 1670 342 1671
rect 302 1668 326 1670
rect 330 1668 342 1670
rect 478 1668 486 1671
rect 546 1668 670 1671
rect 678 1671 681 1678
rect 678 1668 694 1671
rect 722 1668 758 1671
rect 770 1668 894 1671
rect 978 1668 1142 1671
rect 1486 1671 1489 1678
rect 1486 1668 1534 1671
rect 1650 1668 1654 1671
rect 1674 1668 1790 1671
rect 1794 1668 1798 1671
rect 1810 1668 1814 1671
rect 1922 1668 1934 1671
rect 1970 1668 2078 1671
rect 2086 1671 2089 1678
rect 2166 1671 2169 1678
rect 2558 1672 2561 1678
rect 2086 1668 2182 1671
rect 2226 1668 2246 1671
rect 2354 1668 2366 1671
rect 2378 1668 2454 1671
rect 2482 1668 2518 1671
rect 2778 1668 2942 1671
rect 3298 1668 3302 1671
rect 3442 1668 3638 1671
rect 3642 1668 3678 1671
rect 3714 1668 3742 1671
rect 3858 1668 3966 1671
rect 3970 1668 4006 1671
rect 4010 1668 4046 1671
rect 4166 1671 4169 1678
rect 4166 1668 4230 1671
rect 4234 1668 4294 1671
rect 4354 1668 4390 1671
rect 4418 1668 4526 1671
rect 4538 1668 4598 1671
rect 4722 1668 4782 1671
rect 4830 1671 4833 1678
rect 5150 1672 5153 1678
rect 5238 1672 5241 1678
rect 4830 1668 4886 1671
rect 4946 1668 5030 1671
rect 5178 1668 5198 1671
rect 478 1662 481 1668
rect 1598 1662 1601 1668
rect 1822 1662 1825 1668
rect 290 1658 310 1661
rect 314 1658 366 1661
rect 402 1658 422 1661
rect 442 1658 446 1661
rect 618 1658 622 1661
rect 642 1658 686 1661
rect 690 1658 782 1661
rect 850 1658 854 1661
rect 906 1658 918 1661
rect 962 1658 974 1661
rect 1058 1658 1070 1661
rect 1074 1658 1094 1661
rect 1114 1658 1174 1661
rect 1242 1658 1326 1661
rect 1682 1658 1694 1661
rect 1698 1658 1718 1661
rect 1730 1658 1790 1661
rect 1826 1658 1902 1661
rect 1914 1658 1926 1661
rect 2010 1658 2014 1661
rect 2018 1658 2022 1661
rect 2034 1658 2086 1661
rect 2374 1661 2377 1668
rect 2330 1658 2377 1661
rect 2578 1658 2614 1661
rect 2618 1658 2702 1661
rect 2706 1658 2758 1661
rect 2810 1658 2814 1661
rect 2942 1661 2945 1668
rect 2942 1658 3022 1661
rect 3026 1658 3078 1661
rect 4502 1662 4505 1668
rect 3250 1659 3462 1661
rect 3246 1658 3462 1659
rect 3474 1658 3478 1661
rect 3514 1658 3550 1661
rect 3570 1658 3574 1661
rect 4218 1658 4270 1661
rect 4274 1658 4310 1661
rect 4522 1658 4582 1661
rect 4626 1658 4638 1661
rect 4662 1661 4665 1668
rect 4918 1662 4921 1668
rect 5198 1662 5201 1668
rect 4662 1658 4686 1661
rect 4730 1658 4758 1661
rect 4774 1658 4798 1661
rect 5106 1658 5182 1661
rect 5202 1658 5222 1661
rect 5262 1661 5265 1688
rect 5262 1658 5270 1661
rect 5342 1661 5346 1662
rect 5314 1658 5346 1661
rect 3950 1652 3953 1658
rect 4774 1652 4777 1658
rect 170 1648 238 1651
rect 242 1648 262 1651
rect 370 1648 401 1651
rect 570 1648 633 1651
rect 786 1648 846 1651
rect 890 1648 902 1651
rect 946 1648 974 1651
rect 978 1648 1065 1651
rect 1082 1648 1134 1651
rect 1138 1648 1182 1651
rect 1186 1648 1270 1651
rect 1290 1648 1318 1651
rect 1490 1648 1622 1651
rect 1682 1648 1718 1651
rect 1730 1648 1878 1651
rect 1898 1648 1966 1651
rect 1994 1648 2006 1651
rect 2202 1648 2270 1651
rect 2314 1648 2342 1651
rect 2346 1648 2366 1651
rect 2394 1648 2406 1651
rect 2466 1648 2470 1651
rect 2514 1648 2518 1651
rect 2594 1648 2622 1651
rect 2626 1648 2646 1651
rect 2754 1648 2910 1651
rect 3194 1648 3302 1651
rect 3306 1648 3446 1651
rect 3450 1648 3486 1651
rect 3514 1648 3518 1651
rect 3550 1648 3566 1651
rect 3570 1648 3590 1651
rect 3594 1648 3614 1651
rect 4266 1648 4286 1651
rect 4346 1648 4510 1651
rect 4690 1648 4750 1651
rect 4850 1648 5014 1651
rect 5178 1648 5214 1651
rect 398 1642 401 1648
rect 630 1642 633 1648
rect 1062 1642 1065 1648
rect 282 1638 294 1641
rect 578 1638 598 1641
rect 746 1638 750 1641
rect 754 1638 1038 1641
rect 1082 1638 1110 1641
rect 1338 1638 1686 1641
rect 1730 1638 1742 1641
rect 1858 1638 1878 1641
rect 1906 1638 2742 1641
rect 3322 1638 3382 1641
rect 3550 1641 3553 1648
rect 4886 1642 4889 1648
rect 3498 1638 3553 1641
rect 3562 1638 3566 1641
rect 3586 1638 3702 1641
rect 4162 1638 4246 1641
rect 4250 1638 4366 1641
rect 4450 1638 4502 1641
rect 4610 1638 4622 1641
rect 4626 1638 4694 1641
rect 162 1628 510 1631
rect 546 1628 630 1631
rect 802 1628 886 1631
rect 890 1628 1102 1631
rect 1126 1631 1129 1638
rect 1114 1628 1129 1631
rect 1666 1628 1782 1631
rect 1922 1628 1974 1631
rect 2130 1628 2190 1631
rect 2218 1628 2542 1631
rect 2570 1628 3566 1631
rect 3570 1628 3838 1631
rect 3906 1628 4678 1631
rect 26 1618 54 1621
rect 58 1618 278 1621
rect 810 1618 894 1621
rect 938 1618 1398 1621
rect 1498 1618 1846 1621
rect 1962 1618 2166 1621
rect 2402 1618 2854 1621
rect 2922 1618 3118 1621
rect 3122 1618 4190 1621
rect 4194 1618 4302 1621
rect 4658 1618 4790 1621
rect 250 1608 326 1611
rect 650 1608 830 1611
rect 922 1608 961 1611
rect 970 1608 974 1611
rect 1410 1608 1718 1611
rect 1834 1608 1854 1611
rect 2250 1608 2350 1611
rect 2698 1608 2790 1611
rect 3098 1608 3254 1611
rect 3258 1608 3398 1611
rect 3402 1608 3406 1611
rect 3682 1608 3686 1611
rect 3698 1608 4150 1611
rect 4154 1608 4430 1611
rect 344 1603 346 1607
rect 350 1603 353 1607
rect 358 1603 360 1607
rect 818 1598 878 1601
rect 906 1598 950 1601
rect 958 1601 961 1608
rect 1368 1603 1370 1607
rect 1374 1603 1377 1607
rect 1382 1603 1384 1607
rect 2030 1602 2033 1608
rect 2392 1603 2394 1607
rect 2398 1603 2401 1607
rect 2406 1603 2408 1607
rect 3416 1603 3418 1607
rect 3422 1603 3425 1607
rect 3430 1603 3432 1607
rect 4440 1603 4442 1607
rect 4446 1603 4449 1607
rect 4454 1603 4456 1607
rect 958 1598 998 1601
rect 1570 1598 1846 1601
rect 2146 1598 2382 1601
rect 3674 1598 3966 1601
rect 4810 1598 4822 1601
rect 4978 1598 5214 1601
rect 162 1588 998 1591
rect 1162 1588 1334 1591
rect 1338 1588 1702 1591
rect 2010 1588 2262 1591
rect 2310 1588 2318 1591
rect 2322 1588 2446 1591
rect 2634 1588 2646 1591
rect 2978 1588 3134 1591
rect 3138 1588 4126 1591
rect 4146 1588 4662 1591
rect 4802 1588 4814 1591
rect 4818 1588 4910 1591
rect 4914 1588 5134 1591
rect 110 1581 113 1588
rect 98 1578 113 1581
rect 642 1578 681 1581
rect 714 1578 822 1581
rect 1042 1578 1694 1581
rect 1698 1578 2078 1581
rect 2250 1578 2294 1581
rect 2298 1578 2406 1581
rect 4098 1578 4478 1581
rect 4938 1578 5126 1581
rect 678 1572 681 1578
rect 90 1568 134 1571
rect 258 1568 382 1571
rect 386 1568 390 1571
rect 394 1568 414 1571
rect 794 1568 814 1571
rect 970 1568 974 1571
rect 1018 1568 1054 1571
rect 1074 1568 1142 1571
rect 1146 1568 1510 1571
rect 1538 1568 1854 1571
rect 1922 1568 1934 1571
rect 2194 1568 2294 1571
rect 2298 1568 2302 1571
rect 2506 1568 2742 1571
rect 2770 1568 3150 1571
rect 4498 1568 4598 1571
rect 4602 1568 4646 1571
rect 4746 1568 4782 1571
rect 4810 1568 4897 1571
rect 5018 1568 5038 1571
rect 66 1558 158 1561
rect 178 1558 182 1561
rect 298 1558 310 1561
rect 314 1558 318 1561
rect 322 1558 358 1561
rect 562 1558 590 1561
rect 654 1561 657 1568
rect 594 1558 657 1561
rect 818 1558 838 1561
rect 906 1558 910 1561
rect 914 1558 998 1561
rect 1002 1558 1206 1561
rect 1214 1558 1646 1561
rect 1738 1558 1766 1561
rect 1930 1558 1950 1561
rect 1954 1558 1958 1561
rect 2054 1558 2102 1561
rect 2414 1561 2417 1568
rect 4894 1562 4897 1568
rect 2330 1558 2417 1561
rect 2594 1558 2998 1561
rect 3186 1558 3190 1561
rect 3346 1558 3366 1561
rect 3674 1558 3686 1561
rect 4250 1558 4422 1561
rect 4538 1558 4558 1561
rect 4714 1558 4734 1561
rect 4738 1558 4758 1561
rect 4770 1558 4798 1561
rect 4922 1558 4974 1561
rect 5062 1561 5065 1568
rect 5034 1558 5174 1561
rect 5218 1558 5230 1561
rect 50 1548 190 1551
rect 194 1548 214 1551
rect 234 1548 286 1551
rect 290 1548 334 1551
rect 338 1548 374 1551
rect 378 1548 385 1551
rect 434 1548 617 1551
rect 658 1548 662 1551
rect 722 1548 742 1551
rect 770 1548 806 1551
rect 834 1548 870 1551
rect 874 1548 894 1551
rect 930 1548 942 1551
rect 946 1548 950 1551
rect 1002 1548 1006 1551
rect 1130 1548 1166 1551
rect 1214 1551 1217 1558
rect 1686 1552 1689 1558
rect 2054 1552 2057 1558
rect 2278 1552 2281 1558
rect 1170 1548 1217 1551
rect 1322 1548 1502 1551
rect 1582 1548 1614 1551
rect 1754 1548 1758 1551
rect 1826 1548 1942 1551
rect 1962 1548 2054 1551
rect 2098 1548 2134 1551
rect 2210 1548 2222 1551
rect 2290 1548 2294 1551
rect 2370 1548 2446 1551
rect 2674 1548 2678 1551
rect 2754 1548 2822 1551
rect 2826 1548 3022 1551
rect 3026 1548 3038 1551
rect 3086 1551 3089 1558
rect 3134 1551 3137 1558
rect 3086 1548 3137 1551
rect 3154 1548 3254 1551
rect 3258 1548 3302 1551
rect 3306 1548 3342 1551
rect 3346 1548 3422 1551
rect 3522 1548 3526 1551
rect 3630 1548 3646 1551
rect 3758 1551 3761 1558
rect 4478 1552 4481 1558
rect 3722 1548 3761 1551
rect 3786 1548 3918 1551
rect 3978 1548 4014 1551
rect 4018 1548 4022 1551
rect 614 1542 617 1548
rect 18 1538 78 1541
rect 82 1538 102 1541
rect 186 1538 206 1541
rect 210 1538 222 1541
rect 306 1538 342 1541
rect 618 1538 646 1541
rect 650 1538 654 1541
rect 722 1538 726 1541
rect 738 1538 846 1541
rect 918 1541 921 1548
rect 850 1538 921 1541
rect 938 1538 950 1541
rect 954 1538 1022 1541
rect 1078 1541 1081 1548
rect 1582 1542 1585 1548
rect 1050 1538 1081 1541
rect 1090 1538 1094 1541
rect 1122 1538 1134 1541
rect 1146 1538 1150 1541
rect 1170 1538 1174 1541
rect 1254 1538 1310 1541
rect 1682 1538 1686 1541
rect 1754 1538 1766 1541
rect 1770 1538 1982 1541
rect 1994 1538 1998 1541
rect 2042 1538 2062 1541
rect 2066 1538 2073 1541
rect 2090 1538 2158 1541
rect 2162 1538 2174 1541
rect 2370 1538 2582 1541
rect 2606 1541 2609 1548
rect 2702 1542 2705 1548
rect 3630 1542 3633 1548
rect 4210 1548 4214 1551
rect 4386 1548 4406 1551
rect 4514 1548 4542 1551
rect 4578 1548 4686 1551
rect 4770 1548 4798 1551
rect 4802 1548 4814 1551
rect 4858 1548 5054 1551
rect 5058 1548 5065 1551
rect 5090 1548 5158 1551
rect 2606 1538 2702 1541
rect 2878 1538 2974 1541
rect 3034 1538 3038 1541
rect 3250 1538 3262 1541
rect 3266 1538 3310 1541
rect 3362 1538 3382 1541
rect 3394 1538 3414 1541
rect 3418 1538 3462 1541
rect 3678 1538 3702 1541
rect 3706 1538 3822 1541
rect 3906 1538 3974 1541
rect 3978 1538 3990 1541
rect 3994 1538 4014 1541
rect 4246 1541 4249 1548
rect 4162 1538 4249 1541
rect 4358 1541 4361 1548
rect 4358 1538 4374 1541
rect 4418 1538 4486 1541
rect 4546 1538 4582 1541
rect 4826 1538 4918 1541
rect 5018 1538 5046 1541
rect 5050 1538 5054 1541
rect 5082 1538 5097 1541
rect 5210 1538 5238 1541
rect 110 1531 113 1538
rect 478 1532 481 1538
rect 534 1532 537 1538
rect 110 1528 254 1531
rect 322 1528 398 1531
rect 602 1528 654 1531
rect 674 1528 678 1531
rect 722 1528 758 1531
rect 934 1531 937 1538
rect 794 1528 937 1531
rect 1034 1528 1054 1531
rect 1058 1528 1126 1531
rect 1166 1531 1169 1538
rect 1146 1528 1169 1531
rect 1254 1532 1257 1538
rect 1494 1532 1497 1538
rect 2078 1532 2081 1538
rect 2182 1532 2185 1538
rect 2878 1532 2881 1538
rect 3678 1532 3681 1538
rect 1450 1528 1481 1531
rect 1706 1528 1758 1531
rect 1810 1528 1878 1531
rect 1890 1528 1894 1531
rect 1922 1528 1950 1531
rect 1954 1528 1966 1531
rect 1994 1528 2046 1531
rect 2050 1528 2054 1531
rect 2098 1528 2102 1531
rect 2346 1528 2718 1531
rect 3338 1528 3358 1531
rect 4442 1528 4446 1531
rect 4518 1531 4521 1538
rect 4498 1528 4521 1531
rect 4614 1532 4617 1538
rect 5094 1532 5097 1538
rect 4642 1528 4926 1531
rect 4994 1528 5006 1531
rect 5270 1531 5273 1548
rect 5250 1528 5273 1531
rect 42 1518 134 1521
rect 138 1518 510 1521
rect 610 1518 702 1521
rect 782 1521 785 1528
rect 1478 1522 1481 1528
rect 738 1518 785 1521
rect 842 1518 1374 1521
rect 1514 1518 1897 1521
rect 1994 1518 2006 1521
rect 2238 1521 2241 1528
rect 2042 1518 2241 1521
rect 2578 1518 2918 1521
rect 2954 1518 2982 1521
rect 3010 1518 3190 1521
rect 3626 1518 3670 1521
rect 3674 1518 3718 1521
rect 3730 1518 4270 1521
rect 4346 1518 4486 1521
rect 4630 1521 4633 1528
rect 4506 1518 4633 1521
rect 4698 1518 4710 1521
rect 4794 1518 4862 1521
rect 4946 1518 5070 1521
rect 5074 1518 5102 1521
rect 5178 1518 5182 1521
rect 5210 1518 5270 1521
rect 5282 1518 5302 1521
rect 106 1508 158 1511
rect 466 1508 502 1511
rect 690 1508 846 1511
rect 1722 1508 1798 1511
rect 1894 1511 1897 1518
rect 1894 1508 2022 1511
rect 2026 1508 2110 1511
rect 2154 1508 2318 1511
rect 2482 1508 2782 1511
rect 3234 1508 3350 1511
rect 3418 1508 3502 1511
rect 3506 1508 3686 1511
rect 3754 1508 3862 1511
rect 4090 1508 4102 1511
rect 4290 1508 4342 1511
rect 4354 1508 4374 1511
rect 4418 1508 4510 1511
rect 4578 1508 4598 1511
rect 4602 1508 4734 1511
rect 5018 1508 5150 1511
rect 5154 1508 5166 1511
rect 190 1502 193 1508
rect 856 1503 858 1507
rect 862 1503 865 1507
rect 870 1503 872 1507
rect 1872 1503 1874 1507
rect 1878 1503 1881 1507
rect 1886 1503 1888 1507
rect 2904 1503 2906 1507
rect 2910 1503 2913 1507
rect 2918 1503 2920 1507
rect 3928 1503 3930 1507
rect 3934 1503 3937 1507
rect 3942 1503 3944 1507
rect 4952 1503 4954 1507
rect 4958 1503 4961 1507
rect 4966 1503 4968 1507
rect 42 1498 94 1501
rect 626 1498 742 1501
rect 1466 1498 1862 1501
rect 2074 1498 2094 1501
rect 2114 1498 2190 1501
rect 2202 1498 2278 1501
rect 2386 1498 2414 1501
rect 2522 1498 2534 1501
rect 2610 1498 2846 1501
rect 2978 1498 3110 1501
rect 3114 1498 3222 1501
rect 3226 1498 3310 1501
rect 3314 1498 3550 1501
rect 3554 1498 3630 1501
rect 3634 1498 3838 1501
rect 3978 1498 4318 1501
rect 4410 1498 4526 1501
rect 4530 1498 4710 1501
rect 5302 1492 5305 1498
rect 98 1488 198 1491
rect 202 1488 222 1491
rect 282 1488 470 1491
rect 554 1488 710 1491
rect 730 1488 766 1491
rect 850 1488 902 1491
rect 1122 1488 1126 1491
rect 1498 1488 1521 1491
rect 1518 1482 1521 1488
rect 1626 1488 1710 1491
rect 1714 1488 1721 1491
rect 1818 1488 1894 1491
rect 1918 1488 1926 1491
rect 1930 1488 2014 1491
rect 2026 1488 2102 1491
rect 2122 1488 2142 1491
rect 2186 1488 2190 1491
rect 2610 1488 2654 1491
rect 2658 1488 2670 1491
rect 2906 1488 2926 1491
rect 3090 1488 3278 1491
rect 3394 1488 3494 1491
rect 3514 1488 3550 1491
rect 3610 1488 3774 1491
rect 4010 1488 4174 1491
rect 4258 1488 4262 1491
rect 4474 1488 4542 1491
rect 4570 1488 4606 1491
rect 4610 1488 4702 1491
rect 4770 1488 5110 1491
rect 5282 1488 5294 1491
rect 74 1478 177 1481
rect 186 1478 206 1481
rect 250 1478 254 1481
rect 426 1478 486 1481
rect 490 1478 494 1481
rect 690 1478 734 1481
rect 746 1478 774 1481
rect 782 1478 1222 1481
rect 1298 1478 1334 1481
rect 1490 1478 1510 1481
rect 1526 1481 1529 1488
rect 1526 1478 1558 1481
rect 1722 1478 1758 1481
rect 1766 1481 1769 1488
rect 1766 1478 1790 1481
rect 1826 1478 1902 1481
rect 1906 1478 1974 1481
rect 1986 1478 2246 1481
rect 2250 1478 2270 1481
rect 2282 1478 2302 1481
rect 2370 1478 2486 1481
rect 2498 1478 2510 1481
rect 2722 1478 2742 1481
rect 3002 1478 3022 1481
rect 3026 1478 3190 1481
rect 3290 1478 3294 1481
rect 3338 1478 3342 1481
rect 3386 1478 3481 1481
rect 3554 1478 3630 1481
rect 3634 1478 3782 1481
rect 4074 1478 4086 1481
rect 4090 1478 4134 1481
rect 4374 1481 4377 1488
rect 4414 1481 4417 1488
rect 4374 1478 4417 1481
rect 4498 1478 4582 1481
rect 4586 1478 4590 1481
rect 4850 1478 4886 1481
rect 4890 1478 4918 1481
rect 5066 1478 5134 1481
rect 5142 1478 5150 1481
rect 5154 1478 5190 1481
rect 5250 1478 5278 1481
rect 174 1472 177 1478
rect 210 1468 310 1471
rect 698 1468 734 1471
rect 782 1471 785 1478
rect 1342 1472 1345 1478
rect 762 1468 785 1471
rect 878 1468 1158 1471
rect 1250 1468 1302 1471
rect 1482 1468 1502 1471
rect 1522 1468 1566 1471
rect 1738 1468 1750 1471
rect 1754 1468 1862 1471
rect 1914 1468 1934 1471
rect 2002 1468 2006 1471
rect 2026 1468 2030 1471
rect 2034 1468 2038 1471
rect 2106 1468 2118 1471
rect 2138 1468 2166 1471
rect 2482 1468 2494 1471
rect 2714 1468 2758 1471
rect 2862 1471 2865 1478
rect 3478 1472 3481 1478
rect 3894 1472 3897 1478
rect 2862 1468 2926 1471
rect 3018 1468 3046 1471
rect 3218 1468 3246 1471
rect 3250 1468 3406 1471
rect 3482 1468 3518 1471
rect 3522 1468 3574 1471
rect 3586 1468 3606 1471
rect 3682 1468 3726 1471
rect 3898 1468 3918 1471
rect 4458 1468 4478 1471
rect 4514 1468 4542 1471
rect 4554 1468 4582 1471
rect 4806 1471 4809 1478
rect 4786 1468 4809 1471
rect 4818 1468 4846 1471
rect 4922 1468 4942 1471
rect 4978 1468 4982 1471
rect 4990 1471 4993 1478
rect 4990 1468 5030 1471
rect 5050 1468 5054 1471
rect 5142 1471 5145 1478
rect 5106 1468 5145 1471
rect 5150 1468 5158 1471
rect 5162 1468 5174 1471
rect 5234 1468 5246 1471
rect 10 1458 70 1461
rect 106 1458 134 1461
rect 218 1458 326 1461
rect 422 1458 457 1461
rect 646 1461 649 1468
rect 642 1458 649 1461
rect 862 1462 865 1468
rect 878 1462 881 1468
rect 990 1462 993 1468
rect 1110 1462 1113 1468
rect 1190 1462 1193 1468
rect 1302 1462 1305 1468
rect 1026 1458 1030 1461
rect 1094 1458 1102 1461
rect 1310 1461 1313 1468
rect 1310 1458 1334 1461
rect 1514 1458 1518 1461
rect 1706 1458 1710 1461
rect 1746 1458 1750 1461
rect 1826 1458 1862 1461
rect 1914 1458 1958 1461
rect 2010 1458 2030 1461
rect 2090 1458 2198 1461
rect 2202 1459 2222 1461
rect 2278 1462 2281 1468
rect 2202 1458 2225 1459
rect 2466 1458 2486 1461
rect 2498 1458 2774 1461
rect 2778 1458 2782 1461
rect 3002 1458 3038 1461
rect 3042 1458 3094 1461
rect 3178 1458 3958 1461
rect 3974 1461 3977 1468
rect 3974 1458 4089 1461
rect 4150 1461 4153 1468
rect 4662 1462 4665 1468
rect 4122 1458 4153 1461
rect 4202 1458 4206 1461
rect 4298 1458 4318 1461
rect 4682 1458 4694 1461
rect 4754 1458 4774 1461
rect 4778 1458 4894 1461
rect 5002 1458 5030 1461
rect 5114 1458 5142 1461
rect 5154 1458 5174 1461
rect 5210 1458 5254 1461
rect 5270 1461 5273 1468
rect 5270 1458 5310 1461
rect 5342 1461 5346 1462
rect 5314 1458 5346 1461
rect 422 1452 425 1458
rect 454 1452 457 1458
rect 1094 1452 1097 1458
rect 50 1448 230 1451
rect 650 1448 694 1451
rect 1234 1448 1238 1451
rect 1294 1451 1297 1458
rect 1258 1448 1297 1451
rect 1358 1451 1361 1458
rect 1322 1448 1361 1451
rect 1646 1451 1649 1458
rect 2006 1452 2009 1458
rect 2462 1452 2465 1458
rect 2958 1452 2961 1458
rect 4086 1452 4089 1458
rect 1394 1448 1649 1451
rect 1766 1448 1782 1451
rect 1818 1448 1926 1451
rect 1930 1448 1934 1451
rect 2026 1448 2046 1451
rect 2138 1448 2182 1451
rect 2314 1448 2334 1451
rect 2634 1448 2694 1451
rect 2698 1448 2710 1451
rect 2746 1448 2750 1451
rect 3046 1448 3102 1451
rect 3106 1448 3158 1451
rect 3186 1448 3326 1451
rect 3330 1448 3654 1451
rect 3658 1448 3686 1451
rect 3706 1448 3766 1451
rect 3782 1448 3822 1451
rect 4154 1448 4158 1451
rect 4470 1451 4473 1458
rect 4442 1448 4473 1451
rect 4490 1448 4510 1451
rect 4794 1448 4814 1451
rect 4890 1448 5230 1451
rect 226 1438 374 1441
rect 666 1438 806 1441
rect 978 1438 1182 1441
rect 1310 1441 1313 1448
rect 1766 1442 1769 1448
rect 2134 1442 2137 1448
rect 3046 1442 3049 1448
rect 1282 1438 1646 1441
rect 1794 1438 1894 1441
rect 1906 1438 1982 1441
rect 2290 1438 2302 1441
rect 2458 1438 2641 1441
rect 2658 1438 2790 1441
rect 2850 1438 3014 1441
rect 3158 1441 3161 1448
rect 3782 1442 3785 1448
rect 3158 1438 3230 1441
rect 3234 1438 3294 1441
rect 3354 1438 3382 1441
rect 3458 1438 3473 1441
rect 3506 1438 3654 1441
rect 3794 1438 4142 1441
rect 4146 1438 4326 1441
rect 4394 1438 4558 1441
rect 4642 1438 5102 1441
rect 5106 1438 5126 1441
rect 5130 1438 5182 1441
rect 2638 1432 2641 1438
rect 3470 1432 3473 1438
rect 386 1428 534 1431
rect 538 1428 558 1431
rect 1314 1428 1390 1431
rect 1634 1428 1654 1431
rect 1770 1428 1774 1431
rect 1906 1428 1910 1431
rect 1946 1428 2150 1431
rect 2154 1428 2174 1431
rect 2178 1428 2310 1431
rect 2442 1428 2561 1431
rect 3194 1428 3214 1431
rect 3218 1428 3462 1431
rect 3498 1428 3702 1431
rect 3706 1428 3766 1431
rect 3810 1428 4262 1431
rect 4266 1428 4294 1431
rect 4302 1428 4638 1431
rect 4802 1428 4822 1431
rect 4834 1428 4846 1431
rect 4970 1428 5006 1431
rect 5010 1428 5110 1431
rect 22 1421 25 1428
rect 22 1418 222 1421
rect 562 1418 790 1421
rect 962 1418 1022 1421
rect 1690 1418 1822 1421
rect 1842 1418 1870 1421
rect 1874 1418 1918 1421
rect 2066 1418 2214 1421
rect 2218 1418 2526 1421
rect 2538 1418 2550 1421
rect 2558 1421 2561 1428
rect 2558 1418 2870 1421
rect 3370 1418 3558 1421
rect 3626 1418 3646 1421
rect 4302 1421 4305 1428
rect 4050 1418 4305 1421
rect 4314 1418 4470 1421
rect 5002 1418 5062 1421
rect 5178 1418 5214 1421
rect 26 1408 46 1411
rect 746 1408 1158 1411
rect 1714 1408 1950 1411
rect 2146 1408 2174 1411
rect 2682 1408 2862 1411
rect 4154 1408 4198 1411
rect 4914 1408 5190 1411
rect 5194 1408 5262 1411
rect 344 1403 346 1407
rect 350 1403 353 1407
rect 358 1403 360 1407
rect 1368 1403 1370 1407
rect 1374 1403 1377 1407
rect 1382 1403 1384 1407
rect 2392 1403 2394 1407
rect 2398 1403 2401 1407
rect 2406 1403 2408 1407
rect 3416 1403 3418 1407
rect 3422 1403 3425 1407
rect 3430 1403 3432 1407
rect 4440 1403 4442 1407
rect 4446 1403 4449 1407
rect 4454 1403 4456 1407
rect 690 1398 1134 1401
rect 1466 1398 1758 1401
rect 1802 1398 2038 1401
rect 2042 1398 2142 1401
rect 2146 1398 2222 1401
rect 2730 1398 2982 1401
rect 3514 1398 3790 1401
rect 3794 1398 3846 1401
rect 4018 1398 4150 1401
rect 130 1388 1174 1391
rect 1330 1388 1478 1391
rect 1482 1388 1550 1391
rect 1570 1388 1806 1391
rect 1858 1388 1934 1391
rect 1946 1388 1974 1391
rect 1978 1388 2958 1391
rect 2978 1388 3190 1391
rect 3314 1388 3318 1391
rect 3530 1388 3566 1391
rect 4130 1388 4270 1391
rect 4274 1388 4334 1391
rect 4338 1388 4350 1391
rect 4858 1388 4862 1391
rect 98 1378 118 1381
rect 122 1378 278 1381
rect 450 1378 486 1381
rect 490 1378 542 1381
rect 1338 1378 1838 1381
rect 1898 1378 1918 1381
rect 1930 1378 2078 1381
rect 2114 1378 2230 1381
rect 2234 1378 2241 1381
rect 2250 1378 2342 1381
rect 2474 1378 2686 1381
rect 2754 1378 2806 1381
rect 3066 1378 3102 1381
rect 3106 1378 3142 1381
rect 3146 1378 4102 1381
rect 4502 1381 4505 1388
rect 4322 1378 4505 1381
rect 62 1371 65 1378
rect 50 1368 65 1371
rect 430 1371 433 1378
rect 314 1368 433 1371
rect 962 1368 966 1371
rect 1110 1371 1113 1378
rect 1010 1368 1113 1371
rect 1122 1368 1134 1371
rect 1186 1368 1470 1371
rect 1810 1368 1862 1371
rect 1866 1368 4198 1371
rect 4466 1368 4470 1371
rect 4490 1368 4654 1371
rect 4682 1368 4766 1371
rect 5214 1371 5217 1378
rect 5238 1371 5241 1378
rect 5214 1368 5278 1371
rect 50 1358 54 1361
rect 90 1358 110 1361
rect 138 1358 286 1361
rect 302 1361 305 1368
rect 302 1358 366 1361
rect 422 1358 430 1361
rect 434 1358 438 1361
rect 474 1358 494 1361
rect 498 1358 606 1361
rect 634 1358 670 1361
rect 818 1358 822 1361
rect 922 1358 1006 1361
rect 1042 1358 1054 1361
rect 1058 1358 1062 1361
rect 1090 1358 1142 1361
rect 1146 1358 1382 1361
rect 1738 1358 2030 1361
rect 2122 1358 2126 1361
rect 2194 1358 2198 1361
rect 2210 1358 2222 1361
rect 2226 1358 2246 1361
rect 2274 1358 2326 1361
rect 2330 1358 2350 1361
rect 2386 1358 2398 1361
rect 2610 1358 2622 1361
rect 2666 1358 2934 1361
rect 2938 1358 2942 1361
rect 3594 1358 3654 1361
rect 3722 1358 3758 1361
rect 3826 1358 3886 1361
rect 4082 1358 4174 1361
rect 4178 1358 4214 1361
rect 4222 1361 4225 1368
rect 4222 1358 4262 1361
rect 4266 1358 4302 1361
rect 4370 1358 4502 1361
rect 4506 1358 4510 1361
rect 4602 1358 4702 1361
rect 4870 1361 4873 1368
rect 4850 1358 4873 1361
rect 5210 1358 5230 1361
rect 5234 1358 5262 1361
rect 218 1348 254 1351
rect 382 1351 385 1358
rect 362 1348 385 1351
rect 410 1348 518 1351
rect 554 1348 582 1351
rect 586 1348 614 1351
rect 618 1348 662 1351
rect 1010 1348 1014 1351
rect 1050 1348 1070 1351
rect 1138 1348 1166 1351
rect 1170 1348 1174 1351
rect 1770 1348 1878 1351
rect 1882 1348 1918 1351
rect 2018 1348 2150 1351
rect 2186 1348 2190 1351
rect 2250 1348 2254 1351
rect 2282 1348 2406 1351
rect 2554 1348 3030 1351
rect 3246 1351 3249 1358
rect 3534 1352 3537 1358
rect 3210 1348 3249 1351
rect 3442 1348 3518 1351
rect 3546 1348 3966 1351
rect 3970 1348 3985 1351
rect 750 1342 753 1348
rect 74 1338 94 1341
rect 314 1338 366 1341
rect 394 1338 462 1341
rect 490 1338 518 1341
rect 522 1338 558 1341
rect 898 1338 934 1341
rect 938 1338 974 1341
rect 1026 1338 1054 1341
rect 1082 1338 1086 1341
rect 1098 1338 1126 1341
rect 1130 1338 1142 1341
rect 1146 1338 1182 1341
rect 1186 1338 1390 1341
rect 1462 1341 1465 1348
rect 1614 1342 1617 1348
rect 1462 1338 1542 1341
rect 1630 1341 1633 1348
rect 2422 1342 2425 1348
rect 2550 1342 2553 1348
rect 1630 1338 1678 1341
rect 1794 1338 1798 1341
rect 1874 1338 1878 1341
rect 1906 1338 1934 1341
rect 1938 1338 1969 1341
rect 2106 1338 2110 1341
rect 2218 1338 2230 1341
rect 2234 1338 2238 1341
rect 2290 1338 2374 1341
rect 2530 1338 2534 1341
rect 2714 1338 2822 1341
rect 3002 1338 3054 1341
rect 3058 1338 3094 1341
rect 3098 1338 3118 1341
rect 3150 1341 3153 1348
rect 3982 1342 3985 1348
rect 4014 1348 4030 1351
rect 4034 1348 4086 1351
rect 4202 1348 4230 1351
rect 4290 1348 4294 1351
rect 4342 1351 4345 1358
rect 4902 1352 4905 1358
rect 4342 1348 4406 1351
rect 4554 1348 4622 1351
rect 4634 1348 4686 1351
rect 4690 1348 4902 1351
rect 5034 1348 5038 1351
rect 5154 1348 5158 1351
rect 5186 1348 5198 1351
rect 4014 1342 4017 1348
rect 3122 1338 3174 1341
rect 3498 1338 3542 1341
rect 3546 1338 3590 1341
rect 3594 1338 3678 1341
rect 3682 1338 3790 1341
rect 3794 1338 3814 1341
rect 3818 1338 3822 1341
rect 4098 1338 4238 1341
rect 4266 1338 4310 1341
rect 4402 1338 4566 1341
rect 4570 1338 4609 1341
rect 1814 1332 1817 1338
rect 66 1328 78 1331
rect 146 1328 198 1331
rect 202 1328 230 1331
rect 274 1328 318 1331
rect 386 1328 390 1331
rect 482 1328 486 1331
rect 626 1328 902 1331
rect 962 1328 998 1331
rect 1266 1328 1310 1331
rect 1314 1328 1478 1331
rect 1922 1328 1926 1331
rect 1966 1331 1969 1338
rect 2374 1332 2377 1338
rect 2390 1332 2393 1338
rect 4606 1332 4609 1338
rect 4834 1338 4846 1341
rect 4850 1338 4870 1341
rect 4974 1341 4977 1348
rect 4974 1338 5006 1341
rect 5018 1338 5094 1341
rect 5114 1338 5142 1341
rect 5150 1338 5166 1341
rect 4790 1332 4793 1338
rect 5150 1332 5153 1338
rect 1966 1328 2110 1331
rect 2114 1328 2126 1331
rect 2170 1328 2182 1331
rect 2234 1328 2262 1331
rect 2546 1328 2550 1331
rect 2666 1328 2710 1331
rect 2810 1328 2830 1331
rect 2834 1328 2910 1331
rect 2946 1328 2990 1331
rect 3202 1328 3230 1331
rect 3410 1328 3494 1331
rect 3554 1328 3598 1331
rect 3714 1328 3774 1331
rect 3778 1328 3806 1331
rect 4218 1328 4262 1331
rect 4294 1328 4302 1331
rect 4306 1328 4350 1331
rect 4490 1328 4518 1331
rect 4850 1328 4862 1331
rect 4866 1328 4886 1331
rect 4930 1328 4961 1331
rect 5058 1328 5134 1331
rect 5186 1328 5246 1331
rect 5250 1328 5278 1331
rect 270 1321 273 1328
rect 218 1318 273 1321
rect 458 1318 510 1321
rect 558 1321 561 1328
rect 514 1318 561 1321
rect 682 1318 694 1321
rect 706 1318 814 1321
rect 818 1318 838 1321
rect 994 1318 1014 1321
rect 1150 1321 1153 1328
rect 1018 1318 1153 1321
rect 1186 1318 1262 1321
rect 1274 1318 1398 1321
rect 1442 1318 1494 1321
rect 1498 1318 1638 1321
rect 1690 1318 1734 1321
rect 1810 1318 1894 1321
rect 1922 1318 1926 1321
rect 1970 1318 1974 1321
rect 2138 1318 2310 1321
rect 2314 1318 2366 1321
rect 2386 1318 2574 1321
rect 2594 1318 2630 1321
rect 2766 1321 2769 1328
rect 3006 1321 3009 1328
rect 2658 1318 2769 1321
rect 2774 1318 3009 1321
rect 3018 1318 3366 1321
rect 3378 1318 3830 1321
rect 3834 1318 4702 1321
rect 4714 1318 4742 1321
rect 4746 1318 4798 1321
rect 4802 1318 4950 1321
rect 4958 1321 4961 1328
rect 4958 1318 5073 1321
rect 226 1308 310 1311
rect 418 1308 766 1311
rect 890 1308 1422 1311
rect 1702 1308 1798 1311
rect 1962 1308 2190 1311
rect 2194 1308 2294 1311
rect 2346 1308 2382 1311
rect 2466 1308 2470 1311
rect 2774 1311 2777 1318
rect 5070 1312 5073 1318
rect 2478 1308 2777 1311
rect 2978 1308 2998 1311
rect 3650 1308 3662 1311
rect 3666 1308 3694 1311
rect 4170 1308 4246 1311
rect 4698 1308 4742 1311
rect 5130 1308 5278 1311
rect 856 1303 858 1307
rect 862 1303 865 1307
rect 870 1303 872 1307
rect 450 1298 494 1301
rect 498 1298 526 1301
rect 546 1298 550 1301
rect 554 1298 582 1301
rect 946 1298 1030 1301
rect 1354 1298 1374 1301
rect 1702 1301 1705 1308
rect 1846 1302 1849 1308
rect 1872 1303 1874 1307
rect 1878 1303 1881 1307
rect 1886 1303 1888 1307
rect 1378 1298 1705 1301
rect 1722 1298 1734 1301
rect 2050 1298 2334 1301
rect 2478 1301 2481 1308
rect 2904 1303 2906 1307
rect 2910 1303 2913 1307
rect 2918 1303 2920 1307
rect 3928 1303 3930 1307
rect 3934 1303 3937 1307
rect 3942 1303 3944 1307
rect 4952 1303 4954 1307
rect 4958 1303 4961 1307
rect 4966 1303 4968 1307
rect 2338 1298 2481 1301
rect 2602 1298 2630 1301
rect 2778 1298 2798 1301
rect 2802 1298 2886 1301
rect 3546 1298 3558 1301
rect 3562 1298 3670 1301
rect 4162 1298 4334 1301
rect 4338 1298 4382 1301
rect 5066 1298 5134 1301
rect 5138 1298 5222 1301
rect 5234 1298 5254 1301
rect 242 1288 430 1291
rect 506 1288 566 1291
rect 826 1288 854 1291
rect 866 1288 886 1291
rect 1026 1288 1086 1291
rect 1090 1288 1206 1291
rect 1210 1288 1254 1291
rect 1258 1288 1598 1291
rect 1658 1288 2366 1291
rect 2474 1288 2478 1291
rect 2686 1288 2694 1291
rect 2698 1288 2782 1291
rect 3554 1288 3566 1291
rect 3570 1288 3590 1291
rect 3626 1288 3654 1291
rect 3738 1288 3798 1291
rect 3938 1288 3950 1291
rect 3962 1288 4094 1291
rect 4218 1288 4246 1291
rect 4318 1288 4326 1291
rect 4330 1288 4350 1291
rect 5026 1288 5158 1291
rect 5162 1288 5190 1291
rect 122 1278 286 1281
rect 290 1278 350 1281
rect 426 1278 454 1281
rect 458 1278 502 1281
rect 758 1281 761 1288
rect 758 1278 838 1281
rect 850 1278 894 1281
rect 898 1278 942 1281
rect 962 1278 966 1281
rect 994 1278 1022 1281
rect 1130 1278 1182 1281
rect 1186 1278 1214 1281
rect 1234 1278 1246 1281
rect 1346 1278 1350 1281
rect 1522 1278 1534 1281
rect 1538 1278 1545 1281
rect 1654 1281 1657 1288
rect 1554 1278 1657 1281
rect 1674 1278 1678 1281
rect 1738 1278 1766 1281
rect 1854 1278 1910 1281
rect 1986 1278 2054 1281
rect 2074 1278 2150 1281
rect 2178 1278 2182 1281
rect 2202 1278 2286 1281
rect 2314 1278 2326 1281
rect 2862 1281 2865 1288
rect 2826 1278 2865 1281
rect 2962 1278 2982 1281
rect 3102 1281 3105 1288
rect 2986 1278 3105 1281
rect 3262 1281 3265 1288
rect 3234 1278 3265 1281
rect 3394 1278 3462 1281
rect 3546 1278 3558 1281
rect 3690 1278 3702 1281
rect 3798 1281 3801 1288
rect 3798 1278 3894 1281
rect 3922 1278 4494 1281
rect 4514 1278 4646 1281
rect 4654 1281 4657 1288
rect 4654 1278 4774 1281
rect 4794 1278 4830 1281
rect 5018 1278 5062 1281
rect 5146 1278 5150 1281
rect 5226 1278 5238 1281
rect 5250 1278 5302 1281
rect 66 1268 94 1271
rect 98 1268 126 1271
rect 250 1268 414 1271
rect 418 1268 486 1271
rect 590 1271 593 1278
rect 1406 1272 1409 1278
rect 590 1268 614 1271
rect 730 1268 766 1271
rect 770 1268 830 1271
rect 834 1268 902 1271
rect 1058 1268 1062 1271
rect 1098 1268 1118 1271
rect 1122 1268 1134 1271
rect 1202 1268 1222 1271
rect 1298 1268 1310 1271
rect 1338 1268 1350 1271
rect 1474 1268 1558 1271
rect 1626 1268 1638 1271
rect 1666 1268 1678 1271
rect 1754 1268 1774 1271
rect 1778 1268 1782 1271
rect 1790 1271 1793 1278
rect 1838 1272 1841 1278
rect 1854 1272 1857 1278
rect 1790 1268 1822 1271
rect 1890 1268 1942 1271
rect 2058 1268 2086 1271
rect 2090 1268 2102 1271
rect 2114 1268 2126 1271
rect 2162 1268 2174 1271
rect 2258 1268 2294 1271
rect 2298 1268 2310 1271
rect 2498 1268 2670 1271
rect 2718 1271 2721 1278
rect 2718 1268 2758 1271
rect 2786 1268 2790 1271
rect 2882 1268 2910 1271
rect 2914 1268 2966 1271
rect 3042 1268 3054 1271
rect 3058 1268 3070 1271
rect 3082 1268 3158 1271
rect 3246 1268 3294 1271
rect 3314 1268 3358 1271
rect 3482 1268 3558 1271
rect 3618 1268 3638 1271
rect 3718 1271 3721 1278
rect 3658 1268 3721 1271
rect 4138 1268 4273 1271
rect 4314 1268 4342 1271
rect 4346 1268 4358 1271
rect 4642 1268 4662 1271
rect 4778 1268 4809 1271
rect 4938 1268 5006 1271
rect 5066 1268 5070 1271
rect 5178 1268 5198 1271
rect 5202 1268 5262 1271
rect 1606 1262 1609 1268
rect 34 1258 78 1261
rect 226 1258 273 1261
rect 330 1258 361 1261
rect 378 1258 414 1261
rect 418 1258 454 1261
rect 742 1258 777 1261
rect 786 1258 798 1261
rect 802 1258 806 1261
rect 834 1258 998 1261
rect 1002 1258 1222 1261
rect 1250 1258 1254 1261
rect 1306 1258 1326 1261
rect 1394 1258 1550 1261
rect 1586 1258 1606 1261
rect 1634 1258 1654 1261
rect 1706 1258 1710 1261
rect 1762 1258 1782 1261
rect 1786 1258 1790 1261
rect 1802 1258 1825 1261
rect 1882 1258 1910 1261
rect 1922 1259 1998 1261
rect 3246 1262 3249 1268
rect 2002 1259 2046 1261
rect 1922 1258 2046 1259
rect 2274 1258 2278 1261
rect 2282 1258 2302 1261
rect 2338 1258 2390 1261
rect 2618 1258 2718 1261
rect 2754 1258 2790 1261
rect 2794 1258 2814 1261
rect 2890 1258 2902 1261
rect 2906 1258 2942 1261
rect 3002 1258 3006 1261
rect 3050 1258 3094 1261
rect 3098 1258 3158 1261
rect 3390 1261 3393 1268
rect 3346 1258 3393 1261
rect 3402 1258 3406 1261
rect 3682 1258 3782 1261
rect 3894 1261 3897 1268
rect 4270 1262 4273 1268
rect 4806 1262 4809 1268
rect 3894 1258 3950 1261
rect 4202 1258 4246 1261
rect 4298 1258 4318 1261
rect 4358 1258 4366 1261
rect 4370 1258 4441 1261
rect 4522 1258 4718 1261
rect 4906 1258 5070 1261
rect 5074 1258 5081 1261
rect 5154 1258 5190 1261
rect 5242 1258 5246 1261
rect 270 1252 273 1258
rect 358 1252 361 1258
rect 42 1248 54 1251
rect 242 1248 262 1251
rect 274 1248 286 1251
rect 370 1248 710 1251
rect 734 1251 737 1258
rect 742 1252 745 1258
rect 774 1252 777 1258
rect 1822 1252 1825 1258
rect 2134 1252 2137 1258
rect 734 1248 742 1251
rect 866 1248 1006 1251
rect 1146 1248 1206 1251
rect 1322 1248 1334 1251
rect 1490 1248 1518 1251
rect 1546 1248 1606 1251
rect 1650 1248 1662 1251
rect 1762 1248 1766 1251
rect 1770 1248 1782 1251
rect 2050 1248 2086 1251
rect 2174 1251 2177 1258
rect 2558 1252 2561 1258
rect 2174 1248 2214 1251
rect 2314 1248 2406 1251
rect 2642 1248 2670 1251
rect 2850 1248 2889 1251
rect 2954 1248 2974 1251
rect 3022 1251 3025 1258
rect 4438 1252 4441 1258
rect 2978 1248 3025 1251
rect 3034 1248 3062 1251
rect 3498 1248 3502 1251
rect 3586 1248 3606 1251
rect 4578 1248 4582 1251
rect 4642 1248 4662 1251
rect 4754 1248 4782 1251
rect 4786 1248 4798 1251
rect 4834 1248 4838 1251
rect 4890 1248 4990 1251
rect 4994 1248 5054 1251
rect 5058 1248 5062 1251
rect 5066 1248 5174 1251
rect 5262 1248 5281 1251
rect 162 1238 262 1241
rect 266 1238 398 1241
rect 402 1238 486 1241
rect 610 1238 710 1241
rect 714 1238 750 1241
rect 826 1238 1590 1241
rect 1594 1238 1814 1241
rect 1818 1238 2254 1241
rect 2454 1241 2457 1248
rect 2886 1242 2889 1248
rect 5262 1242 5265 1248
rect 5278 1242 5281 1248
rect 2454 1238 2526 1241
rect 2754 1238 2790 1241
rect 2906 1238 3102 1241
rect 4850 1238 4902 1241
rect 5042 1238 5046 1241
rect 5066 1238 5070 1241
rect 5146 1238 5206 1241
rect 162 1228 238 1231
rect 338 1228 406 1231
rect 490 1228 614 1231
rect 618 1228 926 1231
rect 1074 1228 1078 1231
rect 1082 1228 1110 1231
rect 1154 1228 1174 1231
rect 1194 1228 1510 1231
rect 1514 1228 1694 1231
rect 1762 1228 1766 1231
rect 2090 1228 2222 1231
rect 2698 1228 2838 1231
rect 2842 1228 2854 1231
rect 3010 1228 3057 1231
rect 3530 1228 4553 1231
rect 4562 1228 4974 1231
rect 4978 1228 5054 1231
rect 5206 1231 5209 1238
rect 5206 1228 5270 1231
rect 258 1218 838 1221
rect 882 1218 1286 1221
rect 1294 1218 1478 1221
rect 1570 1218 1974 1221
rect 1978 1218 2342 1221
rect 2346 1218 2518 1221
rect 2778 1218 2782 1221
rect 2998 1221 3001 1228
rect 2786 1218 3001 1221
rect 3054 1222 3057 1228
rect 3386 1218 3622 1221
rect 3626 1218 3702 1221
rect 3706 1218 4062 1221
rect 4066 1218 4110 1221
rect 4550 1221 4553 1228
rect 4550 1218 4614 1221
rect 4618 1218 4878 1221
rect 5018 1218 5158 1221
rect 5162 1218 5230 1221
rect 5234 1218 5246 1221
rect 18 1208 46 1211
rect 50 1208 110 1211
rect 314 1208 334 1211
rect 674 1208 710 1211
rect 930 1208 966 1211
rect 1294 1211 1297 1218
rect 970 1208 1297 1211
rect 1898 1208 1958 1211
rect 2666 1208 2678 1211
rect 2682 1208 2702 1211
rect 2762 1208 2774 1211
rect 2778 1208 2918 1211
rect 2962 1208 3006 1211
rect 3338 1208 3390 1211
rect 5106 1208 5214 1211
rect 5218 1208 5222 1211
rect 344 1203 346 1207
rect 350 1203 353 1207
rect 358 1203 360 1207
rect 1368 1203 1370 1207
rect 1374 1203 1377 1207
rect 1382 1203 1384 1207
rect 2392 1203 2394 1207
rect 2398 1203 2401 1207
rect 2406 1203 2408 1207
rect 3416 1203 3418 1207
rect 3422 1203 3425 1207
rect 3430 1203 3432 1207
rect 4440 1203 4442 1207
rect 4446 1203 4449 1207
rect 4454 1203 4456 1207
rect 26 1198 38 1201
rect 218 1198 326 1201
rect 814 1198 990 1201
rect 994 1198 1030 1201
rect 1066 1198 1086 1201
rect 1090 1198 1198 1201
rect 1602 1198 2286 1201
rect 2874 1198 3094 1201
rect 3098 1198 3182 1201
rect 5210 1198 5222 1201
rect 814 1192 817 1198
rect 118 1188 126 1191
rect 130 1188 318 1191
rect 338 1188 462 1191
rect 578 1188 622 1191
rect 730 1188 814 1191
rect 906 1188 1094 1191
rect 1106 1188 1614 1191
rect 2026 1188 2030 1191
rect 2314 1188 2966 1191
rect 3202 1188 4014 1191
rect 4018 1188 4054 1191
rect 4506 1188 4574 1191
rect 4682 1188 5345 1191
rect 290 1178 318 1181
rect 322 1178 438 1181
rect 626 1178 934 1181
rect 1786 1178 1902 1181
rect 2074 1178 2142 1181
rect 2146 1178 2166 1181
rect 2426 1178 2470 1181
rect 2994 1178 3966 1181
rect 4098 1178 4198 1181
rect 4202 1178 4318 1181
rect 4322 1178 4430 1181
rect 4434 1178 4446 1181
rect 4502 1181 4505 1188
rect 5342 1182 5345 1188
rect 4450 1178 4505 1181
rect 5342 1178 5346 1182
rect 162 1168 174 1171
rect 218 1168 534 1171
rect 770 1168 806 1171
rect 826 1168 1142 1171
rect 1258 1168 1262 1171
rect 1598 1171 1601 1178
rect 1598 1168 1606 1171
rect 1610 1168 1646 1171
rect 1906 1168 2086 1171
rect 2098 1168 2190 1171
rect 2330 1168 2446 1171
rect 2450 1168 2478 1171
rect 2690 1168 2734 1171
rect 2906 1168 2966 1171
rect 2970 1168 2998 1171
rect 3002 1168 4102 1171
rect 4154 1168 4166 1171
rect 4234 1168 4238 1171
rect 4274 1168 4678 1171
rect 4818 1168 4902 1171
rect 5106 1168 5126 1171
rect 5246 1171 5249 1178
rect 5130 1168 5249 1171
rect 402 1158 406 1161
rect 418 1158 422 1161
rect 442 1158 510 1161
rect 742 1161 745 1168
rect 562 1158 745 1161
rect 794 1158 822 1161
rect 1218 1158 1238 1161
rect 1242 1158 1246 1161
rect 1498 1158 1502 1161
rect 1682 1158 1686 1161
rect 1810 1158 1830 1161
rect 1850 1158 1854 1161
rect 2042 1158 2054 1161
rect 2058 1158 2094 1161
rect 2154 1158 2198 1161
rect 2210 1158 2230 1161
rect 2234 1158 2270 1161
rect 2274 1158 2294 1161
rect 2298 1158 2502 1161
rect 2570 1158 2606 1161
rect 2686 1161 2689 1168
rect 2626 1158 2689 1161
rect 2962 1158 2990 1161
rect 3506 1158 3558 1161
rect 3562 1158 3590 1161
rect 3610 1158 3742 1161
rect 3746 1158 3774 1161
rect 4002 1158 4038 1161
rect 4242 1158 4294 1161
rect 4298 1158 4342 1161
rect 5122 1158 5142 1161
rect 5162 1158 5174 1161
rect 5178 1158 5182 1161
rect 5342 1161 5346 1162
rect 5314 1158 5346 1161
rect 98 1148 110 1151
rect 114 1148 134 1151
rect 166 1151 169 1158
rect 154 1148 169 1151
rect 178 1148 230 1151
rect 234 1148 462 1151
rect 546 1148 558 1151
rect 562 1148 598 1151
rect 646 1148 678 1151
rect 722 1148 742 1151
rect 746 1148 774 1151
rect 810 1148 830 1151
rect 962 1148 1022 1151
rect 1030 1151 1033 1158
rect 1030 1148 1286 1151
rect 1326 1148 1398 1151
rect 1614 1148 1670 1151
rect 1674 1148 1702 1151
rect 1990 1151 1993 1158
rect 1850 1148 1993 1151
rect 2042 1148 2110 1151
rect 2146 1148 2174 1151
rect 2274 1148 2342 1151
rect 2346 1148 2438 1151
rect 2822 1151 2825 1158
rect 2442 1148 2825 1151
rect 3198 1151 3201 1158
rect 2890 1148 3201 1151
rect 3398 1151 3401 1158
rect 4102 1152 4105 1158
rect 4742 1152 4745 1158
rect 3398 1148 3430 1151
rect 3462 1148 3470 1151
rect 3474 1148 3542 1151
rect 3546 1148 3582 1151
rect 3586 1148 3622 1151
rect 130 1138 190 1141
rect 194 1138 254 1141
rect 290 1138 302 1141
rect 358 1138 414 1141
rect 494 1141 497 1148
rect 646 1142 649 1148
rect 494 1138 574 1141
rect 698 1138 958 1141
rect 1018 1138 1233 1141
rect 1326 1141 1329 1148
rect 1290 1138 1329 1141
rect 1338 1138 1342 1141
rect 1446 1141 1449 1148
rect 1510 1141 1513 1148
rect 1614 1142 1617 1148
rect 3690 1148 3726 1151
rect 3834 1148 3865 1151
rect 3962 1148 3990 1151
rect 4122 1148 4206 1151
rect 4242 1148 4262 1151
rect 4306 1148 4334 1151
rect 4378 1148 4430 1151
rect 4946 1148 4982 1151
rect 5078 1148 5086 1151
rect 5090 1148 5150 1151
rect 5154 1148 5158 1151
rect 5194 1148 5209 1151
rect 3862 1142 3865 1148
rect 5206 1142 5209 1148
rect 1446 1138 1513 1141
rect 1594 1138 1614 1141
rect 1626 1138 1638 1141
rect 1642 1138 1662 1141
rect 1778 1138 1862 1141
rect 1866 1138 1910 1141
rect 1914 1138 1934 1141
rect 1946 1138 1966 1141
rect 1970 1138 1982 1141
rect 2058 1138 2110 1141
rect 2138 1138 2182 1141
rect 2186 1138 2302 1141
rect 2490 1138 2614 1141
rect 2634 1138 2646 1141
rect 2690 1138 2710 1141
rect 2738 1138 2766 1141
rect 2934 1138 2977 1141
rect 3090 1138 3134 1141
rect 3474 1138 3534 1141
rect 3978 1138 4006 1141
rect 4194 1138 4222 1141
rect 4226 1138 4262 1141
rect 4266 1138 4310 1141
rect 4314 1138 4382 1141
rect 5106 1138 5118 1141
rect 5122 1138 5158 1141
rect 358 1132 361 1138
rect 98 1128 166 1131
rect 170 1128 230 1131
rect 410 1128 422 1131
rect 426 1128 542 1131
rect 570 1128 574 1131
rect 582 1131 585 1138
rect 1230 1132 1233 1138
rect 2502 1132 2505 1138
rect 2934 1132 2937 1138
rect 2974 1132 2977 1138
rect 582 1128 702 1131
rect 746 1128 1073 1131
rect 270 1121 273 1128
rect 1070 1122 1073 1128
rect 1234 1128 1238 1131
rect 1242 1128 1302 1131
rect 1402 1128 1454 1131
rect 1466 1128 1798 1131
rect 1818 1128 1846 1131
rect 1938 1128 1961 1131
rect 1986 1128 1990 1131
rect 2034 1128 2038 1131
rect 2106 1128 2454 1131
rect 2610 1128 2630 1131
rect 2706 1128 2718 1131
rect 2722 1128 2750 1131
rect 2866 1128 2910 1131
rect 3466 1128 3494 1131
rect 3618 1128 3729 1131
rect 130 1118 273 1121
rect 530 1118 558 1121
rect 578 1118 758 1121
rect 762 1118 830 1121
rect 838 1118 878 1121
rect 954 1118 974 1121
rect 1182 1121 1185 1128
rect 1958 1122 1961 1128
rect 3726 1122 3729 1128
rect 3914 1128 3958 1131
rect 3962 1128 3998 1131
rect 4050 1128 4182 1131
rect 4210 1128 4230 1131
rect 4442 1128 4566 1131
rect 4758 1128 4814 1131
rect 4910 1131 4913 1138
rect 4910 1128 4966 1131
rect 1170 1118 1185 1121
rect 1394 1118 1422 1121
rect 1442 1118 1550 1121
rect 1794 1118 1798 1121
rect 1818 1118 1830 1121
rect 2114 1118 2254 1121
rect 2330 1118 2398 1121
rect 2458 1118 2478 1121
rect 2642 1118 2670 1121
rect 2674 1118 2726 1121
rect 2734 1118 2862 1121
rect 2866 1118 2982 1121
rect 3002 1118 3062 1121
rect 3482 1118 3502 1121
rect 3782 1121 3785 1128
rect 3738 1118 3785 1121
rect 4354 1118 4558 1121
rect 4758 1121 4761 1128
rect 4594 1118 4761 1121
rect 4770 1118 4886 1121
rect 4890 1118 4910 1121
rect 4914 1118 5030 1121
rect 186 1108 262 1111
rect 266 1108 310 1111
rect 314 1108 326 1111
rect 554 1108 662 1111
rect 838 1111 841 1118
rect 682 1108 841 1111
rect 1130 1108 1150 1111
rect 1458 1108 1654 1111
rect 1954 1108 1990 1111
rect 2002 1108 2014 1111
rect 2018 1108 2166 1111
rect 2266 1108 2382 1111
rect 2734 1111 2737 1118
rect 2674 1108 2737 1111
rect 2842 1108 2870 1111
rect 3362 1108 3406 1111
rect 3506 1108 3526 1111
rect 3530 1108 3574 1111
rect 3578 1108 3798 1111
rect 856 1103 858 1107
rect 862 1103 865 1107
rect 870 1103 872 1107
rect 1872 1103 1874 1107
rect 1878 1103 1881 1107
rect 1886 1103 1888 1107
rect 2904 1103 2906 1107
rect 2910 1103 2913 1107
rect 2918 1103 2920 1107
rect 3928 1103 3930 1107
rect 3934 1103 3937 1107
rect 3942 1103 3944 1107
rect 4622 1102 4625 1108
rect 4952 1103 4954 1107
rect 4958 1103 4961 1107
rect 4966 1103 4968 1107
rect 58 1098 374 1101
rect 522 1098 782 1101
rect 914 1098 942 1101
rect 946 1098 1094 1101
rect 1098 1098 1134 1101
rect 1138 1098 1158 1101
rect 1266 1098 1366 1101
rect 1530 1098 1558 1101
rect 1562 1098 1694 1101
rect 2130 1098 2158 1101
rect 2370 1098 2574 1101
rect 3450 1098 3582 1101
rect 3586 1098 3710 1101
rect 3714 1098 3846 1101
rect 3954 1098 4214 1101
rect 4218 1098 4582 1101
rect 86 1088 222 1091
rect 234 1088 278 1091
rect 286 1088 374 1091
rect 462 1088 470 1091
rect 474 1088 550 1091
rect 834 1088 1062 1091
rect 1138 1088 1430 1091
rect 1458 1088 1462 1091
rect 1634 1088 1654 1091
rect 1914 1088 2006 1091
rect 2058 1088 2142 1091
rect 2170 1088 2969 1091
rect 3186 1088 3310 1091
rect 3642 1088 3742 1091
rect 3746 1088 3830 1091
rect 3890 1088 3974 1091
rect 3978 1088 3990 1091
rect 4026 1088 4126 1091
rect 4130 1088 4206 1091
rect 4210 1088 4238 1091
rect 4242 1088 4326 1091
rect 4690 1088 5006 1091
rect 86 1082 89 1088
rect 74 1078 78 1081
rect 178 1078 214 1081
rect 286 1081 289 1088
rect 274 1078 289 1081
rect 378 1078 406 1081
rect 410 1078 478 1081
rect 482 1078 630 1081
rect 714 1078 734 1081
rect 970 1078 1014 1081
rect 1018 1078 1046 1081
rect 1050 1078 1102 1081
rect 1126 1081 1129 1088
rect 1126 1078 1230 1081
rect 1234 1078 1270 1081
rect 1550 1081 1553 1088
rect 1622 1081 1625 1088
rect 2966 1082 2969 1088
rect 1506 1078 1625 1081
rect 1650 1078 1742 1081
rect 1762 1078 1846 1081
rect 1970 1078 1974 1081
rect 1978 1078 1990 1081
rect 2178 1078 2214 1081
rect 2386 1078 2558 1081
rect 2562 1078 2598 1081
rect 2602 1078 2622 1081
rect 2778 1078 2806 1081
rect 2858 1078 2886 1081
rect 2890 1078 2926 1081
rect 3314 1078 3334 1081
rect 3338 1078 3406 1081
rect 3410 1078 3470 1081
rect 3562 1078 3614 1081
rect 3634 1078 3638 1081
rect 3666 1078 3678 1081
rect 3826 1078 3966 1081
rect 4026 1078 4070 1081
rect 4074 1078 4350 1081
rect 4478 1081 4481 1088
rect 4362 1078 4481 1081
rect 4502 1081 4505 1088
rect 4502 1078 4518 1081
rect 5266 1078 5281 1081
rect 5342 1081 5346 1082
rect 5314 1078 5346 1081
rect 150 1071 153 1078
rect 74 1068 174 1071
rect 282 1068 566 1071
rect 594 1068 598 1071
rect 610 1068 646 1071
rect 702 1071 705 1078
rect 650 1068 705 1071
rect 714 1068 742 1071
rect 826 1068 830 1071
rect 934 1068 1054 1071
rect 1098 1068 1150 1071
rect 1202 1068 1310 1071
rect 1314 1068 1342 1071
rect 1346 1068 1446 1071
rect 1450 1068 1574 1071
rect 1810 1068 1814 1071
rect 1858 1068 1942 1071
rect 1946 1068 1998 1071
rect 2142 1071 2145 1078
rect 2294 1072 2297 1078
rect 2142 1068 2190 1071
rect 2354 1068 2358 1071
rect 2498 1068 2526 1071
rect 2686 1070 2734 1071
rect 38 1061 41 1068
rect 62 1061 65 1068
rect 934 1062 937 1068
rect 38 1058 65 1061
rect 130 1058 142 1061
rect 290 1058 294 1061
rect 298 1058 382 1061
rect 394 1058 430 1061
rect 434 1058 470 1061
rect 474 1058 582 1061
rect 590 1058 630 1061
rect 746 1058 766 1061
rect 770 1058 926 1061
rect 1074 1058 1166 1061
rect 1202 1058 1214 1061
rect 1354 1058 1446 1061
rect 1554 1058 1582 1061
rect 1726 1058 1774 1061
rect 1830 1061 1833 1068
rect 2690 1068 2734 1070
rect 2738 1068 2742 1071
rect 2786 1068 2814 1071
rect 2818 1068 2942 1071
rect 3150 1071 3153 1078
rect 3150 1068 3214 1071
rect 3570 1068 3598 1071
rect 3626 1068 3734 1071
rect 3938 1068 4030 1071
rect 4498 1068 4550 1071
rect 4570 1068 4590 1071
rect 4662 1071 4665 1078
rect 5278 1072 5281 1078
rect 4594 1068 4665 1071
rect 5202 1068 5222 1071
rect 1830 1058 1846 1061
rect 1882 1058 1926 1061
rect 1930 1058 1942 1061
rect 1946 1058 1974 1061
rect 2074 1058 2134 1061
rect 2138 1058 2230 1061
rect 2270 1058 2310 1061
rect 2314 1058 2342 1061
rect 2386 1058 2438 1061
rect 2482 1058 2502 1061
rect 2506 1058 2542 1061
rect 2658 1058 2662 1061
rect 2754 1058 2838 1061
rect 2858 1058 2886 1061
rect 2922 1058 2950 1061
rect 3162 1058 3206 1061
rect 3430 1061 3433 1068
rect 4742 1062 4745 1068
rect 5078 1062 5081 1068
rect 3430 1058 3726 1061
rect 3758 1058 3886 1061
rect 3962 1058 4078 1061
rect 4114 1058 4153 1061
rect 4242 1058 4286 1061
rect 4378 1058 4390 1061
rect 4410 1058 4502 1061
rect 4834 1058 4862 1061
rect 4866 1058 4910 1061
rect 4922 1058 4942 1061
rect 4946 1058 4982 1061
rect 4986 1058 4990 1061
rect 5026 1058 5046 1061
rect 5342 1061 5346 1062
rect 5082 1058 5346 1061
rect 78 1051 81 1058
rect 66 1048 81 1051
rect 154 1048 190 1051
rect 506 1048 534 1051
rect 546 1048 558 1051
rect 590 1051 593 1058
rect 562 1048 593 1051
rect 726 1051 729 1058
rect 634 1048 729 1051
rect 746 1048 750 1051
rect 754 1048 934 1051
rect 994 1048 1030 1051
rect 1034 1048 1070 1051
rect 1114 1048 1142 1051
rect 1214 1048 1270 1051
rect 1274 1048 1286 1051
rect 1306 1048 1414 1051
rect 1470 1051 1473 1058
rect 1726 1052 1729 1058
rect 1426 1048 1510 1051
rect 1730 1048 1734 1051
rect 1842 1048 1910 1051
rect 1914 1048 1966 1051
rect 2166 1048 2174 1051
rect 2270 1051 2273 1058
rect 3758 1052 3761 1058
rect 4150 1052 4153 1058
rect 2178 1048 2273 1051
rect 2306 1048 2574 1051
rect 2578 1048 2606 1051
rect 2666 1048 2702 1051
rect 2746 1048 2769 1051
rect 2778 1048 2801 1051
rect 2842 1048 2854 1051
rect 2858 1048 2862 1051
rect 2890 1048 2982 1051
rect 3202 1048 3262 1051
rect 3650 1048 3702 1051
rect 4186 1048 4222 1051
rect 4290 1048 4350 1051
rect 4426 1048 4518 1051
rect 4574 1051 4577 1058
rect 4522 1048 4577 1051
rect 4918 1051 4921 1058
rect 4898 1048 4921 1051
rect 5154 1048 5254 1051
rect 34 1038 102 1041
rect 106 1038 246 1041
rect 450 1038 454 1041
rect 458 1038 542 1041
rect 626 1038 830 1041
rect 834 1038 950 1041
rect 958 1041 961 1048
rect 1214 1042 1217 1048
rect 958 1038 998 1041
rect 1002 1038 1030 1041
rect 1050 1038 1182 1041
rect 1434 1038 1606 1041
rect 1746 1038 2038 1041
rect 2042 1038 2214 1041
rect 2278 1041 2281 1048
rect 2766 1042 2769 1048
rect 2798 1042 2801 1048
rect 2274 1038 2281 1041
rect 2354 1038 2462 1041
rect 2466 1038 2550 1041
rect 2602 1038 2646 1041
rect 2818 1038 2934 1041
rect 3106 1038 3166 1041
rect 3170 1038 3198 1041
rect 3202 1038 3225 1041
rect 3498 1038 3654 1041
rect 3658 1038 3694 1041
rect 3698 1038 3710 1041
rect 3906 1038 4006 1041
rect 4010 1038 4022 1041
rect 4338 1038 4382 1041
rect 4398 1041 4401 1048
rect 4398 1038 4430 1041
rect 4658 1038 4670 1041
rect 4778 1038 5110 1041
rect 1486 1032 1489 1038
rect 3222 1032 3225 1038
rect 1018 1028 1118 1031
rect 1362 1028 1478 1031
rect 1602 1028 2942 1031
rect 3330 1028 3590 1031
rect 510 1022 513 1028
rect 538 1018 558 1021
rect 562 1018 686 1021
rect 714 1018 846 1021
rect 850 1018 1534 1021
rect 2170 1018 2190 1021
rect 2270 1018 2278 1021
rect 2282 1018 2326 1021
rect 2330 1018 2358 1021
rect 2362 1018 2494 1021
rect 2510 1018 2518 1021
rect 2522 1018 2582 1021
rect 2794 1018 2862 1021
rect 3234 1018 3318 1021
rect 3322 1018 3350 1021
rect 3578 1018 3774 1021
rect 3778 1018 3934 1021
rect 4322 1018 4414 1021
rect 442 1008 598 1011
rect 1498 1008 1510 1011
rect 1522 1008 1614 1011
rect 1618 1008 2102 1011
rect 2106 1008 2230 1011
rect 2362 1008 2382 1011
rect 3858 1008 3910 1011
rect 3994 1008 4062 1011
rect 4490 1008 4582 1011
rect 4586 1008 4606 1011
rect 5034 1008 5270 1011
rect 344 1003 346 1007
rect 350 1003 353 1007
rect 358 1003 360 1007
rect 1368 1003 1370 1007
rect 1374 1003 1377 1007
rect 1382 1003 1384 1007
rect 2392 1003 2394 1007
rect 2398 1003 2401 1007
rect 2406 1003 2408 1007
rect 3416 1003 3418 1007
rect 3422 1003 3425 1007
rect 3430 1003 3432 1007
rect 4440 1003 4442 1007
rect 4446 1003 4449 1007
rect 4454 1003 4456 1007
rect 386 998 518 1001
rect 1418 998 1462 1001
rect 1466 998 1590 1001
rect 2090 998 2318 1001
rect 2746 998 3110 1001
rect 130 988 1134 991
rect 1306 988 1310 991
rect 1314 988 1406 991
rect 1482 988 1537 991
rect 1554 988 1718 991
rect 2322 988 2734 991
rect 3730 988 3990 991
rect 3994 988 4142 991
rect 4146 988 4238 991
rect 4642 988 4857 991
rect 1534 982 1537 988
rect 170 978 198 981
rect 306 978 478 981
rect 846 978 1030 981
rect 1234 978 1430 981
rect 1434 978 1462 981
rect 1538 978 1702 981
rect 1706 978 1750 981
rect 2170 978 2478 981
rect 2962 978 3126 981
rect 3694 981 3697 988
rect 4854 982 4857 988
rect 3694 978 4118 981
rect 4122 978 4254 981
rect 4618 978 4710 981
rect 82 968 246 971
rect 250 968 406 971
rect 418 968 470 971
rect 514 968 518 971
rect 630 971 633 978
rect 846 972 849 978
rect 630 968 646 971
rect 954 968 958 971
rect 978 968 998 971
rect 1050 968 1094 971
rect 1322 968 1566 971
rect 1758 971 1761 978
rect 1578 968 1761 971
rect 2234 968 2342 971
rect 2370 968 2374 971
rect 2546 968 2798 971
rect 2802 968 2870 971
rect 3162 968 3182 971
rect 3370 968 3478 971
rect 3482 968 3614 971
rect 3618 968 3630 971
rect 3650 968 3774 971
rect 3806 968 3822 971
rect 3826 968 3846 971
rect 3858 968 3982 971
rect 3986 968 4022 971
rect 4026 968 4134 971
rect 4322 968 4390 971
rect 4546 968 4574 971
rect 4578 968 4753 971
rect 5098 968 5206 971
rect 5210 968 5238 971
rect 146 958 182 961
rect 202 958 366 961
rect 402 958 438 961
rect 554 958 574 961
rect 678 961 681 968
rect 618 958 681 961
rect 842 958 918 961
rect 922 958 974 961
rect 1014 961 1017 968
rect 1014 958 1086 961
rect 1210 958 1366 961
rect 1526 958 1534 961
rect 1538 958 1542 961
rect 1610 958 1686 961
rect 1722 958 1838 961
rect 2130 958 2142 961
rect 2330 958 2390 961
rect 2466 958 2494 961
rect 2514 958 2678 961
rect 2990 961 2993 968
rect 3806 962 3809 968
rect 4750 962 4753 968
rect 2682 958 2993 961
rect 3154 958 3422 961
rect 3674 958 3806 961
rect 3818 958 3830 961
rect 4402 958 4478 961
rect 4482 958 4654 961
rect 4890 958 4942 961
rect 5242 958 5254 961
rect 510 952 513 958
rect 798 952 801 958
rect 162 948 222 951
rect 546 948 566 951
rect 586 948 638 951
rect 642 948 718 951
rect 930 948 934 951
rect 946 948 966 951
rect 1034 948 1038 951
rect 1066 948 1094 951
rect 1138 948 1174 951
rect 1178 948 1230 951
rect 1374 951 1377 958
rect 1374 948 1390 951
rect 1394 948 1422 951
rect 1438 948 1454 951
rect 1494 951 1497 958
rect 1494 948 1518 951
rect 1690 948 1702 951
rect 1706 948 1734 951
rect 1850 948 1886 951
rect 2022 951 2025 958
rect 2022 948 2030 951
rect 2098 948 2134 951
rect 2214 948 2278 951
rect 2282 948 2334 951
rect 2346 948 2534 951
rect 2538 948 2542 951
rect 2562 948 2606 951
rect 2610 948 2614 951
rect 2626 948 2654 951
rect 2822 948 2974 951
rect 3054 948 3086 951
rect 3138 948 3182 951
rect 3186 948 3214 951
rect 3234 948 3238 951
rect 3298 948 3382 951
rect 3530 948 3590 951
rect 3618 948 3718 951
rect 3762 948 3862 951
rect 3882 948 3894 951
rect 3898 948 3958 951
rect 4150 951 4153 958
rect 4042 948 4153 951
rect 4170 948 4214 951
rect 4342 951 4345 958
rect 4342 948 4438 951
rect 4474 948 4502 951
rect 4522 948 4614 951
rect 4666 948 4678 951
rect 4698 948 4718 951
rect 4786 948 4934 951
rect 4986 948 5062 951
rect 5194 948 5198 951
rect 5342 951 5346 952
rect 5314 948 5346 951
rect 202 938 278 941
rect 414 941 417 948
rect 1438 942 1441 948
rect 2214 942 2217 948
rect 414 938 454 941
rect 530 938 550 941
rect 666 938 678 941
rect 842 938 846 941
rect 906 938 990 941
rect 1042 938 1110 941
rect 1114 938 1142 941
rect 1146 938 1254 941
rect 1274 938 1414 941
rect 1450 938 1574 941
rect 1618 938 1622 941
rect 1786 938 1870 941
rect 1874 938 1934 941
rect 2106 938 2118 941
rect 2122 938 2174 941
rect 2338 938 2342 941
rect 2362 938 2414 941
rect 2418 938 2430 941
rect 2498 938 2518 941
rect 2558 941 2561 948
rect 2546 938 2561 941
rect 2710 942 2713 948
rect 2822 942 2825 948
rect 2974 941 2977 948
rect 3054 942 3057 948
rect 3470 942 3473 948
rect 4222 942 4225 948
rect 2974 938 3046 941
rect 3154 938 3198 941
rect 3498 938 3590 941
rect 3594 938 3622 941
rect 3794 938 3886 941
rect 3890 938 3950 941
rect 3978 938 3998 941
rect 4098 938 4118 941
rect 4138 938 4182 941
rect 4370 938 4385 941
rect 4394 938 4494 941
rect 4570 938 4686 941
rect 4690 938 4742 941
rect 4802 938 4862 941
rect 4874 938 4886 941
rect 4986 938 5046 941
rect 5062 941 5065 948
rect 5126 941 5129 948
rect 5062 938 5129 941
rect 5278 941 5281 948
rect 5234 938 5281 941
rect 226 928 286 931
rect 390 931 393 938
rect 1078 932 1081 938
rect 290 928 393 931
rect 402 928 422 931
rect 426 928 534 931
rect 1514 928 1558 931
rect 1586 928 1606 931
rect 1626 928 1670 931
rect 1762 928 1790 931
rect 1802 928 2054 931
rect 2082 928 2094 931
rect 2262 931 2265 938
rect 2262 928 2438 931
rect 2442 928 2470 931
rect 2490 928 2614 931
rect 2754 928 2758 931
rect 3010 928 3094 931
rect 3098 928 3118 931
rect 3122 928 3142 931
rect 3270 931 3273 938
rect 4382 932 4385 938
rect 4846 932 4849 938
rect 3146 928 3286 931
rect 3506 928 3534 931
rect 3538 928 3726 931
rect 4034 928 4046 931
rect 4130 928 4166 931
rect 4186 928 4190 931
rect 4194 928 4222 931
rect 4306 928 4318 931
rect 4602 928 4630 931
rect 4650 928 4705 931
rect 4970 928 5006 931
rect 5050 928 5070 931
rect 5074 928 5142 931
rect 5178 928 5262 931
rect 274 918 390 921
rect 558 921 561 928
rect 450 918 561 921
rect 1106 918 1246 921
rect 1270 921 1273 928
rect 1470 922 1473 928
rect 1270 918 1422 921
rect 1490 918 1654 921
rect 1658 918 1726 921
rect 1818 918 1966 921
rect 1970 918 2054 921
rect 2074 918 2086 921
rect 2266 918 2462 921
rect 2622 921 2625 928
rect 2610 918 2625 921
rect 2866 918 2870 921
rect 3138 918 3254 921
rect 3258 918 3334 921
rect 3462 921 3465 928
rect 4702 922 4705 928
rect 3394 918 3510 921
rect 3946 918 4174 921
rect 4258 918 4278 921
rect 4546 918 4670 921
rect 4730 918 4790 921
rect 4794 918 4870 921
rect 4890 918 4974 921
rect 5114 918 5118 921
rect 5122 918 5174 921
rect 490 908 502 911
rect 506 908 670 911
rect 1138 908 1145 911
rect 1154 908 1158 911
rect 1170 908 1198 911
rect 1242 908 1278 911
rect 1282 908 1326 911
rect 1922 908 2081 911
rect 2098 908 2286 911
rect 2362 908 2582 911
rect 2626 908 2742 911
rect 2746 908 2870 911
rect 2970 908 3022 911
rect 3522 908 3566 911
rect 4130 908 4302 911
rect 4738 908 4745 911
rect 4770 908 4878 911
rect 856 903 858 907
rect 862 903 865 907
rect 870 903 872 907
rect 474 898 614 901
rect 1098 898 1134 901
rect 1142 901 1145 908
rect 1872 903 1874 907
rect 1878 903 1881 907
rect 1886 903 1888 907
rect 2078 902 2081 908
rect 2904 903 2906 907
rect 2910 903 2913 907
rect 2918 903 2920 907
rect 3928 903 3930 907
rect 3934 903 3937 907
rect 3942 903 3944 907
rect 1142 898 1150 901
rect 1226 898 1302 901
rect 1730 898 1774 901
rect 1778 898 1846 901
rect 2058 898 2062 901
rect 2138 898 2294 901
rect 2298 898 2366 901
rect 2410 898 2430 901
rect 2434 898 2582 901
rect 2586 898 2614 901
rect 3234 898 3262 901
rect 3266 898 3286 901
rect 3330 898 3342 901
rect 3426 898 3518 901
rect 3522 898 3542 901
rect 3642 898 3718 901
rect 3970 898 4078 901
rect 4082 898 4126 901
rect 4722 898 4734 901
rect 4742 901 4745 908
rect 4952 903 4954 907
rect 4958 903 4961 907
rect 4966 903 4968 907
rect 4742 898 4822 901
rect 114 888 206 891
rect 210 888 214 891
rect 446 891 449 898
rect 734 892 737 898
rect 446 888 542 891
rect 674 888 718 891
rect 754 888 774 891
rect 778 888 1358 891
rect 1394 888 1662 891
rect 1882 888 1945 891
rect 1954 888 2110 891
rect 2194 888 2649 891
rect 2730 888 2774 891
rect 2898 888 3030 891
rect 3042 888 3054 891
rect 3210 888 3358 891
rect 3470 888 3478 891
rect 3482 888 3494 891
rect 3874 888 3966 891
rect 4714 888 4814 891
rect 4938 888 5030 891
rect 5178 888 5206 891
rect 5226 888 5262 891
rect 550 882 553 888
rect 558 882 561 888
rect -26 881 -22 882
rect -26 878 6 881
rect 266 878 302 881
rect 338 878 406 881
rect 410 878 446 881
rect 506 878 542 881
rect 610 878 654 881
rect 658 878 710 881
rect 714 878 734 881
rect 866 878 918 881
rect 922 878 966 881
rect 1082 878 1126 881
rect 1138 878 1214 881
rect 1230 878 1238 881
rect 1242 878 1262 881
rect 1306 878 1318 881
rect 1514 878 1902 881
rect 1906 878 1926 881
rect 1942 881 1945 888
rect 2646 882 2649 888
rect 1942 878 1974 881
rect 2146 878 2182 881
rect 2186 878 2214 881
rect 2418 878 2446 881
rect 2450 878 2558 881
rect 2570 878 2598 881
rect 2834 878 2974 881
rect 3026 878 3030 881
rect 3078 881 3081 888
rect 3042 878 3081 881
rect 3162 878 3382 881
rect 3402 878 3430 881
rect 3434 878 3454 881
rect 3458 878 3478 881
rect 3510 881 3513 888
rect 3510 878 3614 881
rect 3698 878 3734 881
rect 3842 878 3881 881
rect 4038 881 4041 888
rect 3994 878 4041 881
rect 4058 878 4126 881
rect 4130 878 4206 881
rect 4466 878 4478 881
rect 4658 878 4702 881
rect 4706 878 4718 881
rect 4750 878 4766 881
rect 66 868 158 871
rect 278 868 297 871
rect 394 868 494 871
rect 498 868 638 871
rect 946 868 958 871
rect 962 868 977 871
rect -26 861 -22 862
rect -26 858 126 861
rect 158 861 161 868
rect 278 862 281 868
rect 294 862 297 868
rect 974 862 977 868
rect 1038 868 1166 871
rect 1198 868 1238 871
rect 1250 868 1262 871
rect 1278 871 1281 878
rect 1414 872 1417 878
rect 1278 868 1342 871
rect 1546 868 1609 871
rect 1666 868 1769 871
rect 1994 868 2030 871
rect 2170 868 2182 871
rect 2222 871 2225 878
rect 2638 872 2641 878
rect 2190 868 2225 871
rect 2298 868 2350 871
rect 2370 868 2494 871
rect 2522 868 2542 871
rect 2586 868 2590 871
rect 2834 868 2942 871
rect 2978 868 3078 871
rect 3082 868 3110 871
rect 3118 868 3121 878
rect 3126 871 3129 878
rect 3766 872 3769 878
rect 3126 868 3222 871
rect 3346 868 3430 871
rect 3482 868 3486 871
rect 3722 868 3766 871
rect 3858 868 3870 871
rect 3878 871 3881 878
rect 3878 868 3886 871
rect 4042 868 4054 871
rect 4410 868 4630 871
rect 4634 868 4654 871
rect 4750 871 4753 878
rect 5302 872 5305 878
rect 4698 868 4753 871
rect 4762 868 4774 871
rect 4866 868 4902 871
rect 4906 868 4934 871
rect 5050 868 5054 871
rect 5250 868 5270 871
rect 1038 862 1041 868
rect 1198 862 1201 868
rect 1606 862 1609 868
rect 1766 862 1769 868
rect 158 858 278 861
rect 306 858 534 861
rect 594 858 646 861
rect 698 858 734 861
rect 738 858 790 861
rect 994 858 1038 861
rect 1058 858 1078 861
rect 1130 858 1158 861
rect 1162 858 1174 861
rect 1234 858 1254 861
rect 1506 858 1550 861
rect 1610 858 1758 861
rect 1802 858 1806 861
rect 1810 858 1910 861
rect 1994 858 1998 861
rect 2018 858 2094 861
rect 2130 858 2142 861
rect 2190 861 2193 868
rect 2146 858 2193 861
rect 2218 858 2254 861
rect 2258 858 2342 861
rect 2386 858 2390 861
rect 2398 858 2422 861
rect 2426 858 2438 861
rect 2466 858 2470 861
rect 2526 858 2566 861
rect 2710 861 2713 868
rect 2710 858 2793 861
rect 2950 858 2958 861
rect 2962 858 3158 861
rect 3226 858 3254 861
rect 3258 858 3294 861
rect 3322 858 3326 861
rect 3466 858 3470 861
rect 3474 858 3662 861
rect 3794 858 3862 861
rect 4022 861 4025 868
rect 3922 858 4025 861
rect 4070 861 4073 868
rect 4070 858 4102 861
rect 4254 861 4257 868
rect 4186 858 4257 861
rect 4482 858 4510 861
rect 4514 858 4566 861
rect 4570 858 4606 861
rect 4850 858 4894 861
rect 5018 858 5070 861
rect 5130 858 5262 861
rect 5282 858 5302 861
rect 602 848 622 851
rect 626 848 686 851
rect 858 848 886 851
rect 890 848 918 851
rect 922 848 950 851
rect 954 848 958 851
rect 1050 848 1094 851
rect 1134 848 1294 851
rect 1306 848 1310 851
rect 1382 851 1385 858
rect 1382 848 1542 851
rect 1562 848 1630 851
rect 1850 848 1974 851
rect 1978 848 2006 851
rect 2042 848 2046 851
rect 2146 848 2150 851
rect 2162 848 2166 851
rect 2398 851 2401 858
rect 2526 852 2529 858
rect 2790 852 2793 858
rect 2338 848 2401 851
rect 2426 848 2454 851
rect 2458 848 2526 851
rect 2994 848 3038 851
rect 3058 848 3302 851
rect 3314 848 3630 851
rect 3690 848 3694 851
rect 3962 848 4062 851
rect 4338 848 4358 851
rect 4362 848 4398 851
rect 4530 848 4582 851
rect 4586 848 4606 851
rect 4794 848 4830 851
rect 4834 848 4846 851
rect 4882 848 4910 851
rect 4918 851 4921 858
rect 5030 852 5033 858
rect 4918 848 5006 851
rect 5010 848 5014 851
rect 362 838 614 841
rect 618 838 662 841
rect 1022 841 1025 848
rect 1134 842 1137 848
rect 1022 838 1086 841
rect 1090 838 1110 841
rect 1162 838 1342 841
rect 1610 838 1646 841
rect 1746 838 1870 841
rect 1898 838 1902 841
rect 2146 838 2158 841
rect 2274 838 2286 841
rect 2314 838 2414 841
rect 2818 838 3134 841
rect 3154 838 3278 841
rect 3282 838 3342 841
rect 3842 838 3854 841
rect 3858 838 3934 841
rect 3938 838 4086 841
rect 4378 838 4414 841
rect 4418 838 4534 841
rect 4546 838 4622 841
rect 4898 838 4926 841
rect 4994 838 5030 841
rect 1010 828 1057 831
rect 1082 828 1166 831
rect 1326 828 1334 831
rect 1338 828 1438 831
rect 1658 828 1742 831
rect 1794 828 1966 831
rect 2042 828 2046 831
rect 2058 828 2766 831
rect 2770 828 2926 831
rect 3106 828 3278 831
rect 3330 828 3374 831
rect 3698 828 4262 831
rect 4266 828 4318 831
rect 4434 828 4646 831
rect 4842 828 4950 831
rect 642 818 1046 821
rect 1054 821 1057 828
rect 1054 818 1094 821
rect 1254 821 1257 828
rect 1254 818 1430 821
rect 2274 818 2278 821
rect 2298 818 2358 821
rect 2618 818 3054 821
rect 3098 818 3326 821
rect 3578 818 3742 821
rect 3746 818 4422 821
rect 4426 818 4574 821
rect 4610 818 4686 821
rect 4690 818 4710 821
rect 4874 818 4982 821
rect 1010 808 1230 811
rect 1234 808 1238 811
rect 1954 808 2222 811
rect 3618 808 4126 811
rect 4274 808 4294 811
rect 4298 808 4334 811
rect 4370 808 4390 811
rect 4570 808 4702 811
rect 344 803 346 807
rect 350 803 353 807
rect 358 803 360 807
rect 1368 803 1370 807
rect 1374 803 1377 807
rect 1382 803 1384 807
rect 2392 803 2394 807
rect 2398 803 2401 807
rect 2406 803 2408 807
rect 3416 803 3418 807
rect 3422 803 3425 807
rect 3430 803 3432 807
rect 4440 803 4442 807
rect 4446 803 4449 807
rect 4454 803 4456 807
rect 1018 798 1142 801
rect 1314 798 1358 801
rect 1434 798 1446 801
rect 1834 798 2006 801
rect 2010 798 2022 801
rect 2450 798 2926 801
rect 2930 798 2934 801
rect 2946 798 3118 801
rect 3122 798 3353 801
rect 3642 798 3726 801
rect 4466 798 4766 801
rect 4770 798 5230 801
rect 3350 792 3353 798
rect 830 788 1710 791
rect 1866 788 2886 791
rect 2914 788 3214 791
rect 3354 788 3366 791
rect 3370 788 3454 791
rect 3722 788 3734 791
rect 5018 788 5134 791
rect 830 782 833 788
rect 298 778 830 781
rect 1046 778 1718 781
rect 1722 778 1926 781
rect 1938 778 1961 781
rect 2298 778 2502 781
rect 2778 778 4454 781
rect 4458 778 4478 781
rect 4514 778 4558 781
rect 4670 778 4678 781
rect 4682 778 4798 781
rect 5114 778 5182 781
rect 418 768 454 771
rect 470 768 478 771
rect 482 768 486 771
rect 1046 771 1049 778
rect 1958 772 1961 778
rect 690 768 1049 771
rect 1058 768 1126 771
rect 1154 768 1166 771
rect 1458 768 1462 771
rect 1506 768 1510 771
rect 1530 768 1534 771
rect 1542 768 1550 771
rect 1554 768 1574 771
rect 1730 768 1862 771
rect 2042 768 2062 771
rect 2138 768 2286 771
rect 2290 768 2326 771
rect 2482 768 2670 771
rect 3430 768 3470 771
rect 3746 768 3822 771
rect 4298 768 4310 771
rect 4322 768 4414 771
rect 4498 768 4582 771
rect 4610 768 4617 771
rect 4634 768 4670 771
rect 4674 768 4678 771
rect 4818 768 4974 771
rect 5022 771 5025 778
rect 4978 768 5025 771
rect 5146 768 5150 771
rect 210 758 238 761
rect 274 758 502 761
rect 522 758 553 761
rect 550 752 553 758
rect 1122 758 1182 761
rect 1342 761 1345 768
rect 1342 758 1406 761
rect 1410 758 1478 761
rect 1482 758 1510 761
rect 1518 761 1521 768
rect 1518 758 1542 761
rect 1794 758 1910 761
rect 1914 758 1926 761
rect 1950 761 1953 768
rect 1950 758 2078 761
rect 2082 758 2110 761
rect 2242 758 2246 761
rect 2250 758 2270 761
rect 2442 758 2470 761
rect 2538 758 2606 761
rect 3034 758 3054 761
rect 3066 758 3198 761
rect 3310 761 3313 768
rect 3430 762 3433 768
rect 3202 758 3390 761
rect 3394 758 3430 761
rect 3502 761 3505 768
rect 3466 758 3505 761
rect 3562 758 3662 761
rect 3666 758 3678 761
rect 3706 758 3726 761
rect 4066 758 4102 761
rect 4282 758 4342 761
rect 4346 758 4374 761
rect 4398 758 4406 761
rect 4410 758 4430 761
rect 4494 761 4497 768
rect 4614 762 4617 768
rect 4450 758 4497 761
rect 4538 758 4558 761
rect 4574 758 4606 761
rect 4642 758 4694 761
rect 4986 758 4998 761
rect 5082 758 5094 761
rect 5098 758 5102 761
rect 5130 758 5150 761
rect 798 752 801 758
rect -26 751 -22 752
rect -26 748 6 751
rect 10 748 38 751
rect 114 748 126 751
rect 186 748 217 751
rect 226 748 230 751
rect 330 748 342 751
rect 346 748 374 751
rect 442 748 510 751
rect 594 748 718 751
rect 818 748 1014 751
rect 1050 748 1150 751
rect 1262 751 1265 758
rect 4198 752 4201 758
rect 4574 752 4577 758
rect 1262 748 1270 751
rect 1314 748 1374 751
rect 1450 748 1454 751
rect 1474 748 1478 751
rect 1490 748 1558 751
rect 1578 748 1590 751
rect 1690 748 1814 751
rect 2090 748 2182 751
rect 2186 748 2206 751
rect 2322 748 2350 751
rect 2434 748 2462 751
rect 2466 748 2694 751
rect 2722 748 2790 751
rect 2906 748 3102 751
rect 3138 748 3166 751
rect 3190 748 3233 751
rect 3338 748 3382 751
rect 3386 748 3414 751
rect 3418 748 3446 751
rect 3450 748 3454 751
rect 3514 748 3526 751
rect 3642 748 3710 751
rect 3842 748 3870 751
rect 3874 748 3902 751
rect 4290 748 4318 751
rect 4386 748 4390 751
rect 4470 748 4486 751
rect 4490 748 4518 751
rect 4638 751 4641 758
rect 4638 748 4654 751
rect 4682 748 4734 751
rect 4790 751 4793 758
rect 4738 748 4793 751
rect 4858 748 4910 751
rect 4982 751 4985 758
rect 4930 748 4985 751
rect 5114 748 5129 751
rect 5202 748 5206 751
rect 5342 751 5346 752
rect 5210 748 5346 751
rect 214 742 217 748
rect 154 738 174 741
rect 318 738 334 741
rect 354 738 593 741
rect 318 732 321 738
rect 590 732 593 738
rect 666 738 710 741
rect 714 738 950 741
rect 1146 738 1174 741
rect 1186 738 1302 741
rect 1306 738 1334 741
rect 1366 738 1542 741
rect 1546 738 1582 741
rect 1662 741 1665 748
rect 1590 738 1665 741
rect 1714 738 2230 741
rect 2282 738 2310 741
rect 2370 738 2374 741
rect 2458 738 2646 741
rect 2838 741 2841 748
rect 2666 738 2841 741
rect 3110 741 3113 748
rect 3190 742 3193 748
rect 3230 742 3233 748
rect 4022 742 4025 748
rect 4470 742 4473 748
rect 5126 742 5129 748
rect 3058 738 3113 741
rect 3154 738 3158 741
rect 3282 738 3310 741
rect 3378 738 3398 741
rect 3522 738 3526 741
rect 4002 738 4022 741
rect 4106 738 4150 741
rect 4374 738 4398 741
rect 4482 738 4510 741
rect 4570 738 4614 741
rect 4618 738 4646 741
rect 4650 738 4710 741
rect 4714 738 4782 741
rect 4874 738 4942 741
rect 5170 738 5249 741
rect 654 732 657 738
rect 1030 732 1033 738
rect 1366 732 1369 738
rect 1590 732 1593 738
rect 1806 732 1809 738
rect 378 728 430 731
rect 450 728 478 731
rect 506 728 526 731
rect 554 728 558 731
rect 794 728 870 731
rect 874 728 990 731
rect 1090 728 1206 731
rect 1322 728 1326 731
rect 1386 728 1414 731
rect 1442 728 1446 731
rect 1482 728 1486 731
rect 1490 728 1494 731
rect 1602 728 1614 731
rect 1906 728 2070 731
rect 2114 728 2158 731
rect 2186 728 2238 731
rect 2258 728 2438 731
rect 2446 731 2449 738
rect 2442 728 2449 731
rect 2454 732 2457 738
rect 2466 728 2470 731
rect 2506 728 2510 731
rect 2622 728 2726 731
rect 2786 728 2934 731
rect 3130 728 3142 731
rect 3330 728 3398 731
rect 3402 728 3430 731
rect 3454 731 3457 738
rect 3582 732 3585 738
rect 4126 732 4129 738
rect 4374 732 4377 738
rect 5246 732 5249 738
rect 3454 728 3478 731
rect 4802 728 5038 731
rect 5042 728 5078 731
rect 94 718 206 721
rect 242 718 438 721
rect 534 721 537 728
rect 1470 722 1473 728
rect 534 718 558 721
rect 570 718 598 721
rect 602 718 630 721
rect 634 718 662 721
rect 930 718 982 721
rect 1018 718 1318 721
rect 1626 718 1686 721
rect 1850 718 1854 721
rect 1890 718 1918 721
rect 2090 718 2150 721
rect 2218 718 2318 721
rect 2378 718 2510 721
rect 2622 721 2625 728
rect 2586 718 2625 721
rect 2634 718 2766 721
rect 2818 718 2830 721
rect 3090 718 3254 721
rect 3266 718 3350 721
rect 3926 721 3929 728
rect 3926 718 3966 721
rect 4866 718 4926 721
rect 4946 718 5158 721
rect 94 712 97 718
rect 178 708 190 711
rect 194 708 278 711
rect 338 708 550 711
rect 922 708 934 711
rect 954 708 1502 711
rect 1578 708 1862 711
rect 2186 708 2214 711
rect 2426 708 2430 711
rect 2554 708 2729 711
rect 2762 708 2806 711
rect 2818 708 2854 711
rect 3130 708 3574 711
rect 3778 708 3814 711
rect 5034 708 5046 711
rect 856 703 858 707
rect 862 703 865 707
rect 870 703 872 707
rect 1872 703 1874 707
rect 1878 703 1881 707
rect 1886 703 1888 707
rect 2726 702 2729 708
rect 2904 703 2906 707
rect 2910 703 2913 707
rect 2918 703 2920 707
rect 3928 703 3930 707
rect 3934 703 3937 707
rect 3942 703 3944 707
rect 4952 703 4954 707
rect 4958 703 4961 707
rect 4966 703 4968 707
rect 234 698 254 701
rect 266 698 358 701
rect 450 698 782 701
rect 786 698 806 701
rect 906 698 1014 701
rect 1026 698 1134 701
rect 1170 698 1774 701
rect 2178 698 2302 701
rect 2466 698 2502 701
rect 2514 698 2590 701
rect 2618 698 2622 701
rect 2626 698 2630 701
rect 2642 698 2718 701
rect 2730 698 2822 701
rect 2970 698 3150 701
rect 3162 698 3254 701
rect 3482 698 3510 701
rect 4170 698 4198 701
rect 4202 698 4230 701
rect 4314 698 4342 701
rect 4426 698 4550 701
rect 4554 698 4766 701
rect 146 688 446 691
rect 546 688 926 691
rect 946 688 1030 691
rect 1074 688 1078 691
rect 1098 688 1150 691
rect 1250 688 1294 691
rect 1306 688 1366 691
rect 1370 688 1606 691
rect 1754 688 2030 691
rect 2034 688 2046 691
rect 2106 688 2118 691
rect 2290 688 2350 691
rect 2354 688 2438 691
rect 2442 688 2486 691
rect 2490 688 2662 691
rect 2670 688 2678 691
rect 2722 688 2782 691
rect 2794 688 2838 691
rect 3058 688 3166 691
rect 3178 688 3302 691
rect 3858 688 4073 691
rect 4154 688 4238 691
rect 4266 688 4486 691
rect 4490 688 4502 691
rect 4730 688 4750 691
rect 5210 688 5254 691
rect 4070 682 4073 688
rect 210 678 262 681
rect 266 678 302 681
rect 358 678 390 681
rect 410 678 470 681
rect 498 678 654 681
rect 874 678 1006 681
rect 1022 678 1310 681
rect 2322 678 2529 681
rect 2610 678 2654 681
rect 2658 678 2782 681
rect 2786 678 2798 681
rect 2866 678 2942 681
rect 3746 678 3774 681
rect 3778 678 3806 681
rect 3890 678 3974 681
rect 3978 678 3998 681
rect 4186 678 4486 681
rect 5086 681 5089 688
rect 5050 678 5089 681
rect 5106 678 5118 681
rect 5146 678 5254 681
rect 5342 681 5346 682
rect 5258 678 5346 681
rect 166 671 169 678
rect 358 672 361 678
rect 138 668 169 671
rect 186 668 190 671
rect 202 668 238 671
rect 254 668 294 671
rect 298 668 310 671
rect 330 668 358 671
rect 386 668 390 671
rect 402 668 518 671
rect 538 668 566 671
rect 702 671 705 678
rect 1022 672 1025 678
rect 1502 672 1505 678
rect 586 668 705 671
rect 842 668 950 671
rect 1042 668 1254 671
rect 1566 668 1614 671
rect 1618 668 1662 671
rect 1726 671 1729 678
rect 1674 668 1729 671
rect 1830 672 1833 678
rect 1866 668 1902 671
rect 2078 671 2081 678
rect 2030 668 2081 671
rect 2282 668 2342 671
rect 2346 668 2430 671
rect 2434 668 2481 671
rect 2490 668 2510 671
rect 2526 671 2529 678
rect 2526 668 2670 671
rect 2674 668 2686 671
rect 2722 668 2734 671
rect 2770 668 2886 671
rect 3086 671 3089 678
rect 3034 668 3089 671
rect 3214 672 3217 678
rect 3738 668 3766 671
rect 3770 668 3782 671
rect 3906 668 3958 671
rect 3970 668 4006 671
rect 4166 671 4169 678
rect 4166 668 4206 671
rect 4258 668 4262 671
rect 4338 668 4366 671
rect 4370 668 4414 671
rect 4570 668 4574 671
rect 4914 668 4974 671
rect 5026 668 5054 671
rect 5194 668 5230 671
rect 154 658 198 661
rect 254 661 257 668
rect 1566 662 1569 668
rect 226 658 257 661
rect 282 658 422 661
rect 530 658 590 661
rect 826 658 862 661
rect 890 658 910 661
rect 970 658 990 661
rect 1026 658 1046 661
rect 1118 658 1166 661
rect 1278 658 1390 661
rect 1634 659 1646 661
rect 1630 658 1646 659
rect 2030 661 2033 668
rect 1810 658 2033 661
rect 2042 658 2134 661
rect 2330 658 2350 661
rect 2370 658 2438 661
rect 2442 658 2462 661
rect 2478 661 2481 668
rect 2478 658 2494 661
rect 2506 658 2518 661
rect 2546 658 2654 661
rect 2658 658 2678 661
rect 2714 658 2726 661
rect 2770 658 2790 661
rect 2882 658 2910 661
rect 2978 658 3022 661
rect 3026 658 3094 661
rect 3154 658 3230 661
rect 3322 658 3326 661
rect 3402 658 3489 661
rect 3714 658 3726 661
rect 3786 658 3814 661
rect 3842 658 3934 661
rect 3954 658 3982 661
rect 4034 658 4038 661
rect 4098 658 4102 661
rect 4106 658 4134 661
rect 4202 658 4230 661
rect 4234 658 4246 661
rect 4622 658 4822 661
rect 4826 658 4862 661
rect 4866 658 4886 661
rect 4946 658 4982 661
rect 4986 658 5102 661
rect 5342 661 5346 662
rect 5162 658 5346 661
rect 114 648 222 651
rect 262 651 265 658
rect 1118 652 1121 658
rect 1278 652 1281 658
rect 3486 652 3489 658
rect 4622 652 4625 658
rect 262 648 286 651
rect 290 648 318 651
rect 338 648 342 651
rect 370 648 398 651
rect 430 648 438 651
rect 442 648 518 651
rect 530 648 534 651
rect 550 648 790 651
rect 1154 648 1182 651
rect 1186 648 1222 651
rect 1426 648 2294 651
rect 2298 648 2358 651
rect 2378 648 2390 651
rect 2442 648 2542 651
rect 2578 648 2734 651
rect 2826 648 2830 651
rect 3002 648 3022 651
rect 3706 648 3838 651
rect 3850 648 3886 651
rect 3962 648 3990 651
rect 3994 648 4014 651
rect 4026 648 4062 651
rect 4066 648 4102 651
rect 4106 648 4158 651
rect 4162 648 4166 651
rect 4314 648 4318 651
rect 4322 648 4358 651
rect 4362 648 4390 651
rect 4394 648 4414 651
rect 4878 648 4918 651
rect 4922 648 4966 651
rect 550 642 553 648
rect 274 638 326 641
rect 498 638 518 641
rect 650 638 902 641
rect 982 641 985 648
rect 982 638 1126 641
rect 1138 638 1198 641
rect 1202 638 1230 641
rect 1234 638 1334 641
rect 1338 638 1438 641
rect 1442 638 1614 641
rect 2066 638 2198 641
rect 2310 638 2318 641
rect 2322 638 2374 641
rect 2510 638 2518 641
rect 2522 638 2558 641
rect 2610 638 2686 641
rect 2762 638 2870 641
rect 2942 641 2945 648
rect 2906 638 2945 641
rect 2950 642 2953 648
rect 2970 638 3558 641
rect 3562 638 3574 641
rect 3682 638 3686 641
rect 3894 641 3897 648
rect 4878 642 4881 648
rect 3894 638 3902 641
rect 4006 638 4030 641
rect 4082 638 4110 641
rect 4114 638 4126 641
rect 4290 638 4654 641
rect 4658 638 4694 641
rect 4698 638 4718 641
rect 4722 638 4742 641
rect 2310 632 2313 638
rect 4006 632 4009 638
rect 226 628 326 631
rect 330 628 414 631
rect 442 628 502 631
rect 802 628 846 631
rect 850 628 942 631
rect 954 628 1126 631
rect 1322 628 1478 631
rect 1498 628 1942 631
rect 1954 628 2286 631
rect 2394 628 2566 631
rect 2578 628 2654 631
rect 2666 628 2886 631
rect 2938 628 2982 631
rect 3698 628 3750 631
rect 4058 628 4078 631
rect 4222 631 4225 638
rect 4082 628 4225 631
rect 418 618 470 621
rect 706 618 886 621
rect 906 618 1102 621
rect 1314 618 1838 621
rect 1930 618 2318 621
rect 2322 618 2758 621
rect 2762 618 3118 621
rect 4030 621 4033 628
rect 3826 618 4033 621
rect 5218 618 5270 621
rect 530 608 766 611
rect 770 608 1046 611
rect 1106 608 1238 611
rect 1450 608 1454 611
rect 1602 608 1958 611
rect 2106 608 2126 611
rect 2466 608 2582 611
rect 2586 608 2630 611
rect 2746 608 3038 611
rect 3578 608 4430 611
rect 344 603 346 607
rect 350 603 353 607
rect 358 603 360 607
rect 1368 603 1370 607
rect 1374 603 1377 607
rect 1382 603 1384 607
rect 2006 602 2009 608
rect 2392 603 2394 607
rect 2398 603 2401 607
rect 2406 603 2408 607
rect 3416 603 3418 607
rect 3422 603 3425 607
rect 3430 603 3432 607
rect 4440 603 4442 607
rect 4446 603 4449 607
rect 4454 603 4456 607
rect 890 598 1022 601
rect 1042 598 1086 601
rect 1098 598 1342 601
rect 1450 598 1494 601
rect 1618 598 1726 601
rect 1762 598 1950 601
rect 2114 598 2118 601
rect 2658 598 2766 601
rect 2818 598 2934 601
rect 2946 598 3030 601
rect 3346 598 3350 601
rect 3786 598 3830 601
rect 4074 598 4102 601
rect 4114 598 4334 601
rect 66 588 982 591
rect 994 588 1302 591
rect 1354 588 2310 591
rect 2314 588 2334 591
rect 2338 588 2374 591
rect 2866 588 3046 591
rect 3050 588 3142 591
rect 3370 588 3574 591
rect 3586 588 3846 591
rect 5282 588 5358 591
rect 682 578 1598 581
rect 1946 578 1982 581
rect 2802 578 2998 581
rect 3674 578 3726 581
rect 3854 581 3857 588
rect 3730 578 3857 581
rect 5146 578 5345 581
rect -26 571 -22 572
rect -26 568 62 571
rect 186 568 206 571
rect 490 568 518 571
rect 522 568 550 571
rect 566 571 569 578
rect 566 568 630 571
rect 818 568 862 571
rect 866 568 966 571
rect 974 568 1070 571
rect 1090 568 1254 571
rect 1410 568 1574 571
rect 1802 568 1830 571
rect 1834 568 1886 571
rect 1978 568 2038 571
rect 2098 568 2174 571
rect 2178 568 2198 571
rect 2430 571 2433 578
rect 2430 568 2534 571
rect 2898 568 2993 571
rect 3114 568 3262 571
rect 3314 568 3614 571
rect 3746 568 3766 571
rect 3770 568 3790 571
rect 3882 568 3894 571
rect 3922 568 3934 571
rect 3970 568 4110 571
rect 4178 568 4182 571
rect 4522 568 4542 571
rect 4570 568 4598 571
rect 5078 571 5081 578
rect 5342 572 5345 578
rect 4602 568 5081 571
rect 5342 568 5346 572
rect 162 558 190 561
rect 410 558 462 561
rect 466 558 502 561
rect 742 561 745 568
rect 742 558 838 561
rect 974 561 977 568
rect 2990 562 2993 568
rect 842 558 977 561
rect 1034 558 1158 561
rect 1234 558 1406 561
rect 1554 558 1662 561
rect 1818 558 1862 561
rect 1866 558 1926 561
rect 1962 558 2070 561
rect 2362 558 2518 561
rect 2522 558 2574 561
rect 2578 558 2614 561
rect 2698 558 2846 561
rect 2850 558 2958 561
rect 2962 558 2974 561
rect 3066 558 3182 561
rect 3242 558 3270 561
rect 3274 558 3390 561
rect 3650 558 3734 561
rect 3754 558 3766 561
rect 3922 558 3958 561
rect 3962 558 3982 561
rect 4818 558 4862 561
rect 5174 561 5177 568
rect 4866 558 5177 561
rect 5242 558 5345 561
rect 710 552 713 558
rect 1494 552 1497 558
rect -26 551 -22 552
rect -26 548 318 551
rect 322 548 326 551
rect 498 548 534 551
rect 634 548 638 551
rect 722 548 774 551
rect 834 548 870 551
rect 914 548 985 551
rect 1026 548 1030 551
rect 1034 548 1182 551
rect 1850 548 1854 551
rect 1890 548 1918 551
rect 2086 551 2089 558
rect 2086 548 2102 551
rect 2258 548 2262 551
rect 2298 548 2414 551
rect 2426 548 2454 551
rect 2526 548 2534 551
rect 2538 548 2542 551
rect 2622 551 2625 558
rect 2622 548 2630 551
rect 2730 548 2774 551
rect 2778 548 2878 551
rect 2954 548 2998 551
rect 3106 548 3150 551
rect 3166 548 3174 551
rect 3178 548 3206 551
rect 3490 548 3510 551
rect 3630 551 3633 558
rect 5342 552 5345 558
rect 3630 548 3654 551
rect 3658 548 3686 551
rect 3786 548 3806 551
rect 3834 548 3870 551
rect 3914 548 3934 551
rect 3994 548 4014 551
rect 4042 548 4134 551
rect 4170 548 4190 551
rect 4198 548 4278 551
rect 4282 548 4310 551
rect 4314 548 4350 551
rect 4530 548 4550 551
rect 4594 548 4622 551
rect 4642 548 4678 551
rect 4682 548 4694 551
rect 4850 548 4870 551
rect 4874 548 4886 551
rect 5010 548 5118 551
rect 5122 548 5214 551
rect 5258 548 5278 551
rect 5342 548 5346 552
rect 518 542 521 548
rect 982 542 985 548
rect 202 538 222 541
rect 690 538 710 541
rect 754 538 782 541
rect 786 538 966 541
rect 1018 538 1078 541
rect 1218 538 1265 541
rect 1414 541 1417 548
rect 1306 538 1417 541
rect 1486 541 1489 548
rect 1486 538 1542 541
rect 1634 538 1694 541
rect 1698 538 1710 541
rect 1974 541 1977 548
rect 1714 538 1977 541
rect 2322 538 2350 541
rect 2354 538 2398 541
rect 2450 538 2486 541
rect 2490 538 2526 541
rect 2530 538 2590 541
rect 2730 538 2734 541
rect 2794 538 2950 541
rect 3014 541 3017 548
rect 3014 538 3054 541
rect 3058 538 3094 541
rect 3474 538 3566 541
rect 3570 538 3614 541
rect 3618 538 3670 541
rect 3762 538 3798 541
rect 3950 541 3953 548
rect 3802 538 3953 541
rect 4198 541 4201 548
rect 4194 538 4201 541
rect 4218 538 4262 541
rect 4266 538 4278 541
rect 4842 538 4854 541
rect 4902 541 4905 548
rect 4858 538 4905 541
rect 4962 538 5054 541
rect 5274 538 5278 541
rect 5298 538 5302 541
rect 514 528 558 531
rect 698 528 726 531
rect 730 528 758 531
rect 802 528 806 531
rect 878 528 886 531
rect 906 528 910 531
rect 982 531 985 538
rect 1014 531 1017 538
rect 1262 532 1265 538
rect 3438 532 3441 538
rect 982 528 1017 531
rect 1026 528 1030 531
rect 1410 528 1494 531
rect 1578 528 1622 531
rect 1626 528 1702 531
rect 1930 528 1950 531
rect 1986 528 2022 531
rect 2418 528 2454 531
rect 2834 528 2878 531
rect 2930 528 3022 531
rect 3082 528 3182 531
rect 3186 528 3334 531
rect 3490 528 3582 531
rect 3586 528 3598 531
rect 3682 528 3718 531
rect 3722 528 3830 531
rect 3842 528 3990 531
rect 3994 528 4001 531
rect 4046 531 4049 538
rect 4018 528 4049 531
rect 4146 528 4166 531
rect 4202 528 4270 531
rect 4274 528 4302 531
rect 4606 531 4609 538
rect 4606 528 4646 531
rect 2798 522 2801 528
rect 4054 522 4057 528
rect 938 518 958 521
rect 962 518 1222 521
rect 1290 518 1302 521
rect 1314 518 1366 521
rect 1466 518 1590 521
rect 1946 518 1982 521
rect 2370 518 2510 521
rect 2514 518 2566 521
rect 2570 518 2606 521
rect 2650 518 2670 521
rect 2882 518 3094 521
rect 3202 518 3238 521
rect 3674 518 3822 521
rect 3830 518 4046 521
rect 4330 518 4334 521
rect 118 512 121 518
rect 666 508 686 511
rect 1074 508 1086 511
rect 1090 508 1318 511
rect 1346 508 1774 511
rect 2562 508 2574 511
rect 2578 508 2726 511
rect 3170 508 3190 511
rect 3194 508 3262 511
rect 3266 508 3342 511
rect 3394 508 3702 511
rect 3762 508 3774 511
rect 3830 511 3833 518
rect 3802 508 3833 511
rect 3978 508 4246 511
rect 38 502 41 508
rect 856 503 858 507
rect 862 503 865 507
rect 870 503 872 507
rect 1872 503 1874 507
rect 1878 503 1881 507
rect 1886 503 1888 507
rect 2904 503 2906 507
rect 2910 503 2913 507
rect 2918 503 2920 507
rect 3928 503 3930 507
rect 3934 503 3937 507
rect 3942 503 3944 507
rect 4952 503 4954 507
rect 4958 503 4961 507
rect 4966 503 4968 507
rect 42 498 294 501
rect 298 498 526 501
rect 770 498 790 501
rect 890 498 1110 501
rect 1162 498 1462 501
rect 2002 498 2094 501
rect 2186 498 2190 501
rect 2274 498 2382 501
rect 2626 498 2766 501
rect 2938 498 3454 501
rect 3658 498 3774 501
rect 3994 498 4006 501
rect 4114 498 4142 501
rect 4146 498 4222 501
rect 4226 498 4262 501
rect 4554 498 4862 501
rect 5074 498 5094 501
rect 162 488 198 491
rect 202 488 222 491
rect 234 488 302 491
rect 306 488 390 491
rect 1194 488 1294 491
rect 1298 488 1438 491
rect 1738 488 1878 491
rect 2002 488 2182 491
rect 2226 488 2230 491
rect 2710 488 2718 491
rect 2722 488 2734 491
rect 2754 488 2782 491
rect 2842 488 2870 491
rect 2882 488 3086 491
rect 3562 488 3638 491
rect 3730 488 3814 491
rect 3858 488 4001 491
rect 4050 488 4070 491
rect 4074 488 4102 491
rect 4106 488 4134 491
rect 4506 488 4534 491
rect 4538 488 4614 491
rect 4626 488 4638 491
rect 4642 488 4662 491
rect 4714 488 4849 491
rect 5034 488 5086 491
rect 610 478 670 481
rect 774 478 798 481
rect 822 481 825 488
rect 822 478 838 481
rect 1170 478 1206 481
rect 1530 478 1558 481
rect 1698 478 1838 481
rect 1922 478 1934 481
rect 1938 478 1990 481
rect 2018 478 2022 481
rect 2074 478 2222 481
rect 2770 478 2870 481
rect 2874 478 2910 481
rect 3314 478 3350 481
rect 3470 481 3473 488
rect 3998 482 4001 488
rect 4846 482 4849 488
rect 3418 478 3473 481
rect 3506 478 3574 481
rect 3594 478 3982 481
rect 4442 478 4486 481
rect 4490 478 4518 481
rect 4594 478 4654 481
rect 4658 478 4742 481
rect 4746 478 4822 481
rect 5074 478 5078 481
rect 774 472 777 478
rect 2758 472 2761 478
rect 186 468 310 471
rect 458 468 678 471
rect 738 468 774 471
rect 794 468 862 471
rect 1226 468 1254 471
rect 1346 468 1353 471
rect 398 462 401 468
rect 210 458 262 461
rect 266 458 278 461
rect 554 458 558 461
rect 626 458 646 461
rect 770 458 798 461
rect 914 458 942 461
rect 946 458 950 461
rect 1142 461 1145 468
rect 1082 458 1145 461
rect 1174 461 1177 468
rect 1350 462 1353 468
rect 1546 468 1550 471
rect 1706 468 1726 471
rect 1850 468 1854 471
rect 2206 468 2281 471
rect 2338 468 2350 471
rect 2354 468 2358 471
rect 2418 468 2462 471
rect 2666 468 2694 471
rect 2770 468 2822 471
rect 2962 468 2974 471
rect 3186 468 3214 471
rect 3310 471 3313 478
rect 3238 468 3313 471
rect 3474 468 3665 471
rect 1454 462 1457 468
rect 1174 458 1182 461
rect 1650 458 1702 461
rect 1706 458 1878 461
rect 1974 461 1977 468
rect 2014 462 2017 468
rect 2206 462 2209 468
rect 2278 462 2281 468
rect 1974 458 1998 461
rect 2338 458 2414 461
rect 2418 458 2446 461
rect 2450 458 2526 461
rect 2530 458 2542 461
rect 2682 458 2702 461
rect 2778 458 2798 461
rect 2806 458 2838 461
rect 2878 461 2881 468
rect 3238 462 3241 468
rect 3566 462 3569 468
rect 3662 462 3665 468
rect 3698 468 3726 471
rect 3762 468 3766 471
rect 3898 468 3926 471
rect 4058 468 4094 471
rect 4610 468 4670 471
rect 4674 468 4718 471
rect 4770 468 4790 471
rect 4866 468 4870 471
rect 4954 468 5006 471
rect 5010 468 5030 471
rect 5054 471 5057 478
rect 5034 468 5057 471
rect 5066 468 5126 471
rect 3678 462 3681 468
rect 2858 458 2881 461
rect 2898 458 3006 461
rect 3010 458 3014 461
rect 3250 458 3254 461
rect 3298 458 3449 461
rect 3522 458 3526 461
rect 3530 458 3550 461
rect 3650 458 3654 461
rect 3790 461 3793 468
rect 3790 458 3838 461
rect 3850 458 3902 461
rect 3938 458 4086 461
rect 4134 461 4137 468
rect 4134 458 4158 461
rect 4162 458 4214 461
rect 4386 458 4494 461
rect 4522 458 4558 461
rect 4562 458 4574 461
rect 4642 458 4662 461
rect 4730 458 4806 461
rect 4894 461 4897 468
rect 4894 458 4934 461
rect 4962 458 4982 461
rect 4986 458 5070 461
rect 5074 458 5174 461
rect 378 448 406 451
rect 410 448 446 451
rect 450 448 470 451
rect 474 448 486 451
rect 610 448 686 451
rect 822 451 825 458
rect 822 448 870 451
rect 874 448 958 451
rect 962 448 1014 451
rect 1294 451 1297 458
rect 2806 452 2809 458
rect 3446 452 3449 458
rect 1234 448 1297 451
rect 1410 448 1422 451
rect 1530 448 1534 451
rect 1714 448 1726 451
rect 2002 448 2038 451
rect 2074 448 2558 451
rect 2834 448 2854 451
rect 3474 448 3478 451
rect 3526 448 3550 451
rect 3554 448 3710 451
rect 3930 448 3974 451
rect 4010 448 4065 451
rect 4130 448 4174 451
rect 4306 448 4382 451
rect 4386 448 4446 451
rect 4554 448 4598 451
rect 4682 448 4718 451
rect 4754 448 4798 451
rect 5038 448 5134 451
rect 5138 448 5166 451
rect 5342 451 5346 452
rect 5250 448 5346 451
rect 314 438 710 441
rect 714 438 758 441
rect 762 438 926 441
rect 930 438 990 441
rect 994 438 1006 441
rect 1178 438 1246 441
rect 1250 438 1270 441
rect 1706 438 1742 441
rect 1950 441 1953 448
rect 1950 438 1958 441
rect 2530 438 2718 441
rect 2722 438 2758 441
rect 2762 438 2814 441
rect 2934 441 2937 448
rect 2898 438 2937 441
rect 3510 441 3513 448
rect 3490 438 3513 441
rect 3526 442 3529 448
rect 3578 438 3622 441
rect 3870 441 3873 448
rect 4062 442 4065 448
rect 3626 438 3873 441
rect 3914 438 3966 441
rect 3986 438 4014 441
rect 4174 441 4177 448
rect 4170 438 4177 441
rect 4362 438 4390 441
rect 4394 438 4454 441
rect 4570 438 4614 441
rect 4926 441 4929 448
rect 5038 442 5041 448
rect 4618 438 4761 441
rect 4926 438 4934 441
rect 4938 438 4998 441
rect 5002 438 5014 441
rect 5058 438 5142 441
rect 4758 432 4761 438
rect 722 428 742 431
rect 746 428 950 431
rect 954 428 998 431
rect 1146 428 1374 431
rect 1682 428 1750 431
rect 1922 428 1974 431
rect 2546 428 2678 431
rect 2698 428 2734 431
rect 2802 428 2806 431
rect 3514 428 3630 431
rect 3906 428 3958 431
rect 3962 428 4054 431
rect 4058 428 4150 431
rect 4890 428 4937 431
rect 658 418 830 421
rect 850 418 894 421
rect 898 418 905 421
rect 914 418 966 421
rect 970 418 974 421
rect 978 418 985 421
rect 1074 418 1078 421
rect 1082 418 1582 421
rect 1858 418 1862 421
rect 1866 418 1886 421
rect 1890 418 1958 421
rect 2634 418 2934 421
rect 3442 418 4270 421
rect 4274 418 4318 421
rect 4674 418 4694 421
rect 4870 421 4873 428
rect 4698 418 4873 421
rect 4934 422 4937 428
rect 522 408 526 411
rect 1394 408 1654 411
rect 1658 408 2014 411
rect 2818 408 2838 411
rect 3922 408 4278 411
rect 4282 408 4406 411
rect 4618 408 4686 411
rect 4858 408 5014 411
rect 344 403 346 407
rect 350 403 353 407
rect 358 403 360 407
rect 1368 403 1370 407
rect 1374 403 1377 407
rect 1382 403 1384 407
rect 2392 403 2394 407
rect 2398 403 2401 407
rect 2406 403 2408 407
rect 3416 403 3418 407
rect 3422 403 3425 407
rect 3430 403 3432 407
rect 4440 403 4442 407
rect 4446 403 4449 407
rect 4454 403 4456 407
rect 1698 398 1798 401
rect 1802 398 1814 401
rect 1818 398 1918 401
rect 2418 398 3262 401
rect 3874 398 4022 401
rect 4546 398 4646 401
rect 402 388 1198 391
rect 1794 388 1910 391
rect 1914 388 1926 391
rect 2598 388 2606 391
rect 2610 388 2638 391
rect 2698 388 2974 391
rect 2978 388 2998 391
rect 3370 388 3822 391
rect 3850 388 3910 391
rect 3914 388 4078 391
rect 4082 388 4086 391
rect 4218 388 4742 391
rect 986 378 1390 381
rect 1502 381 1505 388
rect 1502 378 1542 381
rect 1626 378 1678 381
rect 1754 378 1830 381
rect 2098 378 2446 381
rect 2534 378 2630 381
rect 2658 378 2678 381
rect 2754 378 2758 381
rect 2762 378 2798 381
rect 3346 378 4342 381
rect 4346 378 4422 381
rect 4458 378 4502 381
rect 4506 378 4526 381
rect 4530 378 4598 381
rect 4642 378 4646 381
rect 4650 378 4702 381
rect 4914 378 4966 381
rect 4986 378 5142 381
rect 578 368 718 371
rect 722 368 750 371
rect 762 368 926 371
rect 930 368 1150 371
rect 1550 371 1553 378
rect 1362 368 1553 371
rect 1742 371 1745 378
rect 1586 368 1745 371
rect 1846 371 1849 378
rect 1834 368 1849 371
rect 1938 368 1950 371
rect 2086 371 2089 378
rect 2534 372 2537 378
rect 1954 368 2089 371
rect 2106 368 2126 371
rect 2130 368 2174 371
rect 2226 368 2246 371
rect 2258 368 2486 371
rect 2490 368 2534 371
rect 2610 368 2670 371
rect 2726 368 2734 371
rect 2738 368 2782 371
rect 2802 368 2822 371
rect 2858 368 3182 371
rect 3618 368 3718 371
rect 3978 368 4030 371
rect 4386 368 4502 371
rect 4506 368 4686 371
rect 4894 368 4934 371
rect 4938 368 4990 371
rect 4994 368 5038 371
rect 5266 368 5286 371
rect 3334 362 3337 368
rect 4894 362 4897 368
rect 346 358 534 361
rect 570 358 598 361
rect 602 358 622 361
rect 634 358 662 361
rect 786 358 798 361
rect 802 358 830 361
rect 834 358 854 361
rect 858 358 2934 361
rect 3570 358 3638 361
rect 3722 358 3822 361
rect 4006 358 4086 361
rect 4522 358 4566 361
rect 4610 358 4614 361
rect 4690 358 4710 361
rect 4970 358 5006 361
rect -26 351 -22 352
rect -26 348 62 351
rect 66 348 70 351
rect 202 348 238 351
rect 242 348 310 351
rect 362 348 398 351
rect 134 341 137 348
rect 198 341 201 348
rect 498 348 502 351
rect 546 348 582 351
rect 586 348 598 351
rect 666 348 694 351
rect 710 351 713 358
rect 4006 352 4009 358
rect 698 348 713 351
rect 754 348 878 351
rect 1098 348 1102 351
rect 1274 348 1302 351
rect 1378 348 1510 351
rect 1514 348 1518 351
rect 1530 348 1534 351
rect 1546 348 1606 351
rect 1658 348 1686 351
rect 1714 348 1734 351
rect 1742 348 1766 351
rect 1810 348 1854 351
rect 1858 348 1886 351
rect 1890 348 1894 351
rect 2034 348 2038 351
rect 2082 348 2182 351
rect 2218 348 2238 351
rect 2378 348 2398 351
rect 2514 348 2566 351
rect 2634 348 2638 351
rect 2642 348 2670 351
rect 2754 348 2793 351
rect 2850 348 2878 351
rect 3098 348 3102 351
rect 3138 348 3166 351
rect 3334 348 3438 351
rect 3442 348 3454 351
rect 3474 348 3494 351
rect 3546 348 3606 351
rect 3658 348 3662 351
rect 3730 348 3798 351
rect 3802 348 3862 351
rect 3994 348 4006 351
rect 4242 348 4278 351
rect 4506 348 4657 351
rect 4666 348 4697 351
rect 134 338 201 341
rect 218 338 246 341
rect 250 338 358 341
rect 442 338 446 341
rect 538 338 558 341
rect 562 338 574 341
rect 602 338 702 341
rect 706 340 734 341
rect 706 338 737 340
rect 810 338 838 341
rect 850 338 926 341
rect 1050 338 1102 341
rect 1330 338 1334 341
rect 1338 338 1382 341
rect 1426 338 1430 341
rect 1442 338 1566 341
rect 1578 338 1606 341
rect 1610 338 1670 341
rect 1690 338 1702 341
rect 1742 341 1745 348
rect 1730 338 1745 341
rect 1762 338 1822 341
rect 2062 341 2065 348
rect 2790 342 2793 348
rect 2062 338 2142 341
rect 2146 338 2158 341
rect 2194 338 2222 341
rect 2226 338 2254 341
rect 2402 338 2406 341
rect 2426 338 2558 341
rect 2562 338 2606 341
rect 3334 341 3337 348
rect 3298 338 3337 341
rect 38 332 41 338
rect 1142 332 1145 338
rect 3102 332 3105 338
rect 3334 332 3337 338
rect 3390 338 3462 341
rect 3774 338 3822 341
rect 3826 338 3878 341
rect 3978 338 4022 341
rect 4042 338 4062 341
rect 4406 341 4409 348
rect 4406 338 4486 341
rect 4490 338 4542 341
rect 4578 338 4622 341
rect 4654 341 4657 348
rect 4694 342 4697 348
rect 4842 348 4862 351
rect 4902 351 4905 358
rect 4866 348 4905 351
rect 4914 348 4942 351
rect 4970 348 5022 351
rect 5026 348 5046 351
rect 5114 348 5134 351
rect 5270 351 5273 358
rect 5270 348 5286 351
rect 4654 338 4678 341
rect 4726 341 4729 348
rect 4798 341 4801 348
rect 4726 338 4801 341
rect 4810 340 4822 341
rect 4826 340 4854 341
rect 4810 338 4854 340
rect 4858 338 4982 341
rect 5010 338 5078 341
rect 5174 341 5177 348
rect 5082 338 5177 341
rect 5270 338 5278 341
rect 3390 332 3393 338
rect 178 328 214 331
rect 258 328 294 331
rect 298 328 310 331
rect 586 328 606 331
rect 610 328 646 331
rect 666 328 694 331
rect 698 328 726 331
rect 762 328 814 331
rect 818 328 862 331
rect 1266 328 1270 331
rect 1354 328 1486 331
rect 1490 328 1542 331
rect 1546 328 1582 331
rect 1602 328 1606 331
rect 1634 328 1966 331
rect 1970 328 2230 331
rect 2474 328 2478 331
rect 2518 328 2542 331
rect 2546 328 2574 331
rect 2730 328 2958 331
rect 3566 331 3569 338
rect 3774 332 3777 338
rect 4102 332 4105 338
rect 5270 332 5273 338
rect 3538 328 3569 331
rect 3586 328 3614 331
rect 3618 328 3734 331
rect 3834 328 3862 331
rect 3866 328 3998 331
rect 4338 328 4513 331
rect 4538 328 4582 331
rect 4706 328 4782 331
rect 4794 328 4862 331
rect 4930 328 5086 331
rect 5114 328 5142 331
rect 5146 328 5190 331
rect 5294 331 5297 338
rect 5282 328 5297 331
rect 2518 322 2521 328
rect 4510 322 4513 328
rect 26 318 78 321
rect 842 318 1110 321
rect 1178 318 1190 321
rect 1274 318 1334 321
rect 1434 318 1510 321
rect 1522 318 1590 321
rect 1626 318 1638 321
rect 1642 318 1718 321
rect 1746 318 1790 321
rect 1794 318 1838 321
rect 1842 318 1886 321
rect 1890 318 2134 321
rect 2474 318 2478 321
rect 2538 318 2566 321
rect 2578 318 2806 321
rect 2810 318 2830 321
rect 3010 318 3078 321
rect 3154 318 3366 321
rect 3482 318 3542 321
rect 3546 318 3598 321
rect 3610 318 3750 321
rect 3770 318 3782 321
rect 3982 318 3990 321
rect 3994 318 4014 321
rect 4058 318 4078 321
rect 4082 318 4118 321
rect 4122 318 4142 321
rect 4314 318 4350 321
rect 4778 318 4798 321
rect 5298 318 5310 321
rect 234 308 430 311
rect 754 308 766 311
rect 1202 308 1286 311
rect 1322 308 1470 311
rect 1474 308 1494 311
rect 1718 311 1721 318
rect 1718 308 1758 311
rect 2058 308 2086 311
rect 2090 308 2118 311
rect 2314 308 2590 311
rect 2594 308 2758 311
rect 2762 308 2766 311
rect 3210 308 3342 311
rect 3458 308 3518 311
rect 3594 308 3686 311
rect 4146 308 4182 311
rect 856 303 858 307
rect 862 303 865 307
rect 870 303 872 307
rect 1872 303 1874 307
rect 1878 303 1881 307
rect 1886 303 1888 307
rect 2904 303 2906 307
rect 2910 303 2913 307
rect 2918 303 2920 307
rect 3928 303 3930 307
rect 3934 303 3937 307
rect 3942 303 3944 307
rect 4952 303 4954 307
rect 4958 303 4961 307
rect 4966 303 4968 307
rect 82 298 142 301
rect 354 298 438 301
rect 698 298 726 301
rect 730 298 766 301
rect 770 298 838 301
rect 1050 298 1078 301
rect 1242 298 1246 301
rect 1258 298 1302 301
rect 1330 298 1614 301
rect 2018 298 2078 301
rect 2082 298 2110 301
rect 2166 298 2214 301
rect 2738 298 2750 301
rect 3066 298 3086 301
rect 3090 298 3102 301
rect 3106 298 3142 301
rect 3146 298 3270 301
rect 3306 298 3470 301
rect 3482 298 3542 301
rect 3562 298 3582 301
rect 3674 298 3774 301
rect 3778 298 3846 301
rect 4010 298 4022 301
rect 4082 298 4134 301
rect 4714 298 4758 301
rect 4874 298 4905 301
rect 5210 298 5214 301
rect 418 288 886 291
rect 1198 288 1206 291
rect 1210 288 1414 291
rect 1714 288 1774 291
rect 2166 291 2169 298
rect 2034 288 2169 291
rect 2226 288 2350 291
rect 2454 288 2462 291
rect 2466 288 2550 291
rect 2650 288 2678 291
rect 3010 288 3038 291
rect 3250 288 3270 291
rect 3314 288 3326 291
rect 3330 288 3430 291
rect 3434 288 3510 291
rect 3514 288 4214 291
rect 4234 288 4254 291
rect 4338 288 4350 291
rect 4618 288 4678 291
rect 4690 288 4894 291
rect 4902 291 4905 298
rect 4902 288 4993 291
rect 218 278 270 281
rect 286 281 289 288
rect 286 278 326 281
rect 330 278 350 281
rect 482 278 758 281
rect 986 278 1038 281
rect 1138 278 1310 281
rect 1394 278 1422 281
rect 1570 278 1606 281
rect 1610 278 1678 281
rect 1682 278 1750 281
rect 1754 278 1982 281
rect 2142 278 2206 281
rect 2210 278 2222 281
rect 2250 278 2350 281
rect 2354 278 2358 281
rect 2582 281 2585 288
rect 2546 278 2585 281
rect 2706 278 2758 281
rect 2778 278 2790 281
rect 2794 278 2870 281
rect 2914 278 2974 281
rect 2978 278 3014 281
rect 3070 281 3073 288
rect 4990 282 4993 288
rect 5182 288 5206 291
rect 5210 288 5214 291
rect 3018 278 3073 281
rect 3290 278 3294 281
rect 3306 278 3318 281
rect 3402 278 3446 281
rect 3450 278 3494 281
rect 3674 278 3790 281
rect 4006 278 4494 281
rect 4642 278 4734 281
rect 4738 278 4814 281
rect 4866 278 4886 281
rect 5042 278 5062 281
rect 5134 281 5137 288
rect 5182 282 5185 288
rect 5066 278 5137 281
rect 5170 278 5182 281
rect 1086 272 1089 278
rect 50 268 70 271
rect 234 268 262 271
rect 314 268 414 271
rect 530 268 878 271
rect 1210 268 1270 271
rect 1310 271 1313 278
rect 1290 268 1313 271
rect 1330 268 1334 271
rect 1478 268 1526 271
rect 1546 268 1553 271
rect 1594 268 1598 271
rect 1610 268 1614 271
rect 1618 268 1686 271
rect 1706 268 1766 271
rect 1786 268 1830 271
rect 1854 268 1870 271
rect 2142 271 2145 278
rect 1978 268 2145 271
rect 2230 271 2233 278
rect 2186 268 2233 271
rect 2498 268 2518 271
rect 2770 268 2806 271
rect 2906 268 2950 271
rect 2954 268 3094 271
rect 3254 271 3257 278
rect 3254 268 3382 271
rect 3394 268 3438 271
rect 3442 268 3462 271
rect 3494 271 3497 278
rect 4006 272 4009 278
rect 3482 268 3497 271
rect 3586 268 3638 271
rect 3730 268 3750 271
rect 4002 268 4006 271
rect 4122 268 4166 271
rect 4170 268 4177 271
rect 4590 271 4593 278
rect 4242 268 4585 271
rect 4590 268 4662 271
rect 4666 268 4694 271
rect 4750 268 4798 271
rect 4802 268 4902 271
rect 4962 268 4990 271
rect 4994 268 5046 271
rect 5082 268 5110 271
rect 5138 268 5150 271
rect 5154 268 5222 271
rect 5238 268 5246 271
rect 5250 268 5262 271
rect 114 258 134 261
rect 138 258 222 261
rect 250 258 278 261
rect 306 258 334 261
rect 338 258 366 261
rect 682 258 710 261
rect 714 258 750 261
rect 938 258 958 261
rect 1022 261 1025 268
rect 1478 262 1481 268
rect 978 258 1038 261
rect 1250 258 1254 261
rect 1262 258 1398 261
rect 1466 258 1478 261
rect 1558 261 1561 268
rect 1574 261 1577 268
rect 1854 262 1857 268
rect 2150 262 2153 268
rect 2262 262 2265 268
rect 1558 258 1662 261
rect 1666 258 1814 261
rect 1962 258 1990 261
rect 1994 258 2038 261
rect 2266 258 2278 261
rect 2386 258 2430 261
rect 2434 258 2454 261
rect 2514 258 2550 261
rect 2762 258 2798 261
rect 2802 258 2830 261
rect 3010 258 3038 261
rect 3074 258 3078 261
rect 3090 258 3118 261
rect 3234 258 3238 261
rect 3250 258 3342 261
rect 3346 258 3430 261
rect 3434 258 3486 261
rect 3674 258 3726 261
rect 3730 258 3758 261
rect 3762 258 3817 261
rect 3834 258 3870 261
rect 3938 258 4041 261
rect 4114 258 4126 261
rect 4250 258 4318 261
rect 4466 258 4558 261
rect 4582 261 4585 268
rect 4582 258 4614 261
rect 4710 261 4713 268
rect 4726 261 4729 268
rect 4710 258 4729 261
rect 4750 262 4753 268
rect 5246 262 5249 268
rect 4778 258 4822 261
rect 4914 258 4926 261
rect 4930 258 5094 261
rect 5130 258 5158 261
rect 1262 252 1265 258
rect 66 248 86 251
rect 90 248 102 251
rect 106 248 142 251
rect 170 248 318 251
rect 674 248 921 251
rect 38 241 41 248
rect 38 238 190 241
rect 398 241 401 248
rect 798 242 801 248
rect 918 242 921 248
rect 1402 248 1574 251
rect 1658 248 1726 251
rect 1818 248 1846 251
rect 2466 248 2710 251
rect 2714 248 2718 251
rect 2898 248 2942 251
rect 3086 251 3089 258
rect 3814 252 3817 258
rect 4038 252 4041 258
rect 2946 248 3089 251
rect 3250 248 3262 251
rect 3326 248 3366 251
rect 3378 248 3438 251
rect 3474 248 3526 251
rect 3634 248 3646 251
rect 4042 248 4102 251
rect 4106 248 4174 251
rect 4282 248 4294 251
rect 4378 248 4502 251
rect 4650 248 4686 251
rect 4762 248 4774 251
rect 4842 248 4926 251
rect 394 238 401 241
rect 626 238 638 241
rect 690 238 718 241
rect 722 238 750 241
rect 754 238 782 241
rect 946 238 1094 241
rect 1230 241 1233 248
rect 3326 242 3329 248
rect 1230 238 1246 241
rect 1274 238 1342 241
rect 1346 238 1398 241
rect 1450 238 1462 241
rect 1466 238 1526 241
rect 1562 238 1582 241
rect 1586 238 1638 241
rect 1642 238 1926 241
rect 2178 238 2622 241
rect 2834 238 2854 241
rect 2858 238 3158 241
rect 3178 238 3214 241
rect 3362 238 3390 241
rect 3526 241 3529 248
rect 5278 242 5281 248
rect 3526 238 3910 241
rect 3914 238 4310 241
rect 4666 238 4678 241
rect 4730 238 4862 241
rect 4954 238 5006 241
rect 5010 238 5014 241
rect 5086 238 5102 241
rect 5086 232 5089 238
rect 50 228 150 231
rect 1002 228 1030 231
rect 1034 228 1174 231
rect 1178 228 1214 231
rect 1218 228 2414 231
rect 2498 228 3886 231
rect 4898 228 4910 231
rect 4914 228 5017 231
rect 86 218 94 221
rect 98 218 310 221
rect 726 221 729 228
rect 5014 222 5017 228
rect 726 218 958 221
rect 962 218 1022 221
rect 1026 218 1038 221
rect 1290 218 1326 221
rect 1330 218 1358 221
rect 1362 218 1406 221
rect 1410 218 1494 221
rect 1922 218 2014 221
rect 2018 218 2614 221
rect 2626 218 3126 221
rect 3274 218 3718 221
rect 138 208 214 211
rect 218 208 334 211
rect 586 208 726 211
rect 954 208 1078 211
rect 1082 208 1118 211
rect 1194 208 1326 211
rect 1506 208 2086 211
rect 2098 208 2246 211
rect 2882 208 3022 211
rect 3026 208 3062 211
rect 344 203 346 207
rect 350 203 353 207
rect 358 203 360 207
rect 1368 203 1370 207
rect 1374 203 1377 207
rect 1382 203 1384 207
rect 2392 203 2394 207
rect 2398 203 2401 207
rect 2406 203 2408 207
rect 3416 203 3418 207
rect 3422 203 3425 207
rect 3430 203 3432 207
rect 4440 203 4442 207
rect 4446 203 4449 207
rect 4454 203 4456 207
rect 26 198 270 201
rect 274 198 334 201
rect 754 198 806 201
rect 1050 198 1078 201
rect 1082 198 1126 201
rect 1482 198 1518 201
rect 1530 198 1654 201
rect 1666 198 1710 201
rect 2178 198 2270 201
rect 2306 198 2318 201
rect 3002 198 3350 201
rect 3442 198 4094 201
rect 5050 198 5070 201
rect 242 188 1014 191
rect 1018 188 1222 191
rect 1274 188 1390 191
rect 1466 188 1558 191
rect 1562 188 1686 191
rect 1698 188 1782 191
rect 1794 188 1838 191
rect 1850 188 1942 191
rect 1946 188 1982 191
rect 2002 188 2086 191
rect 2114 188 2358 191
rect 2546 188 2630 191
rect 2634 188 2654 191
rect 2658 188 2686 191
rect 2754 188 2870 191
rect 2874 188 2918 191
rect 2954 188 3006 191
rect 3282 188 3622 191
rect 3642 188 3790 191
rect 4106 188 4134 191
rect 4138 188 4158 191
rect 4306 188 4345 191
rect 4342 182 4345 188
rect 5274 188 5286 191
rect 170 178 230 181
rect 322 178 366 181
rect 562 178 574 181
rect 658 178 790 181
rect 818 178 1350 181
rect 1354 178 2430 181
rect 2434 178 3686 181
rect 3694 178 3742 181
rect 3770 178 3942 181
rect 4690 178 4734 181
rect 4878 181 4881 188
rect 4802 178 4881 181
rect 78 171 81 178
rect 78 168 86 171
rect 122 168 390 171
rect 394 168 470 171
rect 546 168 566 171
rect 638 171 641 178
rect 594 168 702 171
rect 794 168 830 171
rect 914 168 1878 171
rect 1882 168 2486 171
rect 2490 168 3102 171
rect 3154 168 3198 171
rect 3226 168 3310 171
rect 3314 168 3326 171
rect 3530 168 3566 171
rect 3694 171 3697 178
rect 3658 168 3697 171
rect 3754 168 3774 171
rect 3802 168 3822 171
rect 3826 168 3854 171
rect 4218 168 4398 171
rect 4682 168 4710 171
rect 4770 168 4846 171
rect 5062 171 5065 178
rect 5062 168 5070 171
rect 5074 168 5102 171
rect 122 158 126 161
rect 162 158 182 161
rect 194 158 374 161
rect 378 158 398 161
rect 402 158 502 161
rect 522 158 574 161
rect 586 158 598 161
rect 634 158 1486 161
rect 1498 158 1622 161
rect 1658 158 1662 161
rect 1690 158 1718 161
rect 1722 158 1758 161
rect 1770 158 2326 161
rect 2330 158 2558 161
rect 2594 158 2678 161
rect 2682 158 2710 161
rect 2738 158 2742 161
rect 2814 158 2822 161
rect 2826 158 2846 161
rect 2866 158 2889 161
rect 2954 158 2958 161
rect 3050 158 3078 161
rect 3142 161 3145 168
rect 3082 158 3145 161
rect 3234 158 3358 161
rect 3410 158 3462 161
rect 3466 158 3574 161
rect 3634 158 3702 161
rect 3710 161 3713 168
rect 3710 158 3742 161
rect 3746 158 3822 161
rect 4426 158 4430 161
rect 4706 158 4718 161
rect 4786 158 4814 161
rect 4882 158 4886 161
rect 4890 158 4926 161
rect 4930 158 4942 161
rect 2886 152 2889 158
rect 4094 152 4097 158
rect 146 148 246 151
rect 338 148 414 151
rect 490 148 494 151
rect 538 148 542 151
rect 562 148 630 151
rect 634 148 646 151
rect 666 148 710 151
rect 714 148 798 151
rect 914 148 918 151
rect 926 148 1033 151
rect 1106 148 1134 151
rect 1138 148 1190 151
rect 254 141 257 148
rect 58 138 257 141
rect 346 138 446 141
rect 498 138 534 141
rect 546 138 598 141
rect 618 138 654 141
rect 782 138 822 141
rect 826 138 838 141
rect 926 141 929 148
rect 1030 142 1033 148
rect 1290 148 1310 151
rect 1338 148 1902 151
rect 1906 148 2206 151
rect 2770 148 2886 151
rect 2906 148 2950 151
rect 2970 148 2998 151
rect 3146 148 3158 151
rect 3242 148 3246 151
rect 3442 148 3638 151
rect 3706 148 3713 151
rect 3794 148 3822 151
rect 4198 151 4201 158
rect 4106 148 4201 151
rect 4342 152 4345 158
rect 4346 148 4358 151
rect 4594 148 4774 151
rect 4794 148 4838 151
rect 5098 148 5126 151
rect 5130 148 5142 151
rect 5210 148 5214 151
rect 5274 148 5302 151
rect 2478 142 2481 148
rect 3710 142 3713 148
rect 898 138 929 141
rect 938 138 958 141
rect 1098 138 1126 141
rect 1130 138 1166 141
rect 1290 138 1294 141
rect 1394 138 1417 141
rect 1450 138 1462 141
rect 1522 138 1534 141
rect 1554 138 1574 141
rect 1578 138 1582 141
rect 1698 138 1726 141
rect 1746 138 1790 141
rect 1802 138 1806 141
rect 1826 138 1878 141
rect 1882 138 1918 141
rect 2042 138 2062 141
rect 2122 138 2145 141
rect 2170 138 2190 141
rect 2386 138 2390 141
rect 2714 138 2734 141
rect 2786 138 2814 141
rect 2818 138 2830 141
rect 2858 138 2862 141
rect 2874 138 2974 141
rect 2994 138 3022 141
rect 3082 138 3102 141
rect 3354 138 3374 141
rect 3378 138 3462 141
rect 3490 138 3518 141
rect 3594 138 3622 141
rect 3626 138 3654 141
rect 3738 138 3782 141
rect 3826 138 3886 141
rect 3918 138 3982 141
rect 4050 138 4054 141
rect 4650 138 4678 141
rect 4746 138 4806 141
rect 4842 138 4862 141
rect 4986 138 4998 141
rect 5002 138 5078 141
rect 5106 138 5142 141
rect 5242 138 5246 141
rect 14 131 17 138
rect 782 132 785 138
rect 14 128 30 131
rect 126 128 177 131
rect 442 128 481 131
rect 562 128 582 131
rect 602 128 670 131
rect 850 128 918 131
rect 946 128 1030 131
rect 1070 131 1073 138
rect 1414 132 1417 138
rect 2142 132 2145 138
rect 2534 132 2537 138
rect 1034 128 1073 131
rect 1194 128 1222 131
rect 1226 128 1230 131
rect 1442 128 1446 131
rect 1514 128 1526 131
rect 1530 128 1558 131
rect 1586 128 1598 131
rect 1706 128 1742 131
rect 1746 128 1854 131
rect 1874 128 2046 131
rect 2130 128 2134 131
rect 2178 128 2182 131
rect 2210 128 2390 131
rect 2394 128 2473 131
rect 2602 128 2758 131
rect 2762 128 2830 131
rect 2838 131 2841 138
rect 2838 128 2894 131
rect 2986 128 3070 131
rect 3090 128 3230 131
rect 3246 128 3350 131
rect 3370 128 3382 131
rect 3402 128 3406 131
rect 3470 128 3486 131
rect 3558 131 3561 138
rect 3918 132 3921 138
rect 3522 128 3561 131
rect 3586 128 3598 131
rect 3602 128 3822 131
rect 4742 131 4745 138
rect 4714 128 4745 131
rect 4770 128 4918 131
rect 5142 131 5145 138
rect 5174 131 5177 138
rect 4938 128 5001 131
rect 5142 128 5177 131
rect 126 122 129 128
rect 174 122 177 128
rect 478 122 481 128
rect 722 118 854 121
rect 1002 118 1166 121
rect 1170 118 1182 121
rect 1242 118 1246 121
rect 1410 118 1454 121
rect 1610 118 1646 121
rect 1650 118 1702 121
rect 1730 118 1830 121
rect 1842 118 1862 121
rect 1866 118 1910 121
rect 1914 118 2462 121
rect 2470 121 2473 128
rect 3246 122 3249 128
rect 3470 122 3473 128
rect 4998 122 5001 128
rect 2470 118 2614 121
rect 2626 118 2702 121
rect 2706 118 2750 121
rect 2794 118 2822 121
rect 2826 118 2846 121
rect 2850 118 2990 121
rect 2994 118 3078 121
rect 3330 118 3454 121
rect 3482 118 3534 121
rect 3538 118 3606 121
rect 3690 118 3774 121
rect 3922 118 4142 121
rect 4170 118 4262 121
rect 4410 118 4622 121
rect 4722 118 4774 121
rect 762 108 838 111
rect 1042 108 1142 111
rect 1154 108 1222 111
rect 1226 108 1502 111
rect 1634 108 1734 111
rect 1778 108 1790 111
rect 1818 108 1846 111
rect 2034 108 2086 111
rect 2098 108 2118 111
rect 2442 108 2502 111
rect 2666 108 2774 111
rect 2930 108 3126 111
rect 3282 108 3502 111
rect 4298 108 4438 111
rect 4490 108 4558 111
rect 846 102 849 108
rect 856 103 858 107
rect 862 103 865 107
rect 870 103 872 107
rect 250 98 262 101
rect 266 98 302 101
rect 746 98 766 101
rect 1490 98 1633 101
rect 1814 101 1817 108
rect 1872 103 1874 107
rect 1878 103 1881 107
rect 1886 103 1888 107
rect 2904 103 2906 107
rect 2910 103 2913 107
rect 2918 103 2920 107
rect 3928 103 3930 107
rect 3934 103 3937 107
rect 3942 103 3944 107
rect 4952 103 4954 107
rect 4958 103 4961 107
rect 4966 103 4968 107
rect 1786 98 1817 101
rect 1898 98 1958 101
rect 1962 98 2366 101
rect 2370 98 2457 101
rect 2522 98 2526 101
rect 2706 98 2726 101
rect 2730 98 2742 101
rect 2746 98 2790 101
rect 2938 98 3150 101
rect 3154 98 3214 101
rect 3258 98 3262 101
rect 3274 98 3382 101
rect 3394 98 3430 101
rect 3722 98 3798 101
rect 3802 98 3910 101
rect 3914 98 3918 101
rect 4338 98 4374 101
rect 4538 98 4606 101
rect 298 88 422 91
rect 474 88 510 91
rect 550 88 566 91
rect 658 88 758 91
rect 834 88 878 91
rect 946 88 990 91
rect 1058 88 1094 91
rect 1342 91 1345 98
rect 1630 92 1633 98
rect 1338 88 1345 91
rect 1362 88 1406 91
rect 1634 88 1678 91
rect 1682 88 1766 91
rect 1786 88 1806 91
rect 1810 88 2446 91
rect 2454 91 2457 98
rect 3982 92 3985 98
rect 4102 92 4105 98
rect 2454 88 3038 91
rect 3066 88 3070 91
rect 3074 88 3174 91
rect 3202 88 3310 91
rect 3314 88 3438 91
rect 3506 88 3606 91
rect 3634 88 3646 91
rect 3650 88 3814 91
rect 3826 88 3846 91
rect 3858 88 3934 91
rect 4258 88 4262 91
rect 4494 91 4497 98
rect 4354 88 4497 91
rect 4554 88 4558 91
rect 4642 88 4918 91
rect 4986 88 4990 91
rect 4994 88 5030 91
rect 5042 88 5086 91
rect 110 78 126 81
rect 262 81 265 88
rect 550 82 553 88
rect 262 78 318 81
rect 370 78 454 81
rect 466 78 494 81
rect 706 78 766 81
rect 770 78 798 81
rect 810 78 830 81
rect 842 78 902 81
rect 946 78 950 81
rect 1018 78 1030 81
rect 1034 78 1070 81
rect 1098 78 1126 81
rect 1130 78 1134 81
rect 1314 78 1478 81
rect 1502 81 1505 88
rect 1482 78 1505 81
rect 1650 78 1670 81
rect 1730 78 1758 81
rect 1770 78 1814 81
rect 2074 78 2102 81
rect 2674 78 2686 81
rect 2698 78 2750 81
rect 2762 78 2782 81
rect 2786 78 2790 81
rect 2806 78 2870 81
rect 2978 78 3094 81
rect 3202 78 3278 81
rect 3290 78 3350 81
rect 3458 78 3526 81
rect 3666 78 3761 81
rect 3826 78 3878 81
rect 4170 78 4270 81
rect 4318 81 4321 88
rect 4306 78 4321 81
rect 5066 78 5094 81
rect 5158 81 5161 88
rect 5098 78 5161 81
rect 5298 78 5302 81
rect 110 72 113 78
rect 510 72 513 78
rect 142 70 161 71
rect 146 68 161 70
rect 242 68 262 71
rect 314 68 414 71
rect 450 68 486 71
rect 534 71 537 78
rect 518 68 537 71
rect 546 68 753 71
rect 786 68 958 71
rect 978 68 1014 71
rect 1082 68 1110 71
rect 1138 68 1214 71
rect 1302 71 1305 78
rect 1290 68 1305 71
rect 1442 68 1478 71
rect 1538 68 1590 71
rect 1594 68 1686 71
rect 1722 68 1750 71
rect 1770 68 1790 71
rect 1914 68 1918 71
rect 1942 71 1945 78
rect 2446 72 2449 78
rect 2494 72 2497 78
rect 2806 72 2809 78
rect 1942 68 2158 71
rect 2234 68 2262 71
rect 2594 68 2678 71
rect 2682 68 2798 71
rect 2818 68 2822 71
rect 2834 68 2846 71
rect 2858 68 2894 71
rect 2898 68 2918 71
rect 2946 68 2990 71
rect 3002 68 3134 71
rect 3138 68 3150 71
rect 3178 68 3190 71
rect 3194 68 3318 71
rect 3346 68 3350 71
rect 3358 68 3361 78
rect 3366 72 3369 78
rect 3574 72 3577 78
rect 3614 72 3617 78
rect 3758 72 3761 78
rect 3418 68 3422 71
rect 3466 68 3550 71
rect 3626 68 3646 71
rect 3714 68 3734 71
rect 3782 70 3889 71
rect 66 58 94 61
rect 158 61 161 68
rect 518 62 521 68
rect 750 62 753 68
rect 98 58 166 61
rect 170 58 174 61
rect 386 58 398 61
rect 426 58 481 61
rect 530 58 566 61
rect 570 58 590 61
rect 594 58 630 61
rect 634 58 654 61
rect 794 58 966 61
rect 970 58 985 61
rect 478 52 481 58
rect 734 52 737 58
rect 982 52 985 58
rect 1042 58 1046 61
rect 1270 58 1278 61
rect 1282 58 1382 61
rect 1442 58 1446 61
rect 1482 58 1486 61
rect 1578 58 1622 61
rect 1626 58 1630 61
rect 1638 58 1678 61
rect 1690 58 1734 61
rect 1738 58 1958 61
rect 2038 62 2041 68
rect 2158 62 2161 68
rect 2018 59 2022 61
rect 2014 58 2022 59
rect 2190 61 2193 68
rect 3786 68 3889 70
rect 4130 68 4214 71
rect 4290 68 4318 71
rect 4322 68 4334 71
rect 4654 71 4657 78
rect 4562 68 4657 71
rect 5006 71 5009 78
rect 5006 68 5206 71
rect 2190 58 2254 61
rect 2322 58 2510 61
rect 2514 59 2534 61
rect 3886 62 3889 68
rect 5294 62 5297 68
rect 2514 58 2537 59
rect 2674 58 2726 61
rect 2730 58 2854 61
rect 2858 58 2974 61
rect 2978 58 3214 61
rect 3218 58 3225 61
rect 3258 58 3598 61
rect 3602 58 3638 61
rect 3658 58 3694 61
rect 3890 58 3918 61
rect 3934 58 4294 61
rect 4418 58 4473 61
rect 4770 58 4798 61
rect 990 52 993 58
rect 266 48 270 51
rect 482 48 686 51
rect 690 48 718 51
rect 1102 51 1105 58
rect 1082 48 1150 51
rect 1210 48 1238 51
rect 1282 48 1310 51
rect 1638 51 1641 58
rect 1618 48 1641 51
rect 1674 48 1782 51
rect 2082 48 2094 51
rect 2098 48 2406 51
rect 2650 48 2758 51
rect 2762 48 3086 51
rect 3122 48 3302 51
rect 3306 48 3350 51
rect 3594 48 3734 51
rect 3762 48 3766 51
rect 3770 48 3814 51
rect 3818 48 3822 51
rect 3858 48 3870 51
rect 3934 51 3937 58
rect 3874 48 3937 51
rect 4358 51 4361 58
rect 4298 48 4361 51
rect 4470 52 4473 58
rect 4906 48 5030 51
rect 5034 48 5038 51
rect 5074 48 5086 51
rect 5118 51 5121 58
rect 5090 48 5121 51
rect 5270 51 5273 58
rect 5266 48 5273 51
rect 278 41 281 48
rect 278 38 702 41
rect 958 41 961 48
rect 958 38 1134 41
rect 1554 38 1582 41
rect 1586 38 1614 41
rect 1654 41 1657 48
rect 1618 38 1657 41
rect 2042 38 2094 41
rect 2706 38 2713 41
rect 2754 38 2982 41
rect 3010 38 3014 41
rect 3018 38 3142 41
rect 3154 38 3494 41
rect 3682 38 3702 41
rect 3722 38 3742 41
rect 3746 38 4390 41
rect 2710 32 2713 38
rect 2050 28 2078 31
rect 2186 28 2214 31
rect 3006 28 3286 31
rect 1230 22 1233 28
rect 3006 22 3009 28
rect 2066 18 2070 21
rect 2250 18 2310 21
rect 526 12 529 18
rect 558 12 561 18
rect 798 12 801 18
rect 1078 12 1081 18
rect 1278 12 1281 18
rect 1390 12 1393 18
rect 2150 12 2153 18
rect 2198 12 2201 18
rect 2558 12 2561 18
rect 2926 12 2929 18
rect 3182 12 3185 18
rect 3558 12 3561 18
rect 3718 12 3721 18
rect 4094 12 4097 18
rect 4486 12 4489 18
rect 490 8 502 11
rect 1106 8 1110 11
rect 1178 8 1182 11
rect 1218 8 1254 11
rect 1298 8 1310 11
rect 1354 8 1358 11
rect 1458 8 1462 11
rect 1482 8 1494 11
rect 1642 8 1646 11
rect 1682 8 1686 11
rect 1738 8 1742 11
rect 1802 8 1806 11
rect 2034 8 2046 11
rect 2106 8 2126 11
rect 2186 8 2190 11
rect 2250 8 2254 11
rect 2274 8 2294 11
rect 2354 8 2358 11
rect 2418 8 2446 11
rect 2978 8 2982 11
rect 3010 8 3014 11
rect 3090 8 3094 11
rect 3338 8 3342 11
rect 3506 8 3510 11
rect 3882 8 3902 11
rect 4050 8 4054 11
rect 4194 8 4198 11
rect 4426 8 4430 11
rect 5242 8 5246 11
rect 344 3 346 7
rect 350 3 353 7
rect 358 3 360 7
rect 1368 3 1370 7
rect 1374 3 1377 7
rect 1382 3 1384 7
rect 2392 3 2394 7
rect 2398 3 2401 7
rect 2406 3 2408 7
rect 3416 3 3418 7
rect 3422 3 3425 7
rect 3430 3 3432 7
rect 4440 3 4442 7
rect 4446 3 4449 7
rect 4454 3 4456 7
<< m4contact >>
rect 858 3703 862 3707
rect 866 3703 869 3707
rect 869 3703 870 3707
rect 1874 3703 1878 3707
rect 1882 3703 1885 3707
rect 1885 3703 1886 3707
rect 2906 3703 2910 3707
rect 2914 3703 2917 3707
rect 2917 3703 2918 3707
rect 3930 3703 3934 3707
rect 3938 3703 3941 3707
rect 3941 3703 3942 3707
rect 4954 3703 4958 3707
rect 4962 3703 4965 3707
rect 4965 3703 4966 3707
rect 2174 3698 2178 3702
rect 2694 3698 2698 3702
rect 3974 3698 3978 3702
rect 3990 3698 3994 3702
rect 4070 3698 4074 3702
rect 4206 3698 4210 3702
rect 4366 3698 4370 3702
rect 5246 3698 5250 3702
rect 1734 3688 1738 3692
rect 2270 3688 2274 3692
rect 2710 3688 2714 3692
rect 3286 3688 3290 3692
rect 4238 3688 4242 3692
rect 4294 3688 4298 3692
rect 942 3678 946 3682
rect 1742 3678 1746 3682
rect 1982 3678 1986 3682
rect 974 3668 978 3672
rect 1366 3668 1370 3672
rect 1790 3668 1794 3672
rect 2358 3668 2362 3672
rect 1206 3658 1210 3662
rect 1422 3658 1426 3662
rect 1734 3658 1738 3662
rect 2462 3658 2466 3662
rect 2518 3658 2522 3662
rect 3366 3658 3370 3662
rect 5174 3658 5178 3662
rect 1142 3648 1146 3652
rect 1502 3648 1506 3652
rect 1614 3648 1618 3652
rect 1630 3648 1634 3652
rect 4086 3648 4090 3652
rect 5238 3648 5242 3652
rect 5310 3648 5314 3652
rect 1742 3638 1746 3642
rect 1846 3638 1850 3642
rect 2302 3638 2306 3642
rect 4078 3618 4082 3622
rect 5262 3618 5266 3622
rect 1334 3608 1338 3612
rect 2670 3608 2674 3612
rect 346 3603 350 3607
rect 354 3603 357 3607
rect 357 3603 358 3607
rect 1370 3603 1374 3607
rect 1378 3603 1381 3607
rect 1381 3603 1382 3607
rect 2394 3603 2398 3607
rect 2402 3603 2405 3607
rect 2405 3603 2406 3607
rect 3418 3603 3422 3607
rect 3426 3603 3429 3607
rect 3429 3603 3430 3607
rect 4442 3603 4446 3607
rect 4450 3603 4453 3607
rect 4453 3603 4454 3607
rect 1358 3598 1362 3602
rect 3126 3578 3130 3582
rect 5358 3568 5362 3572
rect 446 3558 450 3562
rect 742 3558 746 3562
rect 1150 3558 1154 3562
rect 2670 3558 2674 3562
rect 5310 3558 5314 3562
rect 438 3548 442 3552
rect 1358 3548 1362 3552
rect 1478 3548 1482 3552
rect 1862 3548 1866 3552
rect 3630 3548 3634 3552
rect 4110 3548 4114 3552
rect 4238 3548 4242 3552
rect 4494 3548 4498 3552
rect 5190 3548 5194 3552
rect 5286 3548 5290 3552
rect 1094 3538 1098 3542
rect 1190 3538 1194 3542
rect 166 3528 170 3532
rect 438 3528 442 3532
rect 4302 3538 4306 3542
rect 1862 3528 1866 3532
rect 2302 3528 2306 3532
rect 2342 3528 2346 3532
rect 4886 3528 4890 3532
rect 5206 3528 5210 3532
rect 3094 3518 3098 3522
rect 4742 3518 4746 3522
rect 2414 3508 2418 3512
rect 2894 3508 2898 3512
rect 858 3503 862 3507
rect 866 3503 869 3507
rect 869 3503 870 3507
rect 1874 3503 1878 3507
rect 1882 3503 1885 3507
rect 1885 3503 1886 3507
rect 2906 3503 2910 3507
rect 2914 3503 2917 3507
rect 2917 3503 2918 3507
rect 3930 3503 3934 3507
rect 3938 3503 3941 3507
rect 3941 3503 3942 3507
rect 4954 3503 4958 3507
rect 4962 3503 4965 3507
rect 4965 3503 4966 3507
rect 422 3498 426 3502
rect 2046 3498 2050 3502
rect 2350 3498 2354 3502
rect 1838 3488 1842 3492
rect 2990 3488 2994 3492
rect 750 3468 754 3472
rect 1198 3468 1202 3472
rect 1670 3478 1674 3482
rect 1846 3478 1850 3482
rect 4086 3478 4090 3482
rect 4478 3478 4482 3482
rect 4574 3478 4578 3482
rect 5014 3478 5018 3482
rect 1966 3468 1970 3472
rect 2190 3468 2194 3472
rect 2222 3468 2226 3472
rect 2310 3468 2314 3472
rect 2326 3468 2330 3472
rect 2982 3468 2986 3472
rect 4614 3468 4618 3472
rect 5294 3468 5298 3472
rect 254 3458 258 3462
rect 446 3458 450 3462
rect 1174 3458 1178 3462
rect 2990 3458 2994 3462
rect 4366 3458 4370 3462
rect 4390 3458 4394 3462
rect 4494 3458 4498 3462
rect 4670 3458 4674 3462
rect 4886 3458 4890 3462
rect 1678 3448 1682 3452
rect 2222 3448 2226 3452
rect 2894 3448 2898 3452
rect 5270 3458 5274 3462
rect 3710 3448 3714 3452
rect 4334 3448 4338 3452
rect 1534 3438 1538 3442
rect 1702 3438 1706 3442
rect 1710 3438 1714 3442
rect 3782 3438 3786 3442
rect 4726 3438 4730 3442
rect 5270 3438 5274 3442
rect 5278 3438 5282 3442
rect 646 3428 650 3432
rect 2718 3428 2722 3432
rect 974 3418 978 3422
rect 2486 3418 2490 3422
rect 2726 3408 2730 3412
rect 3534 3408 3538 3412
rect 346 3403 350 3407
rect 354 3403 357 3407
rect 357 3403 358 3407
rect 1370 3403 1374 3407
rect 1378 3403 1381 3407
rect 1381 3403 1382 3407
rect 2394 3403 2398 3407
rect 2402 3403 2405 3407
rect 2405 3403 2406 3407
rect 3418 3403 3422 3407
rect 3426 3403 3429 3407
rect 3429 3403 3430 3407
rect 4442 3403 4446 3407
rect 4450 3403 4453 3407
rect 4453 3403 4454 3407
rect 686 3398 690 3402
rect 1142 3398 1146 3402
rect 2014 3398 2018 3402
rect 3950 3398 3954 3402
rect 4646 3398 4650 3402
rect 62 3388 66 3392
rect 118 3388 122 3392
rect 2094 3388 2098 3392
rect 2982 3388 2986 3392
rect 5014 3388 5018 3392
rect 494 3378 498 3382
rect 2598 3378 2602 3382
rect 2654 3378 2658 3382
rect 462 3368 466 3372
rect 534 3368 538 3372
rect 590 3368 594 3372
rect 702 3368 706 3372
rect 1182 3368 1186 3372
rect 1718 3368 1722 3372
rect 2070 3368 2074 3372
rect 5254 3368 5258 3372
rect 846 3358 850 3362
rect 1022 3358 1026 3362
rect 1070 3358 1074 3362
rect 2358 3358 2362 3362
rect 2606 3358 2610 3362
rect 3846 3358 3850 3362
rect 4102 3358 4106 3362
rect 4686 3358 4690 3362
rect 4998 3358 5002 3362
rect 5302 3358 5306 3362
rect 630 3348 634 3352
rect 1198 3348 1202 3352
rect 1254 3348 1258 3352
rect 1278 3348 1282 3352
rect 1462 3348 1466 3352
rect 1710 3348 1714 3352
rect 2062 3348 2066 3352
rect 2838 3348 2842 3352
rect 3182 3348 3186 3352
rect 3766 3348 3770 3352
rect 4278 3348 4282 3352
rect 4734 3348 4738 3352
rect 5014 3348 5018 3352
rect 5022 3348 5026 3352
rect 5182 3348 5186 3352
rect 230 3338 234 3342
rect 406 3338 410 3342
rect 606 3338 610 3342
rect 686 3338 690 3342
rect 782 3338 786 3342
rect 966 3338 970 3342
rect 1350 3338 1354 3342
rect 1374 3338 1378 3342
rect 1702 3338 1706 3342
rect 1766 3338 1770 3342
rect 1814 3338 1818 3342
rect 2886 3338 2890 3342
rect 4886 3338 4890 3342
rect 4910 3338 4914 3342
rect 5006 3338 5010 3342
rect 5214 3338 5218 3342
rect 486 3328 490 3332
rect 646 3328 650 3332
rect 1454 3328 1458 3332
rect 1518 3328 1522 3332
rect 1670 3328 1674 3332
rect 2094 3328 2098 3332
rect 2478 3328 2482 3332
rect 3062 3328 3066 3332
rect 462 3318 466 3322
rect 1070 3318 1074 3322
rect 1182 3318 1186 3322
rect 1406 3318 1410 3322
rect 1422 3318 1426 3322
rect 4550 3318 4554 3322
rect 622 3308 626 3312
rect 942 3308 946 3312
rect 950 3308 954 3312
rect 958 3308 962 3312
rect 3366 3308 3370 3312
rect 858 3303 862 3307
rect 866 3303 869 3307
rect 869 3303 870 3307
rect 486 3298 490 3302
rect 910 3298 914 3302
rect 1874 3303 1878 3307
rect 1882 3303 1885 3307
rect 1885 3303 1886 3307
rect 2906 3303 2910 3307
rect 2914 3303 2917 3307
rect 2917 3303 2918 3307
rect 3930 3303 3934 3307
rect 3938 3303 3941 3307
rect 3941 3303 3942 3307
rect 4954 3303 4958 3307
rect 4962 3303 4965 3307
rect 4965 3303 4966 3307
rect 990 3298 994 3302
rect 1190 3298 1194 3302
rect 1710 3298 1714 3302
rect 2038 3298 2042 3302
rect 3086 3298 3090 3302
rect 3350 3298 3354 3302
rect 3542 3298 3546 3302
rect 710 3288 714 3292
rect 806 3288 810 3292
rect 1062 3288 1066 3292
rect 1262 3288 1266 3292
rect 2182 3288 2186 3292
rect 3038 3288 3042 3292
rect 3070 3288 3074 3292
rect 3846 3288 3850 3292
rect 4670 3288 4674 3292
rect 4870 3288 4874 3292
rect 4950 3288 4954 3292
rect 5246 3288 5250 3292
rect 1686 3278 1690 3282
rect 1742 3278 1746 3282
rect 2726 3278 2730 3282
rect 4886 3278 4890 3282
rect 4942 3278 4946 3282
rect 4958 3278 4962 3282
rect 126 3268 130 3272
rect 782 3268 786 3272
rect 1678 3268 1682 3272
rect 3070 3268 3074 3272
rect 4718 3268 4722 3272
rect 4918 3268 4922 3272
rect 14 3258 18 3262
rect 422 3258 426 3262
rect 790 3258 794 3262
rect 1038 3258 1042 3262
rect 1798 3258 1802 3262
rect 2054 3258 2058 3262
rect 2518 3258 2522 3262
rect 3398 3258 3402 3262
rect 4110 3258 4114 3262
rect 902 3248 906 3252
rect 1966 3248 1970 3252
rect 2038 3248 2042 3252
rect 2142 3248 2146 3252
rect 2182 3248 2186 3252
rect 2286 3248 2290 3252
rect 3190 3248 3194 3252
rect 4270 3258 4274 3262
rect 4742 3258 4746 3262
rect 5286 3258 5290 3262
rect 174 3238 178 3242
rect 478 3238 482 3242
rect 502 3238 506 3242
rect 1526 3238 1530 3242
rect 2838 3238 2842 3242
rect 3086 3238 3090 3242
rect 4734 3238 4738 3242
rect 1566 3228 1570 3232
rect 2342 3228 2346 3232
rect 4558 3228 4562 3232
rect 5278 3228 5282 3232
rect 438 3218 442 3222
rect 5182 3218 5186 3222
rect 2718 3208 2722 3212
rect 346 3203 350 3207
rect 354 3203 357 3207
rect 357 3203 358 3207
rect 1370 3203 1374 3207
rect 1378 3203 1381 3207
rect 1381 3203 1382 3207
rect 2394 3203 2398 3207
rect 2402 3203 2405 3207
rect 2405 3203 2406 3207
rect 3418 3203 3422 3207
rect 3426 3203 3429 3207
rect 3429 3203 3430 3207
rect 4442 3203 4446 3207
rect 4450 3203 4453 3207
rect 4453 3203 4454 3207
rect 918 3198 922 3202
rect 2702 3198 2706 3202
rect 2822 3198 2826 3202
rect 2550 3188 2554 3192
rect 3950 3188 3954 3192
rect 4910 3188 4914 3192
rect 5294 3188 5298 3192
rect 1790 3178 1794 3182
rect 3342 3178 3346 3182
rect 4870 3178 4874 3182
rect 5294 3178 5298 3182
rect 438 3168 442 3172
rect 3198 3168 3202 3172
rect 4302 3168 4306 3172
rect 486 3158 490 3162
rect 966 3158 970 3162
rect 4878 3158 4882 3162
rect 5254 3158 5258 3162
rect 1510 3148 1514 3152
rect 2014 3148 2018 3152
rect 2190 3148 2194 3152
rect 3014 3148 3018 3152
rect 3086 3148 3090 3152
rect 3406 3148 3410 3152
rect 3870 3148 3874 3152
rect 422 3138 426 3142
rect 558 3138 562 3142
rect 574 3138 578 3142
rect 630 3138 634 3142
rect 638 3138 642 3142
rect 686 3138 690 3142
rect 750 3138 754 3142
rect 2822 3138 2826 3142
rect 3054 3138 3058 3142
rect 3366 3138 3370 3142
rect 3726 3138 3730 3142
rect 1510 3128 1514 3132
rect 1526 3128 1530 3132
rect 2070 3128 2074 3132
rect 2558 3128 2562 3132
rect 3774 3128 3778 3132
rect 4270 3128 4274 3132
rect 182 3118 186 3122
rect 422 3118 426 3122
rect 646 3118 650 3122
rect 670 3118 674 3122
rect 982 3118 986 3122
rect 2718 3118 2722 3122
rect 454 3108 458 3112
rect 606 3108 610 3112
rect 614 3108 618 3112
rect 1750 3108 1754 3112
rect 2238 3108 2242 3112
rect 2310 3108 2314 3112
rect 2550 3108 2554 3112
rect 2702 3108 2706 3112
rect 2926 3108 2930 3112
rect 3390 3108 3394 3112
rect 858 3103 862 3107
rect 866 3103 869 3107
rect 869 3103 870 3107
rect 1874 3103 1878 3107
rect 1882 3103 1885 3107
rect 1885 3103 1886 3107
rect 2906 3103 2910 3107
rect 2914 3103 2917 3107
rect 2917 3103 2918 3107
rect 3930 3103 3934 3107
rect 3938 3103 3941 3107
rect 3941 3103 3942 3107
rect 4954 3103 4958 3107
rect 4962 3103 4965 3107
rect 4965 3103 4966 3107
rect 406 3098 410 3102
rect 838 3098 842 3102
rect 1406 3098 1410 3102
rect 1606 3098 1610 3102
rect 3358 3098 3362 3102
rect 3910 3098 3914 3102
rect 1614 3088 1618 3092
rect 1718 3088 1722 3092
rect 1982 3088 1986 3092
rect 3246 3088 3250 3092
rect 4654 3088 4658 3092
rect 4942 3088 4946 3092
rect 454 3078 458 3082
rect 1950 3078 1954 3082
rect 2414 3078 2418 3082
rect 2982 3078 2986 3082
rect 3118 3078 3122 3082
rect 670 3068 674 3072
rect 918 3068 922 3072
rect 1214 3068 1218 3072
rect 2662 3068 2666 3072
rect 3030 3068 3034 3072
rect 3446 3068 3450 3072
rect 3846 3068 3850 3072
rect 3910 3068 3914 3072
rect 574 3058 578 3062
rect 1230 3058 1234 3062
rect 1718 3058 1722 3062
rect 1854 3058 1858 3062
rect 2366 3058 2370 3062
rect 3214 3058 3218 3062
rect 3870 3058 3874 3062
rect 5302 3058 5306 3062
rect 1214 3048 1218 3052
rect 1326 3048 1330 3052
rect 1982 3048 1986 3052
rect 3982 3048 3986 3052
rect 4278 3048 4282 3052
rect 5230 3048 5234 3052
rect 1830 3038 1834 3042
rect 3198 3038 3202 3042
rect 2374 3028 2378 3032
rect 3614 3028 3618 3032
rect 4110 3028 4114 3032
rect 5054 3028 5058 3032
rect 230 3018 234 3022
rect 974 3018 978 3022
rect 2046 3018 2050 3022
rect 2606 3018 2610 3022
rect 3382 3018 3386 3022
rect 3046 3008 3050 3012
rect 3398 3008 3402 3012
rect 346 3003 350 3007
rect 354 3003 357 3007
rect 357 3003 358 3007
rect 1370 3003 1374 3007
rect 1378 3003 1381 3007
rect 1381 3003 1382 3007
rect 2394 3003 2398 3007
rect 2402 3003 2405 3007
rect 2405 3003 2406 3007
rect 3418 3003 3422 3007
rect 3426 3003 3429 3007
rect 3429 3003 3430 3007
rect 4442 3003 4446 3007
rect 4450 3003 4453 3007
rect 4453 3003 4454 3007
rect 1478 2998 1482 3002
rect 3030 2998 3034 3002
rect 3406 2998 3410 3002
rect 478 2988 482 2992
rect 846 2988 850 2992
rect 1518 2988 1522 2992
rect 3366 2988 3370 2992
rect 3486 2988 3490 2992
rect 878 2958 882 2962
rect 3126 2958 3130 2962
rect 3222 2958 3226 2962
rect 3406 2958 3410 2962
rect 3582 2958 3586 2962
rect 3622 2958 3626 2962
rect 366 2948 370 2952
rect 662 2948 666 2952
rect 862 2948 866 2952
rect 1006 2948 1010 2952
rect 1078 2948 1082 2952
rect 1294 2948 1298 2952
rect 782 2938 786 2942
rect 1654 2948 1658 2952
rect 1710 2948 1714 2952
rect 2038 2948 2042 2952
rect 3430 2948 3434 2952
rect 3438 2948 3442 2952
rect 3718 2948 3722 2952
rect 5238 2948 5242 2952
rect 1198 2938 1202 2942
rect 2582 2938 2586 2942
rect 3198 2938 3202 2942
rect 3470 2938 3474 2942
rect 3718 2938 3722 2942
rect 3734 2938 3738 2942
rect 5270 2938 5274 2942
rect 550 2928 554 2932
rect 1006 2928 1010 2932
rect 3238 2928 3242 2932
rect 3438 2928 3442 2932
rect 5222 2928 5226 2932
rect 54 2918 58 2922
rect 366 2918 370 2922
rect 3382 2918 3386 2922
rect 3462 2918 3466 2922
rect 4214 2918 4218 2922
rect 14 2908 18 2912
rect 502 2908 506 2912
rect 2350 2908 2354 2912
rect 858 2903 862 2907
rect 866 2903 869 2907
rect 869 2903 870 2907
rect 1874 2903 1878 2907
rect 1882 2903 1885 2907
rect 1885 2903 1886 2907
rect 2906 2903 2910 2907
rect 2914 2903 2917 2907
rect 2917 2903 2918 2907
rect 3930 2903 3934 2907
rect 3938 2903 3941 2907
rect 3941 2903 3942 2907
rect 4954 2903 4958 2907
rect 4962 2903 4965 2907
rect 4965 2903 4966 2907
rect 254 2898 258 2902
rect 742 2898 746 2902
rect 2638 2898 2642 2902
rect 3734 2898 3738 2902
rect 1238 2888 1242 2892
rect 1406 2888 1410 2892
rect 1582 2888 1586 2892
rect 2558 2888 2562 2892
rect 3582 2878 3586 2882
rect 2246 2868 2250 2872
rect 2566 2868 2570 2872
rect 2678 2868 2682 2872
rect 398 2858 402 2862
rect 430 2858 434 2862
rect 902 2858 906 2862
rect 1006 2858 1010 2862
rect 1606 2858 1610 2862
rect 1766 2858 1770 2862
rect 1966 2858 1970 2862
rect 2022 2858 2026 2862
rect 2582 2858 2586 2862
rect 3134 2858 3138 2862
rect 3262 2858 3266 2862
rect 4374 2858 4378 2862
rect 1390 2848 1394 2852
rect 2670 2848 2674 2852
rect 3022 2848 3026 2852
rect 3198 2848 3202 2852
rect 3382 2848 3386 2852
rect 686 2838 690 2842
rect 2038 2838 2042 2842
rect 2822 2838 2826 2842
rect 414 2828 418 2832
rect 670 2828 674 2832
rect 1294 2828 1298 2832
rect 4070 2828 4074 2832
rect 4886 2828 4890 2832
rect 3614 2818 3618 2822
rect 2510 2808 2514 2812
rect 3022 2808 3026 2812
rect 346 2803 350 2807
rect 354 2803 357 2807
rect 357 2803 358 2807
rect 1370 2803 1374 2807
rect 1378 2803 1381 2807
rect 1381 2803 1382 2807
rect 2394 2803 2398 2807
rect 2402 2803 2405 2807
rect 2405 2803 2406 2807
rect 3418 2803 3422 2807
rect 3426 2803 3429 2807
rect 3429 2803 3430 2807
rect 4442 2803 4446 2807
rect 4450 2803 4453 2807
rect 4453 2803 4454 2807
rect 910 2798 914 2802
rect 2598 2798 2602 2802
rect 2926 2798 2930 2802
rect 3750 2798 3754 2802
rect 166 2788 170 2792
rect 1334 2788 1338 2792
rect 1766 2788 1770 2792
rect 2054 2788 2058 2792
rect 1646 2778 1650 2782
rect 2470 2778 2474 2782
rect 3214 2778 3218 2782
rect 1134 2768 1138 2772
rect 3126 2768 3130 2772
rect 5134 2768 5138 2772
rect 2470 2758 2474 2762
rect 3406 2758 3410 2762
rect 3598 2758 3602 2762
rect 710 2748 714 2752
rect 782 2748 786 2752
rect 974 2748 978 2752
rect 1518 2748 1522 2752
rect 2182 2748 2186 2752
rect 886 2738 890 2742
rect 1118 2738 1122 2742
rect 2126 2738 2130 2742
rect 3390 2748 3394 2752
rect 3622 2748 3626 2752
rect 3750 2748 3754 2752
rect 3870 2748 3874 2752
rect 3966 2748 3970 2752
rect 4294 2748 4298 2752
rect 2638 2738 2642 2742
rect 2718 2738 2722 2742
rect 3342 2738 3346 2742
rect 3486 2738 3490 2742
rect 3558 2738 3562 2742
rect 3894 2738 3898 2742
rect 4502 2748 4506 2752
rect 5102 2748 5106 2752
rect 4550 2738 4554 2742
rect 4902 2738 4906 2742
rect 718 2728 722 2732
rect 1446 2728 1450 2732
rect 1798 2728 1802 2732
rect 1934 2728 1938 2732
rect 2062 2728 2066 2732
rect 2134 2728 2138 2732
rect 2678 2728 2682 2732
rect 3030 2728 3034 2732
rect 3598 2728 3602 2732
rect 5022 2728 5026 2732
rect 1830 2718 1834 2722
rect 2654 2718 2658 2722
rect 3558 2718 3562 2722
rect 3726 2718 3730 2722
rect 398 2708 402 2712
rect 886 2708 890 2712
rect 974 2708 978 2712
rect 1718 2708 1722 2712
rect 4710 2708 4714 2712
rect 858 2703 862 2707
rect 866 2703 869 2707
rect 869 2703 870 2707
rect 1874 2703 1878 2707
rect 1882 2703 1885 2707
rect 1885 2703 1886 2707
rect 2906 2703 2910 2707
rect 2914 2703 2917 2707
rect 2917 2703 2918 2707
rect 3930 2703 3934 2707
rect 3938 2703 3941 2707
rect 3941 2703 3942 2707
rect 4954 2703 4958 2707
rect 4962 2703 4965 2707
rect 4965 2703 4966 2707
rect 1174 2698 1178 2702
rect 1814 2698 1818 2702
rect 1902 2698 1906 2702
rect 150 2688 154 2692
rect 1126 2688 1130 2692
rect 1734 2688 1738 2692
rect 2302 2688 2306 2692
rect 3222 2698 3226 2702
rect 4678 2698 4682 2702
rect 4734 2698 4738 2702
rect 5270 2698 5274 2702
rect 3054 2688 3058 2692
rect 3446 2688 3450 2692
rect 3470 2688 3474 2692
rect 3590 2688 3594 2692
rect 5302 2688 5306 2692
rect 678 2678 682 2682
rect 982 2678 986 2682
rect 998 2678 1002 2682
rect 1062 2678 1066 2682
rect 2262 2678 2266 2682
rect 2590 2678 2594 2682
rect 2654 2678 2658 2682
rect 3382 2678 3386 2682
rect 5302 2678 5306 2682
rect 166 2668 170 2672
rect 1094 2668 1098 2672
rect 2070 2668 2074 2672
rect 2382 2668 2386 2672
rect 3614 2668 3618 2672
rect 4878 2668 4882 2672
rect 5294 2668 5298 2672
rect 806 2658 810 2662
rect 1126 2658 1130 2662
rect 1982 2658 1986 2662
rect 2366 2658 2370 2662
rect 2702 2658 2706 2662
rect 2974 2658 2978 2662
rect 3526 2658 3530 2662
rect 3694 2658 3698 2662
rect 5150 2658 5154 2662
rect 5294 2658 5298 2662
rect 2446 2648 2450 2652
rect 166 2638 170 2642
rect 4742 2638 4746 2642
rect 5270 2648 5274 2652
rect 5102 2638 5106 2642
rect 526 2628 530 2632
rect 542 2628 546 2632
rect 1990 2628 1994 2632
rect 2582 2628 2586 2632
rect 3326 2628 3330 2632
rect 3998 2628 4002 2632
rect 5142 2628 5146 2632
rect 5294 2628 5298 2632
rect 2406 2618 2410 2622
rect 14 2608 18 2612
rect 1126 2608 1130 2612
rect 1390 2608 1394 2612
rect 346 2603 350 2607
rect 354 2603 357 2607
rect 357 2603 358 2607
rect 1370 2603 1374 2607
rect 1378 2603 1381 2607
rect 1381 2603 1382 2607
rect 2394 2603 2398 2607
rect 2402 2603 2405 2607
rect 2405 2603 2406 2607
rect 3418 2603 3422 2607
rect 3426 2603 3429 2607
rect 3429 2603 3430 2607
rect 4442 2603 4446 2607
rect 4450 2603 4453 2607
rect 4453 2603 4454 2607
rect 3014 2598 3018 2602
rect 366 2588 370 2592
rect 998 2588 1002 2592
rect 1606 2588 1610 2592
rect 1750 2588 1754 2592
rect 1950 2588 1954 2592
rect 2142 2588 2146 2592
rect 2462 2588 2466 2592
rect 2662 2588 2666 2592
rect 3590 2588 3594 2592
rect 3702 2588 3706 2592
rect 1118 2578 1122 2582
rect 1654 2578 1658 2582
rect 1958 2578 1962 2582
rect 2262 2578 2266 2582
rect 4678 2578 4682 2582
rect 902 2568 906 2572
rect 630 2558 634 2562
rect 862 2558 866 2562
rect 3678 2558 3682 2562
rect 4030 2558 4034 2562
rect 4718 2558 4722 2562
rect 5294 2558 5298 2562
rect 14 2548 18 2552
rect 414 2548 418 2552
rect 662 2548 666 2552
rect 1070 2548 1074 2552
rect 1822 2548 1826 2552
rect 134 2538 138 2542
rect 206 2538 210 2542
rect 510 2538 514 2542
rect 2022 2548 2026 2552
rect 2294 2548 2298 2552
rect 2302 2548 2306 2552
rect 2870 2548 2874 2552
rect 3198 2548 3202 2552
rect 3542 2548 3546 2552
rect 3638 2548 3642 2552
rect 4126 2548 4130 2552
rect 4526 2548 4530 2552
rect 4838 2548 4842 2552
rect 5094 2548 5098 2552
rect 1646 2538 1650 2542
rect 1678 2538 1682 2542
rect 2158 2538 2162 2542
rect 2254 2538 2258 2542
rect 2478 2538 2482 2542
rect 2494 2538 2498 2542
rect 2774 2538 2778 2542
rect 2814 2538 2818 2542
rect 4246 2538 4250 2542
rect 5166 2538 5170 2542
rect 5302 2538 5306 2542
rect 150 2528 154 2532
rect 494 2528 498 2532
rect 1310 2528 1314 2532
rect 1334 2528 1338 2532
rect 1702 2528 1706 2532
rect 2150 2528 2154 2532
rect 2790 2528 2794 2532
rect 3702 2528 3706 2532
rect 3950 2528 3954 2532
rect 4734 2528 4738 2532
rect 5014 2528 5018 2532
rect 5302 2528 5306 2532
rect 118 2518 122 2522
rect 678 2518 682 2522
rect 1318 2518 1322 2522
rect 2638 2518 2642 2522
rect 3750 2518 3754 2522
rect 430 2508 434 2512
rect 1334 2508 1338 2512
rect 1526 2508 1530 2512
rect 1670 2508 1674 2512
rect 1894 2508 1898 2512
rect 3246 2508 3250 2512
rect 3342 2508 3346 2512
rect 3950 2508 3954 2512
rect 4614 2508 4618 2512
rect 4982 2508 4986 2512
rect 5278 2508 5282 2512
rect 5294 2508 5298 2512
rect 858 2503 862 2507
rect 866 2503 869 2507
rect 869 2503 870 2507
rect 1874 2503 1878 2507
rect 1882 2503 1885 2507
rect 1885 2503 1886 2507
rect 2906 2503 2910 2507
rect 2914 2503 2917 2507
rect 2917 2503 2918 2507
rect 3930 2503 3934 2507
rect 3938 2503 3941 2507
rect 3941 2503 3942 2507
rect 4954 2503 4958 2507
rect 4962 2503 4965 2507
rect 4965 2503 4966 2507
rect 670 2498 674 2502
rect 1798 2498 1802 2502
rect 2142 2498 2146 2502
rect 2182 2498 2186 2502
rect 2238 2498 2242 2502
rect 3038 2498 3042 2502
rect 4022 2498 4026 2502
rect 4190 2498 4194 2502
rect 3286 2488 3290 2492
rect 2678 2478 2682 2482
rect 5086 2478 5090 2482
rect 406 2468 410 2472
rect 1446 2468 1450 2472
rect 1486 2468 1490 2472
rect 1950 2468 1954 2472
rect 2142 2468 2146 2472
rect 3246 2468 3250 2472
rect 1046 2458 1050 2462
rect 1070 2458 1074 2462
rect 1806 2458 1810 2462
rect 3534 2468 3538 2472
rect 3982 2468 3986 2472
rect 4502 2468 4506 2472
rect 5286 2468 5290 2472
rect 1886 2458 1890 2462
rect 1966 2458 1970 2462
rect 2070 2458 2074 2462
rect 278 2448 282 2452
rect 486 2448 490 2452
rect 1310 2448 1314 2452
rect 1318 2448 1322 2452
rect 2014 2448 2018 2452
rect 2310 2448 2314 2452
rect 2670 2448 2674 2452
rect 3534 2448 3538 2452
rect 4398 2448 4402 2452
rect 5126 2448 5130 2452
rect 1038 2438 1042 2442
rect 1590 2438 1594 2442
rect 2510 2438 2514 2442
rect 2622 2438 2626 2442
rect 2982 2438 2986 2442
rect 5086 2438 5090 2442
rect 1766 2428 1770 2432
rect 3326 2428 3330 2432
rect 4190 2428 4194 2432
rect 846 2418 850 2422
rect 2126 2418 2130 2422
rect 2846 2418 2850 2422
rect 5198 2418 5202 2422
rect 14 2408 18 2412
rect 2142 2408 2146 2412
rect 2150 2408 2154 2412
rect 2182 2408 2186 2412
rect 4014 2408 4018 2412
rect 346 2403 350 2407
rect 354 2403 357 2407
rect 357 2403 358 2407
rect 1370 2403 1374 2407
rect 1378 2403 1381 2407
rect 1381 2403 1382 2407
rect 2394 2403 2398 2407
rect 2402 2403 2405 2407
rect 2405 2403 2406 2407
rect 3418 2403 3422 2407
rect 3426 2403 3429 2407
rect 3429 2403 3430 2407
rect 4442 2403 4446 2407
rect 4450 2403 4453 2407
rect 4453 2403 4454 2407
rect 1710 2398 1714 2402
rect 2118 2398 2122 2402
rect 2190 2398 2194 2402
rect 2374 2398 2378 2402
rect 2830 2398 2834 2402
rect 670 2388 674 2392
rect 1486 2388 1490 2392
rect 1822 2388 1826 2392
rect 2606 2388 2610 2392
rect 3342 2388 3346 2392
rect 4318 2388 4322 2392
rect 4822 2388 4826 2392
rect 1054 2378 1058 2382
rect 2382 2378 2386 2382
rect 118 2368 122 2372
rect 1070 2368 1074 2372
rect 1398 2368 1402 2372
rect 1606 2368 1610 2372
rect 3982 2368 3986 2372
rect 5062 2368 5066 2372
rect 646 2358 650 2362
rect 1006 2358 1010 2362
rect 1990 2358 1994 2362
rect 2694 2358 2698 2362
rect 3134 2358 3138 2362
rect 3270 2358 3274 2362
rect 3342 2358 3346 2362
rect 4246 2358 4250 2362
rect 4830 2358 4834 2362
rect 86 2348 90 2352
rect 1462 2348 1466 2352
rect 1494 2348 1498 2352
rect 1758 2348 1762 2352
rect 1814 2348 1818 2352
rect 1846 2348 1850 2352
rect 1902 2348 1906 2352
rect 1942 2348 1946 2352
rect 2214 2348 2218 2352
rect 2246 2348 2250 2352
rect 2510 2348 2514 2352
rect 2830 2348 2834 2352
rect 110 2338 114 2342
rect 174 2338 178 2342
rect 502 2338 506 2342
rect 1550 2338 1554 2342
rect 1630 2338 1634 2342
rect 1718 2338 1722 2342
rect 2198 2338 2202 2342
rect 2350 2338 2354 2342
rect 5078 2348 5082 2352
rect 5214 2348 5218 2352
rect 4710 2338 4714 2342
rect 4798 2338 4802 2342
rect 4838 2338 4842 2342
rect 5006 2338 5010 2342
rect 718 2328 722 2332
rect 902 2328 906 2332
rect 950 2328 954 2332
rect 1190 2328 1194 2332
rect 1870 2328 1874 2332
rect 1886 2328 1890 2332
rect 2030 2328 2034 2332
rect 2046 2328 2050 2332
rect 2190 2328 2194 2332
rect 4054 2328 4058 2332
rect 4942 2328 4946 2332
rect 510 2318 514 2322
rect 526 2318 530 2322
rect 2038 2318 2042 2322
rect 2214 2318 2218 2322
rect 3598 2318 3602 2322
rect 5158 2318 5162 2322
rect 190 2308 194 2312
rect 846 2308 850 2312
rect 1574 2308 1578 2312
rect 1734 2308 1738 2312
rect 2214 2308 2218 2312
rect 2894 2308 2898 2312
rect 3678 2308 3682 2312
rect 3774 2308 3778 2312
rect 4038 2308 4042 2312
rect 182 2298 186 2302
rect 858 2303 862 2307
rect 866 2303 869 2307
rect 869 2303 870 2307
rect 1874 2303 1878 2307
rect 1882 2303 1885 2307
rect 1885 2303 1886 2307
rect 2906 2303 2910 2307
rect 2914 2303 2917 2307
rect 2917 2303 2918 2307
rect 3930 2303 3934 2307
rect 3938 2303 3941 2307
rect 3941 2303 3942 2307
rect 4954 2303 4958 2307
rect 4962 2303 4965 2307
rect 4965 2303 4966 2307
rect 782 2298 786 2302
rect 1726 2298 1730 2302
rect 1742 2298 1746 2302
rect 3078 2298 3082 2302
rect 4894 2298 4898 2302
rect 118 2288 122 2292
rect 806 2288 810 2292
rect 1038 2288 1042 2292
rect 1134 2288 1138 2292
rect 1862 2288 1866 2292
rect 2054 2288 2058 2292
rect 2174 2288 2178 2292
rect 2846 2288 2850 2292
rect 3534 2288 3538 2292
rect 3774 2288 3778 2292
rect 4630 2288 4634 2292
rect 5150 2288 5154 2292
rect 182 2278 186 2282
rect 270 2278 274 2282
rect 1134 2278 1138 2282
rect 1590 2278 1594 2282
rect 1894 2278 1898 2282
rect 2366 2278 2370 2282
rect 4678 2278 4682 2282
rect 4734 2278 4738 2282
rect 5310 2278 5314 2282
rect 54 2268 58 2272
rect 238 2268 242 2272
rect 406 2268 410 2272
rect 470 2268 474 2272
rect 1510 2268 1514 2272
rect 1526 2268 1530 2272
rect 1750 2268 1754 2272
rect 1942 2268 1946 2272
rect 2094 2268 2098 2272
rect 2278 2268 2282 2272
rect 2358 2268 2362 2272
rect 2638 2268 2642 2272
rect 3582 2268 3586 2272
rect 4382 2268 4386 2272
rect 4798 2268 4802 2272
rect 406 2258 410 2262
rect 422 2258 426 2262
rect 958 2258 962 2262
rect 1102 2258 1106 2262
rect 1198 2258 1202 2262
rect 1710 2258 1714 2262
rect 1974 2258 1978 2262
rect 2254 2258 2258 2262
rect 2294 2258 2298 2262
rect 2806 2258 2810 2262
rect 3142 2258 3146 2262
rect 3502 2258 3506 2262
rect 4110 2258 4114 2262
rect 4574 2258 4578 2262
rect 4726 2258 4730 2262
rect 4910 2258 4914 2262
rect 110 2248 114 2252
rect 174 2248 178 2252
rect 422 2248 426 2252
rect 1038 2248 1042 2252
rect 2430 2248 2434 2252
rect 2710 2248 2714 2252
rect 2798 2248 2802 2252
rect 4014 2248 4018 2252
rect 5006 2248 5010 2252
rect 5238 2248 5242 2252
rect 950 2238 954 2242
rect 1334 2238 1338 2242
rect 1638 2238 1642 2242
rect 1646 2238 1650 2242
rect 1734 2238 1738 2242
rect 2126 2238 2130 2242
rect 2318 2238 2322 2242
rect 2854 2238 2858 2242
rect 4286 2238 4290 2242
rect 4382 2238 4386 2242
rect 1638 2228 1642 2232
rect 4390 2228 4394 2232
rect 486 2218 490 2222
rect 1062 2218 1066 2222
rect 3174 2218 3178 2222
rect 4158 2218 4162 2222
rect 5182 2218 5186 2222
rect 1398 2208 1402 2212
rect 1630 2208 1634 2212
rect 1638 2208 1642 2212
rect 2134 2208 2138 2212
rect 2142 2208 2146 2212
rect 2974 2208 2978 2212
rect 4038 2208 4042 2212
rect 346 2203 350 2207
rect 354 2203 357 2207
rect 357 2203 358 2207
rect 1370 2203 1374 2207
rect 1378 2203 1381 2207
rect 1381 2203 1382 2207
rect 14 2198 18 2202
rect 2078 2198 2082 2202
rect 2086 2198 2090 2202
rect 2394 2203 2398 2207
rect 2402 2203 2405 2207
rect 2405 2203 2406 2207
rect 3418 2203 3422 2207
rect 3426 2203 3429 2207
rect 3429 2203 3430 2207
rect 4442 2203 4446 2207
rect 4450 2203 4453 2207
rect 4453 2203 4454 2207
rect 2222 2198 2226 2202
rect 3630 2198 3634 2202
rect 4958 2198 4962 2202
rect 5206 2198 5210 2202
rect 1414 2188 1418 2192
rect 1422 2188 1426 2192
rect 1630 2188 1634 2192
rect 2142 2188 2146 2192
rect 166 2178 170 2182
rect 1478 2178 1482 2182
rect 1638 2178 1642 2182
rect 1958 2178 1962 2182
rect 3534 2178 3538 2182
rect 1670 2168 1674 2172
rect 1862 2168 1866 2172
rect 1990 2168 1994 2172
rect 3438 2168 3442 2172
rect 1622 2158 1626 2162
rect 1686 2158 1690 2162
rect 2054 2158 2058 2162
rect 2990 2158 2994 2162
rect 3574 2158 3578 2162
rect 5198 2158 5202 2162
rect 782 2148 786 2152
rect 1190 2148 1194 2152
rect 1254 2148 1258 2152
rect 1494 2148 1498 2152
rect 1542 2148 1546 2152
rect 1742 2148 1746 2152
rect 2078 2148 2082 2152
rect 2126 2148 2130 2152
rect 2486 2148 2490 2152
rect 2822 2148 2826 2152
rect 2830 2148 2834 2152
rect 3030 2148 3034 2152
rect 3142 2148 3146 2152
rect 3270 2148 3274 2152
rect 3326 2148 3330 2152
rect 3598 2148 3602 2152
rect 3910 2148 3914 2152
rect 5062 2148 5066 2152
rect 5302 2148 5306 2152
rect 1502 2138 1506 2142
rect 1614 2138 1618 2142
rect 2142 2138 2146 2142
rect 2630 2138 2634 2142
rect 2646 2138 2650 2142
rect 2774 2138 2778 2142
rect 2934 2138 2938 2142
rect 1086 2128 1090 2132
rect 1486 2128 1490 2132
rect 1670 2128 1674 2132
rect 1750 2128 1754 2132
rect 2982 2138 2986 2142
rect 3102 2138 3106 2142
rect 4958 2138 4962 2142
rect 5310 2138 5314 2142
rect 2126 2128 2130 2132
rect 2142 2128 2146 2132
rect 2262 2128 2266 2132
rect 2326 2128 2330 2132
rect 2518 2128 2522 2132
rect 2798 2128 2802 2132
rect 3822 2128 3826 2132
rect 102 2118 106 2122
rect 110 2118 114 2122
rect 782 2118 786 2122
rect 998 2118 1002 2122
rect 1086 2118 1090 2122
rect 1998 2118 2002 2122
rect 2294 2118 2298 2122
rect 3462 2118 3466 2122
rect 5302 2128 5306 2132
rect 5358 2128 5362 2132
rect 4902 2118 4906 2122
rect 414 2108 418 2112
rect 1606 2108 1610 2112
rect 1630 2108 1634 2112
rect 1902 2108 1906 2112
rect 2046 2108 2050 2112
rect 2646 2108 2650 2112
rect 3510 2108 3514 2112
rect 4142 2108 4146 2112
rect 4478 2108 4482 2112
rect 4526 2108 4530 2112
rect 858 2103 862 2107
rect 866 2103 869 2107
rect 869 2103 870 2107
rect 1874 2103 1878 2107
rect 1882 2103 1885 2107
rect 1885 2103 1886 2107
rect 2906 2103 2910 2107
rect 2914 2103 2917 2107
rect 2917 2103 2918 2107
rect 3930 2103 3934 2107
rect 3938 2103 3941 2107
rect 3941 2103 3942 2107
rect 4954 2103 4958 2107
rect 4962 2103 4965 2107
rect 4965 2103 4966 2107
rect 478 2098 482 2102
rect 1046 2098 1050 2102
rect 1542 2098 1546 2102
rect 1566 2088 1570 2092
rect 2166 2088 2170 2092
rect 2870 2088 2874 2092
rect 3062 2088 3066 2092
rect 3710 2088 3714 2092
rect 4982 2088 4986 2092
rect 582 2078 586 2082
rect 1742 2078 1746 2082
rect 3406 2078 3410 2082
rect 4374 2078 4378 2082
rect 270 2068 274 2072
rect 310 2068 314 2072
rect 1414 2068 1418 2072
rect 1766 2068 1770 2072
rect 1934 2068 1938 2072
rect 2094 2068 2098 2072
rect 2118 2068 2122 2072
rect 2174 2068 2178 2072
rect 2206 2068 2210 2072
rect 2294 2068 2298 2072
rect 2830 2068 2834 2072
rect 3222 2068 3226 2072
rect 3486 2068 3490 2072
rect 3630 2068 3634 2072
rect 4054 2068 4058 2072
rect 4494 2068 4498 2072
rect 4550 2068 4554 2072
rect 4718 2068 4722 2072
rect 4766 2068 4770 2072
rect 414 2058 418 2062
rect 1246 2058 1250 2062
rect 1334 2058 1338 2062
rect 1470 2058 1474 2062
rect 2070 2058 2074 2062
rect 2822 2058 2826 2062
rect 2974 2058 2978 2062
rect 3294 2058 3298 2062
rect 3982 2058 3986 2062
rect 4238 2058 4242 2062
rect 4342 2058 4346 2062
rect 4406 2058 4410 2062
rect 1662 2048 1666 2052
rect 1870 2048 1874 2052
rect 2062 2048 2066 2052
rect 2182 2048 2186 2052
rect 2510 2048 2514 2052
rect 2622 2048 2626 2052
rect 2782 2048 2786 2052
rect 2790 2048 2794 2052
rect 2814 2048 2818 2052
rect 2854 2048 2858 2052
rect 3222 2048 3226 2052
rect 4798 2048 4802 2052
rect 5310 2048 5314 2052
rect 214 2038 218 2042
rect 1166 2038 1170 2042
rect 1622 2038 1626 2042
rect 1670 2038 1674 2042
rect 1726 2038 1730 2042
rect 2478 2038 2482 2042
rect 3182 2038 3186 2042
rect 3222 2038 3226 2042
rect 5238 2038 5242 2042
rect 238 2028 242 2032
rect 270 2028 274 2032
rect 478 2028 482 2032
rect 1534 2028 1538 2032
rect 4510 2028 4514 2032
rect 4630 2028 4634 2032
rect 5174 2028 5178 2032
rect 422 2018 426 2022
rect 1734 2018 1738 2022
rect 2110 2018 2114 2022
rect 2158 2018 2162 2022
rect 2950 2018 2954 2022
rect 4398 2018 4402 2022
rect 5166 2018 5170 2022
rect 918 2008 922 2012
rect 1566 2008 1570 2012
rect 2142 2008 2146 2012
rect 2558 2008 2562 2012
rect 3246 2008 3250 2012
rect 346 2003 350 2007
rect 354 2003 357 2007
rect 357 2003 358 2007
rect 1370 2003 1374 2007
rect 1378 2003 1381 2007
rect 1381 2003 1382 2007
rect 2394 2003 2398 2007
rect 2402 2003 2405 2007
rect 2405 2003 2406 2007
rect 3418 2003 3422 2007
rect 3426 2003 3429 2007
rect 3429 2003 3430 2007
rect 4442 2003 4446 2007
rect 4450 2003 4453 2007
rect 4453 2003 4454 2007
rect 1622 1998 1626 2002
rect 2526 1998 2530 2002
rect 3438 1998 3442 2002
rect 518 1988 522 1992
rect 4430 1988 4434 1992
rect 4934 1988 4938 1992
rect 5126 1988 5130 1992
rect 294 1978 298 1982
rect 2278 1978 2282 1982
rect 3390 1978 3394 1982
rect 5150 1978 5154 1982
rect 3574 1968 3578 1972
rect 3894 1968 3898 1972
rect 4070 1968 4074 1972
rect 5246 1968 5250 1972
rect 1614 1958 1618 1962
rect 2134 1958 2138 1962
rect 2478 1958 2482 1962
rect 5190 1958 5194 1962
rect 38 1948 42 1952
rect 1982 1948 1986 1952
rect 1998 1948 2002 1952
rect 2774 1948 2778 1952
rect 2998 1948 3002 1952
rect 3022 1948 3026 1952
rect 3870 1948 3874 1952
rect 286 1938 290 1942
rect 478 1938 482 1942
rect 1390 1938 1394 1942
rect 1590 1938 1594 1942
rect 1654 1938 1658 1942
rect 2006 1938 2010 1942
rect 2086 1938 2090 1942
rect 2102 1938 2106 1942
rect 2230 1938 2234 1942
rect 2550 1938 2554 1942
rect 2646 1938 2650 1942
rect 2854 1938 2858 1942
rect 3350 1938 3354 1942
rect 3534 1938 3538 1942
rect 3742 1938 3746 1942
rect 5182 1948 5186 1952
rect 4182 1938 4186 1942
rect 4710 1938 4714 1942
rect 5030 1938 5034 1942
rect 5206 1938 5210 1942
rect 1286 1928 1290 1932
rect 1646 1928 1650 1932
rect 1902 1928 1906 1932
rect 2286 1928 2290 1932
rect 2318 1928 2322 1932
rect 2934 1928 2938 1932
rect 2998 1928 3002 1932
rect 3590 1928 3594 1932
rect 4734 1928 4738 1932
rect 590 1918 594 1922
rect 1694 1918 1698 1922
rect 1822 1918 1826 1922
rect 2390 1918 2394 1922
rect 2622 1918 2626 1922
rect 2798 1918 2802 1922
rect 2942 1918 2946 1922
rect 3086 1918 3090 1922
rect 3310 1918 3314 1922
rect 3582 1918 3586 1922
rect 3710 1918 3714 1922
rect 222 1908 226 1912
rect 910 1908 914 1912
rect 1454 1908 1458 1912
rect 1710 1908 1714 1912
rect 2158 1908 2162 1912
rect 2638 1908 2642 1912
rect 2926 1908 2930 1912
rect 4694 1908 4698 1912
rect 4702 1908 4706 1912
rect 858 1903 862 1907
rect 866 1903 869 1907
rect 869 1903 870 1907
rect 1874 1903 1878 1907
rect 1882 1903 1885 1907
rect 1885 1903 1886 1907
rect 2906 1903 2910 1907
rect 2914 1903 2917 1907
rect 2917 1903 2918 1907
rect 3930 1903 3934 1907
rect 3938 1903 3941 1907
rect 3941 1903 3942 1907
rect 4954 1903 4958 1907
rect 4962 1903 4965 1907
rect 4965 1903 4966 1907
rect 1102 1898 1106 1902
rect 1614 1898 1618 1902
rect 2182 1898 2186 1902
rect 2222 1898 2226 1902
rect 2366 1898 2370 1902
rect 2702 1898 2706 1902
rect 3294 1898 3298 1902
rect 4142 1898 4146 1902
rect 4630 1898 4634 1902
rect 982 1888 986 1892
rect 1622 1888 1626 1892
rect 2302 1888 2306 1892
rect 2430 1888 2434 1892
rect 2622 1888 2626 1892
rect 3078 1888 3082 1892
rect 4358 1888 4362 1892
rect 1494 1878 1498 1882
rect 2174 1878 2178 1882
rect 2422 1878 2426 1882
rect 3174 1878 3178 1882
rect 5150 1878 5154 1882
rect 5190 1878 5194 1882
rect 430 1868 434 1872
rect 694 1868 698 1872
rect 1158 1868 1162 1872
rect 1622 1868 1626 1872
rect 1998 1868 2002 1872
rect 638 1858 642 1862
rect 2278 1868 2282 1872
rect 2286 1868 2290 1872
rect 2766 1868 2770 1872
rect 4158 1868 4162 1872
rect 4302 1868 4306 1872
rect 4822 1868 4826 1872
rect 4894 1868 4898 1872
rect 4910 1868 4914 1872
rect 5014 1868 5018 1872
rect 5022 1868 5026 1872
rect 5126 1868 5130 1872
rect 5254 1868 5258 1872
rect 1550 1858 1554 1862
rect 1926 1858 1930 1862
rect 2142 1858 2146 1862
rect 3078 1858 3082 1862
rect 3702 1858 3706 1862
rect 4350 1858 4354 1862
rect 4638 1858 4642 1862
rect 4798 1858 4802 1862
rect 5006 1858 5010 1862
rect 38 1848 42 1852
rect 542 1848 546 1852
rect 1150 1848 1154 1852
rect 1678 1848 1682 1852
rect 2350 1848 2354 1852
rect 2502 1848 2506 1852
rect 3110 1848 3114 1852
rect 3158 1848 3162 1852
rect 3326 1848 3330 1852
rect 4606 1848 4610 1852
rect 4886 1848 4890 1852
rect 5174 1848 5178 1852
rect 174 1838 178 1842
rect 1310 1838 1314 1842
rect 1358 1838 1362 1842
rect 1670 1838 1674 1842
rect 1942 1838 1946 1842
rect 2014 1838 2018 1842
rect 2126 1838 2130 1842
rect 2294 1838 2298 1842
rect 2646 1838 2650 1842
rect 2830 1838 2834 1842
rect 3014 1838 3018 1842
rect 1454 1828 1458 1832
rect 2638 1828 2642 1832
rect 2854 1828 2858 1832
rect 4406 1828 4410 1832
rect 5206 1828 5210 1832
rect 582 1818 586 1822
rect 1510 1818 1514 1822
rect 1606 1818 1610 1822
rect 1894 1818 1898 1822
rect 2110 1818 2114 1822
rect 4054 1818 4058 1822
rect 4254 1818 4258 1822
rect 3406 1808 3410 1812
rect 4246 1808 4250 1812
rect 346 1803 350 1807
rect 354 1803 357 1807
rect 357 1803 358 1807
rect 1370 1803 1374 1807
rect 1378 1803 1381 1807
rect 1381 1803 1382 1807
rect 2394 1803 2398 1807
rect 2402 1803 2405 1807
rect 2405 1803 2406 1807
rect 3418 1803 3422 1807
rect 3426 1803 3429 1807
rect 3429 1803 3430 1807
rect 4442 1803 4446 1807
rect 4450 1803 4453 1807
rect 4453 1803 4454 1807
rect 878 1798 882 1802
rect 1654 1798 1658 1802
rect 1702 1798 1706 1802
rect 2118 1798 2122 1802
rect 158 1788 162 1792
rect 2494 1788 2498 1792
rect 1174 1778 1178 1782
rect 1894 1778 1898 1782
rect 2078 1778 2082 1782
rect 4526 1778 4530 1782
rect 4750 1778 4754 1782
rect 5198 1778 5202 1782
rect 910 1768 914 1772
rect 1150 1768 1154 1772
rect 1654 1768 1658 1772
rect 2222 1768 2226 1772
rect 2230 1768 2234 1772
rect 2430 1768 2434 1772
rect 2558 1768 2562 1772
rect 3710 1768 3714 1772
rect 5198 1768 5202 1772
rect 894 1758 898 1762
rect 1238 1758 1242 1762
rect 1742 1758 1746 1762
rect 1862 1758 1866 1762
rect 1990 1758 1994 1762
rect 2526 1758 2530 1762
rect 2654 1758 2658 1762
rect 2942 1758 2946 1762
rect 3462 1758 3466 1762
rect 4350 1758 4354 1762
rect 4366 1758 4370 1762
rect 4638 1758 4642 1762
rect 5062 1758 5066 1762
rect 86 1748 90 1752
rect 438 1748 442 1752
rect 494 1748 498 1752
rect 1166 1748 1170 1752
rect 1214 1748 1218 1752
rect 1382 1748 1386 1752
rect 1494 1748 1498 1752
rect 1606 1748 1610 1752
rect 2350 1748 2354 1752
rect 2646 1748 2650 1752
rect 2878 1748 2882 1752
rect 3334 1748 3338 1752
rect 3550 1748 3554 1752
rect 4102 1748 4106 1752
rect 4358 1748 4362 1752
rect 4758 1748 4762 1752
rect 4982 1748 4986 1752
rect 5214 1748 5218 1752
rect 5238 1748 5242 1752
rect 190 1738 194 1742
rect 406 1738 410 1742
rect 502 1738 506 1742
rect 614 1738 618 1742
rect 694 1738 698 1742
rect 1310 1738 1314 1742
rect 1694 1738 1698 1742
rect 2110 1738 2114 1742
rect 2230 1738 2234 1742
rect 2470 1738 2474 1742
rect 534 1728 538 1732
rect 1422 1728 1426 1732
rect 1678 1728 1682 1732
rect 1798 1728 1802 1732
rect 1846 1728 1850 1732
rect 2270 1728 2274 1732
rect 2502 1728 2506 1732
rect 2894 1738 2898 1742
rect 2926 1738 2930 1742
rect 3094 1738 3098 1742
rect 4366 1738 4370 1742
rect 4606 1738 4610 1742
rect 5166 1738 5170 1742
rect 2614 1728 2618 1732
rect 4526 1728 4530 1732
rect 182 1718 186 1722
rect 542 1718 546 1722
rect 1774 1718 1778 1722
rect 1926 1718 1930 1722
rect 2806 1718 2810 1722
rect 5286 1718 5290 1722
rect 926 1708 930 1712
rect 1862 1708 1866 1712
rect 1894 1708 1898 1712
rect 2478 1708 2482 1712
rect 2870 1708 2874 1712
rect 2934 1708 2938 1712
rect 3958 1708 3962 1712
rect 5174 1708 5178 1712
rect 5246 1708 5250 1712
rect 858 1703 862 1707
rect 866 1703 869 1707
rect 869 1703 870 1707
rect 1874 1703 1878 1707
rect 1882 1703 1885 1707
rect 1885 1703 1886 1707
rect 2906 1703 2910 1707
rect 2914 1703 2917 1707
rect 2917 1703 2918 1707
rect 3930 1703 3934 1707
rect 3938 1703 3941 1707
rect 3941 1703 3942 1707
rect 4954 1703 4958 1707
rect 4962 1703 4965 1707
rect 4965 1703 4966 1707
rect 486 1698 490 1702
rect 646 1698 650 1702
rect 1454 1698 1458 1702
rect 1814 1698 1818 1702
rect 1910 1698 1914 1702
rect 2062 1698 2066 1702
rect 2438 1698 2442 1702
rect 2454 1698 2458 1702
rect 3966 1698 3970 1702
rect 5150 1698 5154 1702
rect 5246 1698 5250 1702
rect 494 1688 498 1692
rect 702 1688 706 1692
rect 726 1688 730 1692
rect 902 1688 906 1692
rect 1630 1688 1634 1692
rect 1734 1688 1738 1692
rect 1950 1688 1954 1692
rect 1966 1688 1970 1692
rect 2046 1688 2050 1692
rect 2990 1688 2994 1692
rect 3822 1688 3826 1692
rect 4126 1688 4130 1692
rect 310 1678 314 1682
rect 366 1678 370 1682
rect 694 1678 698 1682
rect 1582 1678 1586 1682
rect 2054 1678 2058 1682
rect 2102 1678 2106 1682
rect 2502 1678 2506 1682
rect 2638 1678 2642 1682
rect 4350 1688 4354 1692
rect 4582 1688 4586 1692
rect 5238 1688 5242 1692
rect 4686 1678 4690 1682
rect 5214 1678 5218 1682
rect 166 1668 170 1672
rect 486 1668 490 1672
rect 766 1668 770 1672
rect 1598 1668 1602 1672
rect 1646 1668 1650 1672
rect 1670 1668 1674 1672
rect 1790 1668 1794 1672
rect 1806 1668 1810 1672
rect 1822 1668 1826 1672
rect 1918 1668 1922 1672
rect 2078 1668 2082 1672
rect 2246 1668 2250 1672
rect 2558 1668 2562 1672
rect 5030 1668 5034 1672
rect 5150 1668 5154 1672
rect 5198 1668 5202 1672
rect 5238 1668 5242 1672
rect 438 1658 442 1662
rect 622 1658 626 1662
rect 854 1658 858 1662
rect 1110 1658 1114 1662
rect 1238 1658 1242 1662
rect 1718 1658 1722 1662
rect 1902 1658 1906 1662
rect 2014 1658 2018 1662
rect 2030 1658 2034 1662
rect 2806 1658 2810 1662
rect 3470 1658 3474 1662
rect 3566 1658 3570 1662
rect 3950 1658 3954 1662
rect 4918 1658 4922 1662
rect 5310 1658 5314 1662
rect 366 1648 370 1652
rect 1622 1648 1626 1652
rect 2510 1648 2514 1652
rect 2750 1648 2754 1652
rect 5014 1648 5018 1652
rect 5174 1648 5178 1652
rect 598 1638 602 1642
rect 750 1638 754 1642
rect 1110 1638 1114 1642
rect 1686 1638 1690 1642
rect 1854 1638 1858 1642
rect 1902 1638 1906 1642
rect 3566 1638 3570 1642
rect 1662 1628 1666 1632
rect 2190 1628 2194 1632
rect 2566 1628 2570 1632
rect 54 1618 58 1622
rect 934 1618 938 1622
rect 1846 1618 1850 1622
rect 1958 1618 1962 1622
rect 2854 1618 2858 1622
rect 974 1608 978 1612
rect 1406 1608 1410 1612
rect 1830 1608 1834 1612
rect 3686 1608 3690 1612
rect 3694 1608 3698 1612
rect 4430 1608 4434 1612
rect 346 1603 350 1607
rect 354 1603 357 1607
rect 357 1603 358 1607
rect 1370 1603 1374 1607
rect 1378 1603 1381 1607
rect 1381 1603 1382 1607
rect 2394 1603 2398 1607
rect 2402 1603 2405 1607
rect 2405 1603 2406 1607
rect 3418 1603 3422 1607
rect 3426 1603 3429 1607
rect 3429 1603 3430 1607
rect 4442 1603 4446 1607
rect 4450 1603 4453 1607
rect 4453 1603 4454 1607
rect 1846 1598 1850 1602
rect 2030 1598 2034 1602
rect 4974 1598 4978 1602
rect 998 1588 1002 1592
rect 1158 1588 1162 1592
rect 1702 1588 1706 1592
rect 2446 1588 2450 1592
rect 2646 1588 2650 1592
rect 94 1578 98 1582
rect 4478 1578 4482 1582
rect 1534 1568 1538 1572
rect 1918 1568 1922 1572
rect 2190 1568 2194 1572
rect 2302 1568 2306 1572
rect 182 1558 186 1562
rect 310 1558 314 1562
rect 1686 1558 1690 1562
rect 1734 1558 1738 1562
rect 1958 1558 1962 1562
rect 3182 1558 3186 1562
rect 430 1548 434 1552
rect 654 1548 658 1552
rect 950 1548 954 1552
rect 998 1548 1002 1552
rect 1750 1548 1754 1552
rect 2278 1548 2282 1552
rect 2286 1548 2290 1552
rect 2678 1548 2682 1552
rect 3022 1548 3026 1552
rect 3526 1548 3530 1552
rect 3974 1548 3978 1552
rect 4014 1548 4018 1552
rect 102 1538 106 1542
rect 478 1538 482 1542
rect 534 1538 538 1542
rect 646 1538 650 1542
rect 718 1538 722 1542
rect 1094 1538 1098 1542
rect 1142 1538 1146 1542
rect 1166 1538 1170 1542
rect 1678 1538 1682 1542
rect 1982 1538 1986 1542
rect 1998 1538 2002 1542
rect 2062 1538 2066 1542
rect 2078 1538 2082 1542
rect 2174 1538 2178 1542
rect 2182 1538 2186 1542
rect 2366 1538 2370 1542
rect 4214 1548 4218 1552
rect 4478 1548 4482 1552
rect 4854 1548 4858 1552
rect 2702 1538 2706 1542
rect 3030 1538 3034 1542
rect 3382 1538 3386 1542
rect 4158 1538 4162 1542
rect 4374 1538 4378 1542
rect 4542 1538 4546 1542
rect 4614 1538 4618 1542
rect 5046 1538 5050 1542
rect 5206 1538 5210 1542
rect 654 1528 658 1532
rect 1494 1528 1498 1532
rect 1894 1528 1898 1532
rect 1950 1528 1954 1532
rect 2054 1528 2058 1532
rect 2094 1528 2098 1532
rect 3334 1528 3338 1532
rect 4438 1528 4442 1532
rect 4638 1528 4642 1532
rect 734 1518 738 1522
rect 838 1518 842 1522
rect 2006 1518 2010 1522
rect 2038 1518 2042 1522
rect 3190 1518 3194 1522
rect 3726 1518 3730 1522
rect 4710 1518 4714 1522
rect 4790 1518 4794 1522
rect 5182 1518 5186 1522
rect 5302 1518 5306 1522
rect 190 1508 194 1512
rect 502 1508 506 1512
rect 846 1508 850 1512
rect 2150 1508 2154 1512
rect 2782 1508 2786 1512
rect 4342 1508 4346 1512
rect 5166 1508 5170 1512
rect 858 1503 862 1507
rect 866 1503 869 1507
rect 869 1503 870 1507
rect 1874 1503 1878 1507
rect 1882 1503 1885 1507
rect 1885 1503 1886 1507
rect 2906 1503 2910 1507
rect 2914 1503 2917 1507
rect 2917 1503 2918 1507
rect 3930 1503 3934 1507
rect 3938 1503 3941 1507
rect 3941 1503 3942 1507
rect 4954 1503 4958 1507
rect 4962 1503 4965 1507
rect 4965 1503 4966 1507
rect 94 1498 98 1502
rect 1862 1498 1866 1502
rect 2190 1498 2194 1502
rect 2198 1498 2202 1502
rect 2414 1498 2418 1502
rect 2606 1498 2610 1502
rect 3974 1498 3978 1502
rect 710 1488 714 1492
rect 846 1488 850 1492
rect 1126 1488 1130 1492
rect 1766 1488 1770 1492
rect 1926 1488 1930 1492
rect 2014 1488 2018 1492
rect 2022 1488 2026 1492
rect 2190 1488 2194 1492
rect 3510 1488 3514 1492
rect 4254 1488 4258 1492
rect 5302 1488 5306 1492
rect 246 1478 250 1482
rect 494 1478 498 1482
rect 734 1478 738 1482
rect 1558 1478 1562 1482
rect 1982 1478 1986 1482
rect 2246 1478 2250 1482
rect 2486 1478 2490 1482
rect 2742 1478 2746 1482
rect 3294 1478 3298 1482
rect 3894 1478 3898 1482
rect 4582 1478 4586 1482
rect 5134 1478 5138 1482
rect 5190 1478 5194 1482
rect 174 1468 178 1472
rect 1342 1468 1346 1472
rect 1566 1468 1570 1472
rect 1862 1468 1866 1472
rect 1998 1468 2002 1472
rect 2030 1468 2034 1472
rect 2278 1468 2282 1472
rect 3918 1468 3922 1472
rect 4662 1468 4666 1472
rect 4982 1468 4986 1472
rect 862 1458 866 1462
rect 1022 1458 1026 1462
rect 1102 1458 1106 1462
rect 1190 1458 1194 1462
rect 1302 1458 1306 1462
rect 1518 1458 1522 1462
rect 1702 1458 1706 1462
rect 1750 1458 1754 1462
rect 2006 1458 2010 1462
rect 2086 1458 2090 1462
rect 2462 1458 2466 1462
rect 2782 1458 2786 1462
rect 2958 1458 2962 1462
rect 3958 1458 3962 1462
rect 4198 1458 4202 1462
rect 5030 1458 5034 1462
rect 5310 1458 5314 1462
rect 1318 1448 1322 1452
rect 1782 1448 1786 1452
rect 1814 1448 1818 1452
rect 1934 1448 1938 1452
rect 2046 1448 2050 1452
rect 2134 1448 2138 1452
rect 2742 1448 2746 1452
rect 3702 1448 3706 1452
rect 222 1438 226 1442
rect 806 1438 810 1442
rect 1902 1438 1906 1442
rect 3502 1438 3506 1442
rect 3790 1438 3794 1442
rect 4326 1438 4330 1442
rect 382 1428 386 1432
rect 534 1428 538 1432
rect 1390 1428 1394 1432
rect 1766 1428 1770 1432
rect 1902 1428 1906 1432
rect 1942 1428 1946 1432
rect 2310 1428 2314 1432
rect 3462 1428 3466 1432
rect 4638 1428 4642 1432
rect 958 1418 962 1422
rect 1822 1418 1826 1422
rect 1918 1418 1922 1422
rect 2214 1418 2218 1422
rect 2534 1418 2538 1422
rect 1158 1408 1162 1412
rect 2142 1408 2146 1412
rect 5190 1408 5194 1412
rect 346 1403 350 1407
rect 354 1403 357 1407
rect 357 1403 358 1407
rect 1370 1403 1374 1407
rect 1378 1403 1381 1407
rect 1381 1403 1382 1407
rect 2394 1403 2398 1407
rect 2402 1403 2405 1407
rect 2405 1403 2406 1407
rect 3418 1403 3422 1407
rect 3426 1403 3429 1407
rect 3429 1403 3430 1407
rect 4442 1403 4446 1407
rect 4450 1403 4453 1407
rect 4453 1403 4454 1407
rect 1462 1398 1466 1402
rect 1550 1388 1554 1392
rect 2958 1388 2962 1392
rect 2974 1388 2978 1392
rect 3310 1388 3314 1392
rect 4862 1388 4866 1392
rect 486 1378 490 1382
rect 542 1378 546 1382
rect 1894 1378 1898 1382
rect 1006 1368 1010 1372
rect 1118 1368 1122 1372
rect 1182 1368 1186 1372
rect 1806 1368 1810 1372
rect 4198 1368 4202 1372
rect 1054 1358 1058 1362
rect 1734 1358 1738 1362
rect 2126 1358 2130 1362
rect 2190 1358 2194 1362
rect 2206 1358 2210 1362
rect 2222 1358 2226 1362
rect 2622 1358 2626 1362
rect 3534 1358 3538 1362
rect 1006 1348 1010 1352
rect 1166 1348 1170 1352
rect 1614 1348 1618 1352
rect 1766 1348 1770 1352
rect 2150 1348 2154 1352
rect 2254 1348 2258 1352
rect 2278 1348 2282 1352
rect 3206 1348 3210 1352
rect 3518 1348 3522 1352
rect 3542 1348 3546 1352
rect 750 1338 754 1342
rect 1094 1338 1098 1342
rect 1790 1338 1794 1342
rect 1814 1338 1818 1342
rect 1870 1338 1874 1342
rect 2102 1338 2106 1342
rect 2230 1338 2234 1342
rect 2422 1338 2426 1342
rect 2526 1338 2530 1342
rect 2550 1338 2554 1342
rect 2998 1338 3002 1342
rect 4294 1348 4298 1352
rect 4630 1348 4634 1352
rect 4902 1348 4906 1352
rect 5030 1348 5034 1352
rect 5158 1348 5162 1352
rect 3678 1338 3682 1342
rect 4398 1338 4402 1342
rect 478 1328 482 1332
rect 1310 1328 1314 1332
rect 4790 1338 4794 1342
rect 2110 1328 2114 1332
rect 2230 1328 2234 1332
rect 2374 1328 2378 1332
rect 2390 1328 2394 1332
rect 2542 1328 2546 1332
rect 3494 1328 3498 1332
rect 1270 1318 1274 1322
rect 1494 1318 1498 1322
rect 1686 1318 1690 1322
rect 1926 1318 1930 1322
rect 1974 1318 1978 1322
rect 2134 1318 2138 1322
rect 2366 1318 2370 1322
rect 2382 1318 2386 1322
rect 2590 1318 2594 1322
rect 3374 1318 3378 1322
rect 4702 1318 4706 1322
rect 4742 1318 4746 1322
rect 414 1308 418 1312
rect 1798 1308 1802 1312
rect 1846 1308 1850 1312
rect 2190 1308 2194 1312
rect 2462 1308 2466 1312
rect 858 1303 862 1307
rect 866 1303 869 1307
rect 869 1303 870 1307
rect 542 1298 546 1302
rect 1350 1298 1354 1302
rect 1874 1303 1878 1307
rect 1882 1303 1885 1307
rect 1885 1303 1886 1307
rect 1734 1298 1738 1302
rect 2906 1303 2910 1307
rect 2914 1303 2917 1307
rect 2917 1303 2918 1307
rect 3930 1303 3934 1307
rect 3938 1303 3941 1307
rect 3941 1303 3942 1307
rect 4954 1303 4958 1307
rect 4962 1303 4965 1307
rect 4965 1303 4966 1307
rect 3558 1298 3562 1302
rect 5230 1298 5234 1302
rect 1022 1288 1026 1292
rect 1598 1288 1602 1292
rect 2470 1288 2474 1292
rect 3950 1288 3954 1292
rect 4214 1288 4218 1292
rect 5022 1288 5026 1292
rect 1246 1278 1250 1282
rect 1342 1278 1346 1282
rect 1550 1278 1554 1282
rect 1670 1278 1674 1282
rect 1910 1278 1914 1282
rect 1982 1278 1986 1282
rect 2150 1278 2154 1282
rect 2174 1278 2178 1282
rect 3918 1278 3922 1282
rect 4510 1278 4514 1282
rect 5238 1278 5242 1282
rect 5246 1278 5250 1282
rect 1406 1268 1410 1272
rect 1782 1268 1786 1272
rect 1822 1268 1826 1272
rect 1838 1268 1842 1272
rect 1886 1268 1890 1272
rect 2174 1268 2178 1272
rect 2790 1268 2794 1272
rect 3078 1268 3082 1272
rect 3310 1268 3314 1272
rect 5062 1268 5066 1272
rect 374 1258 378 1262
rect 798 1258 802 1262
rect 1246 1258 1250 1262
rect 1550 1258 1554 1262
rect 1606 1258 1610 1262
rect 1702 1258 1706 1262
rect 1790 1258 1794 1262
rect 1798 1258 1802 1262
rect 1918 1258 1922 1262
rect 2134 1258 2138 1262
rect 2174 1258 2178 1262
rect 2278 1258 2282 1262
rect 2334 1258 2338 1262
rect 2558 1258 2562 1262
rect 2998 1258 3002 1262
rect 3398 1258 3402 1262
rect 4198 1258 4202 1262
rect 4294 1258 4298 1262
rect 4902 1258 4906 1262
rect 5238 1258 5242 1262
rect 366 1248 370 1252
rect 862 1248 866 1252
rect 1758 1248 1762 1252
rect 2310 1248 2314 1252
rect 3494 1248 3498 1252
rect 4574 1248 4578 1252
rect 4662 1248 4666 1252
rect 5054 1248 5058 1252
rect 822 1238 826 1242
rect 1814 1238 1818 1242
rect 2790 1238 2794 1242
rect 2902 1238 2906 1242
rect 5038 1238 5042 1242
rect 5070 1238 5074 1242
rect 926 1228 930 1232
rect 1510 1228 1514 1232
rect 1766 1228 1770 1232
rect 2222 1228 2226 1232
rect 5054 1228 5058 1232
rect 838 1218 842 1222
rect 878 1218 882 1222
rect 1974 1218 1978 1222
rect 3702 1218 3706 1222
rect 4878 1218 4882 1222
rect 5158 1218 5162 1222
rect 334 1208 338 1212
rect 2958 1208 2962 1212
rect 3390 1208 3394 1212
rect 5222 1208 5226 1212
rect 346 1203 350 1207
rect 354 1203 357 1207
rect 357 1203 358 1207
rect 1370 1203 1374 1207
rect 1378 1203 1381 1207
rect 1381 1203 1382 1207
rect 2394 1203 2398 1207
rect 2402 1203 2405 1207
rect 2405 1203 2406 1207
rect 3418 1203 3422 1207
rect 3426 1203 3429 1207
rect 3429 1203 3430 1207
rect 4442 1203 4446 1207
rect 4450 1203 4453 1207
rect 4453 1203 4454 1207
rect 1598 1198 1602 1202
rect 2870 1198 2874 1202
rect 3094 1198 3098 1202
rect 334 1188 338 1192
rect 574 1188 578 1192
rect 1094 1188 1098 1192
rect 1102 1188 1106 1192
rect 2030 1188 2034 1192
rect 2966 1188 2970 1192
rect 4014 1188 4018 1192
rect 2142 1178 2146 1182
rect 3966 1178 3970 1182
rect 1254 1168 1258 1172
rect 2086 1168 2090 1172
rect 4102 1168 4106 1172
rect 4238 1168 4242 1172
rect 4270 1168 4274 1172
rect 398 1158 402 1162
rect 422 1158 426 1162
rect 1214 1158 1218 1162
rect 1246 1158 1250 1162
rect 1502 1158 1506 1162
rect 1678 1158 1682 1162
rect 1846 1158 1850 1162
rect 2038 1158 2042 1162
rect 2294 1158 2298 1162
rect 4238 1158 4242 1162
rect 5310 1158 5314 1162
rect 542 1148 546 1152
rect 1022 1148 1026 1152
rect 2886 1148 2890 1152
rect 958 1138 962 1142
rect 1342 1138 1346 1142
rect 4102 1148 4106 1152
rect 4742 1148 4746 1152
rect 1934 1138 1938 1142
rect 1982 1138 1986 1142
rect 2302 1138 2306 1142
rect 166 1128 170 1132
rect 406 1128 410 1132
rect 574 1128 578 1132
rect 1238 1128 1242 1132
rect 1462 1128 1466 1132
rect 1846 1128 1850 1132
rect 1990 1128 1994 1132
rect 2030 1128 2034 1132
rect 2102 1128 2106 1132
rect 2862 1128 2866 1132
rect 3462 1128 3466 1132
rect 950 1118 954 1122
rect 1550 1118 1554 1122
rect 1798 1118 1802 1122
rect 2254 1118 2258 1122
rect 3502 1118 3506 1122
rect 3734 1118 3738 1122
rect 4886 1118 4890 1122
rect 1990 1108 1994 1112
rect 1998 1108 2002 1112
rect 3406 1108 3410 1112
rect 858 1103 862 1107
rect 866 1103 869 1107
rect 869 1103 870 1107
rect 1874 1103 1878 1107
rect 1882 1103 1885 1107
rect 1885 1103 1886 1107
rect 2906 1103 2910 1107
rect 2914 1103 2917 1107
rect 2917 1103 2918 1107
rect 3930 1103 3934 1107
rect 3938 1103 3941 1107
rect 3941 1103 3942 1107
rect 4954 1103 4958 1107
rect 4962 1103 4965 1107
rect 4965 1103 4966 1107
rect 374 1098 378 1102
rect 3950 1098 3954 1102
rect 4582 1098 4586 1102
rect 4622 1098 4626 1102
rect 222 1088 226 1092
rect 550 1088 554 1092
rect 1454 1088 1458 1092
rect 1910 1088 1914 1092
rect 5006 1088 5010 1092
rect 70 1078 74 1082
rect 710 1078 714 1082
rect 1646 1078 1650 1082
rect 1974 1078 1978 1082
rect 2382 1078 2386 1082
rect 4022 1078 4026 1082
rect 5310 1078 5314 1082
rect 598 1068 602 1072
rect 742 1068 746 1072
rect 822 1068 826 1072
rect 1806 1068 1810 1072
rect 1998 1068 2002 1072
rect 2294 1068 2298 1072
rect 382 1058 386 1062
rect 1774 1058 1778 1062
rect 3214 1068 3218 1072
rect 3734 1068 3738 1072
rect 1974 1058 1978 1062
rect 2662 1058 2666 1062
rect 4742 1058 4746 1062
rect 4910 1058 4914 1062
rect 5022 1058 5026 1062
rect 5078 1058 5082 1062
rect 742 1048 746 1052
rect 934 1048 938 1052
rect 1734 1048 1738 1052
rect 2774 1048 2778 1052
rect 2862 1048 2866 1052
rect 2982 1048 2986 1052
rect 950 1038 954 1042
rect 2598 1038 2602 1042
rect 2942 1028 2946 1032
rect 510 1018 514 1022
rect 558 1018 562 1022
rect 2166 1018 2170 1022
rect 1510 1008 1514 1012
rect 1518 1008 1522 1012
rect 1614 1008 1618 1012
rect 2230 1008 2234 1012
rect 2382 1008 2386 1012
rect 5030 1008 5034 1012
rect 346 1003 350 1007
rect 354 1003 357 1007
rect 357 1003 358 1007
rect 1370 1003 1374 1007
rect 1378 1003 1381 1007
rect 1381 1003 1382 1007
rect 2394 1003 2398 1007
rect 2402 1003 2405 1007
rect 2405 1003 2406 1007
rect 3418 1003 3422 1007
rect 3426 1003 3429 1007
rect 3429 1003 3430 1007
rect 4442 1003 4446 1007
rect 4450 1003 4453 1007
rect 4453 1003 4454 1007
rect 2086 998 2090 1002
rect 3110 998 3114 1002
rect 1134 988 1138 992
rect 1310 988 1314 992
rect 1550 988 1554 992
rect 4238 988 4242 992
rect 1462 978 1466 982
rect 78 968 82 972
rect 406 968 410 972
rect 1574 968 1578 972
rect 2542 968 2546 972
rect 4390 968 4394 972
rect 5206 968 5210 972
rect 366 958 370 962
rect 510 958 514 962
rect 1366 958 1370 962
rect 2510 958 2514 962
rect 5238 958 5242 962
rect 798 948 802 952
rect 934 948 938 952
rect 1038 948 1042 952
rect 1094 948 1098 952
rect 1390 948 1394 952
rect 1422 948 1426 952
rect 1518 948 1522 952
rect 2030 948 2034 952
rect 2334 948 2338 952
rect 2342 948 2346 952
rect 2534 948 2538 952
rect 2614 948 2618 952
rect 2622 948 2626 952
rect 3470 948 3474 952
rect 4222 948 4226 952
rect 5198 948 5202 952
rect 5310 948 5314 952
rect 1574 938 1578 942
rect 1622 938 1626 942
rect 2174 938 2178 942
rect 2334 938 2338 942
rect 2710 938 2714 942
rect 4390 938 4394 942
rect 5230 938 5234 942
rect 1798 928 1802 932
rect 2094 928 2098 932
rect 2750 928 2754 932
rect 4166 928 4170 932
rect 5174 928 5178 932
rect 1470 918 1474 922
rect 1726 918 1730 922
rect 1966 918 1970 922
rect 2054 918 2058 922
rect 2086 918 2090 922
rect 1158 908 1162 912
rect 2286 908 2290 912
rect 2622 908 2626 912
rect 2870 908 2874 912
rect 4126 908 4130 912
rect 858 903 862 907
rect 866 903 869 907
rect 869 903 870 907
rect 1874 903 1878 907
rect 1882 903 1885 907
rect 1885 903 1886 907
rect 2906 903 2910 907
rect 2914 903 2917 907
rect 2917 903 2918 907
rect 3930 903 3934 907
rect 3938 903 3941 907
rect 3941 903 3942 907
rect 2062 898 2066 902
rect 2078 898 2082 902
rect 3326 898 3330 902
rect 4954 903 4958 907
rect 4962 903 4965 907
rect 4965 903 4966 907
rect 542 888 546 892
rect 734 888 738 892
rect 750 888 754 892
rect 1358 888 1362 892
rect 1662 888 1666 892
rect 3038 888 3042 892
rect 6 878 10 882
rect 302 878 306 882
rect 550 878 554 882
rect 558 878 562 882
rect 734 878 738 882
rect 1126 878 1130 882
rect 1262 878 1266 882
rect 1926 878 1930 882
rect 2142 878 2146 882
rect 2598 878 2602 882
rect 3022 878 3026 882
rect 3118 878 3122 882
rect 3766 878 3770 882
rect 5302 878 5306 882
rect 1414 868 1418 872
rect 1542 868 1546 872
rect 1662 868 1666 872
rect 2350 868 2354 872
rect 2590 868 2594 872
rect 2638 868 2642 872
rect 3486 868 3490 872
rect 5054 868 5058 872
rect 5246 868 5250 872
rect 302 858 306 862
rect 1126 858 1130 862
rect 1550 858 1554 862
rect 1758 858 1762 862
rect 1806 858 1810 862
rect 1910 858 1914 862
rect 1990 858 1994 862
rect 2342 858 2346 862
rect 2382 858 2386 862
rect 2470 858 2474 862
rect 3326 858 3330 862
rect 3470 858 3474 862
rect 5126 858 5130 862
rect 5302 858 5306 862
rect 958 848 962 852
rect 1310 848 1314 852
rect 2142 848 2146 852
rect 2158 848 2162 852
rect 614 838 618 842
rect 662 838 666 842
rect 1158 838 1162 842
rect 1742 838 1746 842
rect 1902 838 1906 842
rect 4622 838 4626 842
rect 1654 828 1658 832
rect 1790 828 1794 832
rect 2046 828 2050 832
rect 2054 828 2058 832
rect 2926 828 2930 832
rect 1046 818 1050 822
rect 2278 818 2282 822
rect 3742 818 3746 822
rect 4574 818 4578 822
rect 1238 808 1242 812
rect 1950 808 1954 812
rect 4126 808 4130 812
rect 346 803 350 807
rect 354 803 357 807
rect 357 803 358 807
rect 1370 803 1374 807
rect 1378 803 1381 807
rect 1381 803 1382 807
rect 2394 803 2398 807
rect 2402 803 2405 807
rect 2405 803 2406 807
rect 3418 803 3422 807
rect 3426 803 3429 807
rect 3429 803 3430 807
rect 4442 803 4446 807
rect 4450 803 4453 807
rect 4453 803 4454 807
rect 2446 798 2450 802
rect 2926 798 2930 802
rect 4766 798 4770 802
rect 3718 788 3722 792
rect 1926 778 1930 782
rect 1510 768 1514 772
rect 1534 768 1538 772
rect 1726 768 1730 772
rect 2062 768 2066 772
rect 5150 768 5154 772
rect 3054 758 3058 762
rect 4606 758 4610 762
rect 5094 758 5098 762
rect 6 748 10 752
rect 230 748 234 752
rect 326 748 330 752
rect 798 748 802 752
rect 1270 748 1274 752
rect 1454 748 1458 752
rect 1478 748 1482 752
rect 1574 748 1578 752
rect 2790 748 2794 752
rect 3102 748 3106 752
rect 3510 748 3514 752
rect 4198 748 4202 752
rect 4678 748 4682 752
rect 5206 748 5210 752
rect 654 738 658 742
rect 662 738 666 742
rect 1030 738 1034 742
rect 2366 738 2370 742
rect 2454 738 2458 742
rect 3054 738 3058 742
rect 3526 738 3530 742
rect 3582 738 3586 742
rect 3998 738 4002 742
rect 4022 738 4026 742
rect 5166 738 5170 742
rect 430 728 434 732
rect 550 728 554 732
rect 1318 728 1322 732
rect 1470 728 1474 732
rect 1478 728 1482 732
rect 1494 728 1498 732
rect 1614 728 1618 732
rect 2470 728 2474 732
rect 2510 728 2514 732
rect 3326 728 3330 732
rect 558 718 562 722
rect 1014 718 1018 722
rect 1622 718 1626 722
rect 1846 718 1850 722
rect 1918 718 1922 722
rect 2086 718 2090 722
rect 3254 718 3258 722
rect 4942 718 4946 722
rect 1502 708 1506 712
rect 1862 708 1866 712
rect 2214 708 2218 712
rect 2430 708 2434 712
rect 2806 708 2810 712
rect 2814 708 2818 712
rect 858 703 862 707
rect 866 703 869 707
rect 869 703 870 707
rect 1874 703 1878 707
rect 1882 703 1885 707
rect 1885 703 1886 707
rect 2906 703 2910 707
rect 2914 703 2917 707
rect 2917 703 2918 707
rect 3930 703 3934 707
rect 3938 703 3941 707
rect 3941 703 3942 707
rect 4954 703 4958 707
rect 4962 703 4965 707
rect 4965 703 4966 707
rect 254 698 258 702
rect 1014 698 1018 702
rect 2622 698 2626 702
rect 4550 698 4554 702
rect 1070 688 1074 692
rect 1294 688 1298 692
rect 1302 688 1306 692
rect 2046 688 2050 692
rect 2118 688 2122 692
rect 2678 688 2682 692
rect 2790 688 2794 692
rect 3166 688 3170 692
rect 4262 688 4266 692
rect 4486 688 4490 692
rect 5254 688 5258 692
rect 2942 678 2946 682
rect 5142 678 5146 682
rect 190 668 194 672
rect 382 668 386 672
rect 1502 668 1506 672
rect 1662 668 1666 672
rect 1830 668 1834 672
rect 1862 668 1866 672
rect 3214 668 3218 672
rect 3958 668 3962 672
rect 4262 668 4266 672
rect 4574 668 4578 672
rect 5190 668 5194 672
rect 1646 658 1650 662
rect 2038 658 2042 662
rect 3326 658 3330 662
rect 4030 658 4034 662
rect 342 648 346 652
rect 534 648 538 652
rect 2950 648 2954 652
rect 4022 648 4026 652
rect 4318 648 4322 652
rect 326 638 330 642
rect 1614 638 1618 642
rect 2966 638 2970 642
rect 3558 638 3562 642
rect 950 628 954 632
rect 1318 628 1322 632
rect 1942 628 1946 632
rect 2574 628 2578 632
rect 2662 628 2666 632
rect 2934 628 2938 632
rect 1310 618 1314 622
rect 1926 618 1930 622
rect 2758 618 2762 622
rect 5214 618 5218 622
rect 526 608 530 612
rect 1454 608 1458 612
rect 1598 608 1602 612
rect 2006 608 2010 612
rect 346 603 350 607
rect 354 603 357 607
rect 357 603 358 607
rect 1370 603 1374 607
rect 1378 603 1381 607
rect 1381 603 1382 607
rect 2394 603 2398 607
rect 2402 603 2405 607
rect 2405 603 2406 607
rect 3418 603 3422 607
rect 3426 603 3429 607
rect 3429 603 3430 607
rect 4442 603 4446 607
rect 4450 603 4453 607
rect 4453 603 4454 607
rect 1086 598 1090 602
rect 1094 598 1098 602
rect 1494 598 1498 602
rect 1614 598 1618 602
rect 1758 598 1762 602
rect 2110 598 2114 602
rect 2934 598 2938 602
rect 2942 598 2946 602
rect 3342 598 3346 602
rect 982 588 986 592
rect 1302 588 1306 592
rect 1598 578 1602 582
rect 2798 578 2802 582
rect 1086 568 1090 572
rect 2038 568 2042 572
rect 2094 568 2098 572
rect 2198 568 2202 572
rect 3614 568 3618 572
rect 3966 568 3970 572
rect 4174 568 4178 572
rect 1230 558 1234 562
rect 1406 558 1410 562
rect 3982 558 3986 562
rect 318 548 322 552
rect 710 548 714 552
rect 1030 548 1034 552
rect 1494 548 1498 552
rect 2102 548 2106 552
rect 2254 548 2258 552
rect 5254 548 5258 552
rect 1302 538 1306 542
rect 2950 538 2954 542
rect 3438 538 3442 542
rect 3470 538 3474 542
rect 5054 538 5058 542
rect 5270 538 5274 542
rect 5302 538 5306 542
rect 806 528 810 532
rect 886 528 890 532
rect 1022 528 1026 532
rect 2798 528 2802 532
rect 3838 528 3842 532
rect 4054 528 4058 532
rect 118 518 122 522
rect 1302 518 1306 522
rect 2878 518 2882 522
rect 858 503 862 507
rect 866 503 869 507
rect 869 503 870 507
rect 1874 503 1878 507
rect 1882 503 1885 507
rect 1885 503 1886 507
rect 2906 503 2910 507
rect 2914 503 2917 507
rect 2917 503 2918 507
rect 3930 503 3934 507
rect 3938 503 3941 507
rect 3941 503 3942 507
rect 4954 503 4958 507
rect 4962 503 4965 507
rect 4965 503 4966 507
rect 38 498 42 502
rect 2094 498 2098 502
rect 2190 498 2194 502
rect 2382 498 2386 502
rect 2766 498 2770 502
rect 2934 498 2938 502
rect 4262 498 4266 502
rect 230 488 234 492
rect 1294 488 1298 492
rect 1998 488 2002 492
rect 2182 488 2186 492
rect 2230 488 2234 492
rect 2022 478 2026 482
rect 2758 478 2762 482
rect 2766 478 2770 482
rect 3350 478 3354 482
rect 5070 478 5074 482
rect 398 468 402 472
rect 1342 468 1346 472
rect 550 458 554 462
rect 2014 468 2018 472
rect 2334 468 2338 472
rect 2350 468 2354 472
rect 2414 468 2418 472
rect 3214 468 3218 472
rect 1182 458 1186 462
rect 1454 458 1458 462
rect 2526 458 2530 462
rect 2678 458 2682 462
rect 3678 468 3682 472
rect 3758 468 3762 472
rect 4870 468 4874 472
rect 5062 468 5066 472
rect 2894 458 2898 462
rect 3006 458 3010 462
rect 3254 458 3258 462
rect 3550 458 3554 462
rect 3646 458 3650 462
rect 3838 458 3842 462
rect 4934 458 4938 462
rect 2070 448 2074 452
rect 2558 448 2562 452
rect 3470 448 3474 452
rect 1142 428 1146 432
rect 2678 428 2682 432
rect 2798 428 2802 432
rect 4054 428 4058 432
rect 1078 418 1082 422
rect 1582 418 1586 422
rect 2630 418 2634 422
rect 3438 418 3442 422
rect 526 408 530 412
rect 2014 408 2018 412
rect 3918 408 3922 412
rect 4614 408 4618 412
rect 346 403 350 407
rect 354 403 357 407
rect 357 403 358 407
rect 1370 403 1374 407
rect 1378 403 1381 407
rect 1381 403 1382 407
rect 2394 403 2398 407
rect 2402 403 2405 407
rect 2405 403 2406 407
rect 3418 403 3422 407
rect 3426 403 3429 407
rect 3429 403 3430 407
rect 4442 403 4446 407
rect 4450 403 4453 407
rect 4453 403 4454 407
rect 398 388 402 392
rect 2694 388 2698 392
rect 2974 388 2978 392
rect 3366 388 3370 392
rect 4086 388 4090 392
rect 2758 378 2762 382
rect 4342 378 4346 382
rect 758 368 762 372
rect 1150 368 1154 372
rect 2222 368 2226 372
rect 2854 368 2858 372
rect 3182 368 3186 372
rect 5262 368 5266 372
rect 2934 358 2938 362
rect 3334 358 3338 362
rect 4614 358 4618 362
rect 5270 358 5274 362
rect 62 348 66 352
rect 38 338 42 342
rect 502 348 506 352
rect 1102 348 1106 352
rect 1510 348 1514 352
rect 1526 348 1530 352
rect 1606 348 1610 352
rect 1894 348 1898 352
rect 2038 348 2042 352
rect 2078 348 2082 352
rect 3094 348 3098 352
rect 3438 348 3442 352
rect 846 338 850 342
rect 1142 338 1146 342
rect 1430 338 1434 342
rect 2158 338 2162 342
rect 2398 338 2402 342
rect 3102 338 3106 342
rect 3294 338 3298 342
rect 5278 338 5282 342
rect 1606 328 1610 332
rect 2478 328 2482 332
rect 3734 328 3738 332
rect 4102 328 4106 332
rect 3606 318 3610 322
rect 5310 318 5314 322
rect 1286 308 1290 312
rect 3590 308 3594 312
rect 4142 308 4146 312
rect 858 303 862 307
rect 866 303 869 307
rect 869 303 870 307
rect 1874 303 1878 307
rect 1882 303 1885 307
rect 1885 303 1886 307
rect 2906 303 2910 307
rect 2914 303 2917 307
rect 2917 303 2918 307
rect 3930 303 3934 307
rect 3938 303 3941 307
rect 3941 303 3942 307
rect 4954 303 4958 307
rect 4962 303 4965 307
rect 4965 303 4966 307
rect 1246 298 1250 302
rect 1254 298 1258 302
rect 1326 298 1330 302
rect 3470 298 3474 302
rect 3478 298 3482 302
rect 4022 298 4026 302
rect 4078 298 4082 302
rect 5206 298 5210 302
rect 3246 288 3250 292
rect 4230 288 4234 292
rect 4334 288 4338 292
rect 2222 278 2226 282
rect 2246 278 2250 282
rect 2358 278 2362 282
rect 2758 278 2762 282
rect 3294 278 3298 282
rect 3790 278 3794 282
rect 526 268 530 272
rect 878 268 882 272
rect 1086 268 1090 272
rect 1270 268 1274 272
rect 1326 268 1330 272
rect 1526 268 1530 272
rect 1542 268 1546 272
rect 1598 268 1602 272
rect 2262 268 2266 272
rect 3998 268 4002 272
rect 1254 258 1258 262
rect 1398 258 1402 262
rect 2150 258 2154 262
rect 2382 258 2386 262
rect 3078 258 3082 262
rect 3230 258 3234 262
rect 4558 258 4562 262
rect 3374 248 3378 252
rect 3470 248 3474 252
rect 4174 248 4178 252
rect 5278 248 5282 252
rect 1270 238 1274 242
rect 2622 238 2626 242
rect 3174 238 3178 242
rect 2494 228 2498 232
rect 2014 218 2018 222
rect 2622 218 2626 222
rect 1502 208 1506 212
rect 2094 208 2098 212
rect 346 203 350 207
rect 354 203 357 207
rect 357 203 358 207
rect 1370 203 1374 207
rect 1378 203 1381 207
rect 1381 203 1382 207
rect 2394 203 2398 207
rect 2402 203 2405 207
rect 2405 203 2406 207
rect 3418 203 3422 207
rect 3426 203 3429 207
rect 3429 203 3430 207
rect 4442 203 4446 207
rect 4450 203 4453 207
rect 4453 203 4454 207
rect 334 198 338 202
rect 1518 198 1522 202
rect 1526 198 1530 202
rect 2174 198 2178 202
rect 3438 198 3442 202
rect 1222 188 1226 192
rect 1694 188 1698 192
rect 1790 188 1794 192
rect 1998 188 2002 192
rect 4102 188 4106 192
rect 5286 188 5290 192
rect 3102 168 3106 172
rect 3150 168 3154 172
rect 3854 168 3858 172
rect 118 158 122 162
rect 1662 158 1666 162
rect 2734 158 2738 162
rect 2846 158 2850 162
rect 2950 158 2954 162
rect 4094 158 4098 162
rect 4342 158 4346 162
rect 4422 158 4426 162
rect 494 148 498 152
rect 542 148 546 152
rect 662 148 666 152
rect 614 138 618 142
rect 1310 148 1314 152
rect 2206 148 2210 152
rect 5206 148 5210 152
rect 5302 148 5306 152
rect 1294 138 1298 142
rect 1574 138 1578 142
rect 1798 138 1802 142
rect 2382 138 2386 142
rect 2478 138 2482 142
rect 2534 138 2538 142
rect 2854 138 2858 142
rect 2990 138 2994 142
rect 4046 138 4050 142
rect 5246 138 5250 142
rect 1222 128 1226 132
rect 1438 128 1442 132
rect 1870 128 1874 132
rect 2126 128 2130 132
rect 2174 128 2178 132
rect 2206 128 2210 132
rect 2830 128 2834 132
rect 3070 128 3074 132
rect 3086 128 3090 132
rect 3350 128 3354 132
rect 3398 128 3402 132
rect 4142 118 4146 122
rect 838 108 842 112
rect 846 108 850 112
rect 1502 108 1506 112
rect 1790 108 1794 112
rect 2094 108 2098 112
rect 858 103 862 107
rect 866 103 869 107
rect 869 103 870 107
rect 262 98 266 102
rect 1342 98 1346 102
rect 1874 103 1878 107
rect 1882 103 1885 107
rect 1885 103 1886 107
rect 2906 103 2910 107
rect 2914 103 2917 107
rect 2917 103 2918 107
rect 3930 103 3934 107
rect 3938 103 3941 107
rect 3941 103 3942 107
rect 4954 103 4958 107
rect 4962 103 4965 107
rect 4965 103 4966 107
rect 1894 98 1898 102
rect 2518 98 2522 102
rect 3262 98 3266 102
rect 3270 98 3274 102
rect 3918 98 3922 102
rect 4102 98 4106 102
rect 758 88 762 92
rect 3062 88 3066 92
rect 3854 88 3858 92
rect 3982 88 3986 92
rect 4262 88 4266 92
rect 4550 88 4554 92
rect 510 78 514 82
rect 534 78 538 82
rect 838 78 842 82
rect 942 78 946 82
rect 1126 78 1130 82
rect 2750 78 2754 82
rect 2790 78 2794 82
rect 3350 78 3354 82
rect 3358 78 3362 82
rect 5302 78 5306 82
rect 542 68 546 72
rect 958 68 962 72
rect 1286 68 1290 72
rect 1478 68 1482 72
rect 1910 68 1914 72
rect 2230 68 2234 72
rect 2446 68 2450 72
rect 2494 68 2498 72
rect 2814 68 2818 72
rect 2942 68 2946 72
rect 3350 68 3354 72
rect 3366 68 3370 72
rect 3414 68 3418 72
rect 3574 68 3578 72
rect 3614 68 3618 72
rect 3622 68 3626 72
rect 398 58 402 62
rect 734 58 738 62
rect 1046 58 1050 62
rect 1438 58 1442 62
rect 1478 58 1482 62
rect 2022 58 2026 62
rect 2158 58 2162 62
rect 5294 68 5298 72
rect 2254 58 2258 62
rect 2318 58 2322 62
rect 3254 58 3258 62
rect 3654 58 3658 62
rect 262 48 266 52
rect 990 48 994 52
rect 5262 48 5266 52
rect 2038 38 2042 42
rect 2750 38 2754 42
rect 3150 38 3154 42
rect 1230 28 1234 32
rect 2046 28 2050 32
rect 2182 28 2186 32
rect 526 18 530 22
rect 558 18 562 22
rect 798 18 802 22
rect 1078 18 1082 22
rect 1278 18 1282 22
rect 1390 18 1394 22
rect 2070 18 2074 22
rect 2150 18 2154 22
rect 2198 18 2202 22
rect 2558 18 2562 22
rect 2926 18 2930 22
rect 3182 18 3186 22
rect 3558 18 3562 22
rect 3718 18 3722 22
rect 4094 18 4098 22
rect 4486 18 4490 22
rect 502 8 506 12
rect 1102 8 1106 12
rect 1182 8 1186 12
rect 1214 8 1218 12
rect 1310 8 1314 12
rect 1350 8 1354 12
rect 1454 8 1458 12
rect 1494 8 1498 12
rect 1646 8 1650 12
rect 1686 8 1690 12
rect 1742 8 1746 12
rect 1806 8 1810 12
rect 2030 8 2034 12
rect 2102 8 2106 12
rect 2190 8 2194 12
rect 2254 8 2258 12
rect 2350 8 2354 12
rect 2414 8 2418 12
rect 2974 8 2978 12
rect 3014 8 3018 12
rect 3094 8 3098 12
rect 3334 8 3338 12
rect 3510 8 3514 12
rect 4054 8 4058 12
rect 4198 8 4202 12
rect 4430 8 4434 12
rect 5238 8 5242 12
rect 346 3 350 7
rect 354 3 357 7
rect 357 3 358 7
rect 1370 3 1374 7
rect 1378 3 1381 7
rect 1381 3 1382 7
rect 2394 3 2398 7
rect 2402 3 2405 7
rect 2405 3 2406 7
rect 3418 3 3422 7
rect 3426 3 3429 7
rect 3429 3 3430 7
rect 4442 3 4446 7
rect 4450 3 4453 7
rect 4453 3 4454 7
<< metal4 >>
rect 856 3703 858 3707
rect 862 3703 865 3707
rect 870 3703 872 3707
rect 1872 3703 1874 3707
rect 1878 3703 1881 3707
rect 1886 3703 1888 3707
rect 2904 3703 2906 3707
rect 2910 3703 2913 3707
rect 2918 3703 2920 3707
rect 3928 3703 3930 3707
rect 3934 3703 3937 3707
rect 3942 3703 3944 3707
rect 4952 3703 4954 3707
rect 4958 3703 4961 3707
rect 4966 3703 4968 3707
rect 3994 3698 4001 3701
rect 4074 3698 4081 3701
rect 4210 3698 4217 3701
rect 4370 3698 4377 3701
rect 942 3672 945 3678
rect 970 3668 974 3671
rect 1362 3668 1366 3671
rect 1206 3662 1209 3668
rect 1734 3662 1737 3688
rect 1978 3678 1982 3681
rect 344 3603 346 3607
rect 350 3603 353 3607
rect 358 3603 360 3607
rect 438 3532 441 3548
rect 54 3388 62 3391
rect 14 2912 17 3258
rect 54 2922 57 3388
rect 118 3271 121 3388
rect 118 3268 126 3271
rect 166 2792 169 3528
rect 178 3238 185 3241
rect 182 3122 185 3238
rect 230 3022 233 3338
rect 254 2902 257 3458
rect 344 3403 346 3407
rect 350 3403 353 3407
rect 358 3403 360 3407
rect 344 3203 346 3207
rect 350 3203 353 3207
rect 358 3203 360 3207
rect 406 3102 409 3338
rect 422 3262 425 3498
rect 446 3462 449 3558
rect 486 3378 494 3381
rect 462 3322 465 3368
rect 486 3332 489 3378
rect 530 3368 534 3371
rect 586 3368 590 3371
rect 438 3172 441 3218
rect 422 3122 425 3138
rect 454 3082 457 3108
rect 344 3003 346 3007
rect 350 3003 353 3007
rect 358 3003 360 3007
rect 478 2992 481 3238
rect 486 3162 489 3298
rect 366 2922 369 2948
rect 344 2803 346 2807
rect 350 2803 353 2807
rect 358 2803 360 2807
rect 18 2608 22 2611
rect 14 2412 17 2548
rect 110 2521 113 2598
rect 138 2538 142 2541
rect 150 2532 153 2688
rect 166 2642 169 2668
rect 344 2603 346 2607
rect 350 2603 353 2607
rect 358 2603 360 2607
rect 366 2592 369 2918
rect 502 2912 505 3238
rect 562 3138 566 3141
rect 574 3062 577 3138
rect 606 3112 609 3338
rect 614 3308 622 3311
rect 614 3112 617 3308
rect 630 3142 633 3348
rect 646 3332 649 3428
rect 686 3342 689 3398
rect 706 3368 713 3371
rect 638 3132 641 3138
rect 646 3122 649 3328
rect 710 3292 713 3368
rect 670 3072 673 3118
rect 542 2928 550 2931
rect 398 2712 401 2858
rect 414 2552 417 2828
rect 202 2538 206 2541
rect 110 2518 118 2521
rect 430 2512 433 2858
rect 542 2632 545 2928
rect 662 2742 665 2948
rect 670 2832 673 3068
rect 686 2842 689 3138
rect 742 2902 745 3558
rect 1094 3542 1097 3548
rect 856 3503 858 3507
rect 862 3503 865 3507
rect 870 3503 872 3507
rect 750 3142 753 3468
rect 782 3272 785 3338
rect 810 3288 814 3291
rect 782 2942 785 3268
rect 782 2752 785 2938
rect 502 2538 510 2541
rect 270 2448 278 2451
rect 18 2198 22 2201
rect 54 2072 57 2268
rect 38 1852 41 1948
rect 54 1622 57 2068
rect 86 1752 89 2348
rect 118 2341 121 2368
rect 114 2338 121 2341
rect 102 2122 105 2128
rect 110 2122 113 2248
rect 118 2212 121 2288
rect 174 2252 177 2338
rect 182 2282 185 2298
rect 190 2292 193 2308
rect 270 2282 273 2448
rect 344 2403 346 2407
rect 350 2403 353 2407
rect 358 2403 360 2407
rect 158 2178 166 2181
rect 158 1792 161 2178
rect 174 1842 177 2248
rect 182 1722 185 2278
rect 406 2272 409 2468
rect 474 2268 481 2271
rect 218 2038 225 2041
rect 222 1912 225 2038
rect 238 2032 241 2268
rect 406 2262 409 2268
rect 344 2203 346 2207
rect 350 2203 353 2207
rect 358 2203 360 2207
rect 306 2068 310 2071
rect 270 2032 273 2068
rect 344 2003 346 2007
rect 350 2003 353 2007
rect 358 2003 360 2007
rect 294 1941 297 1978
rect 290 1938 297 1941
rect 344 1803 346 1807
rect 350 1803 353 1807
rect 358 1803 360 1807
rect 94 1502 97 1578
rect 102 1542 105 1558
rect 166 1132 169 1668
rect 178 1558 182 1561
rect 190 1512 193 1738
rect 366 1682 369 2118
rect 406 1742 409 2258
rect 422 2252 425 2258
rect 414 2062 417 2108
rect 422 2022 425 2248
rect 478 2102 481 2268
rect 486 2222 489 2448
rect 494 2162 497 2528
rect 502 2342 505 2538
rect 526 2322 529 2628
rect 630 2562 633 2578
rect 662 2552 665 2558
rect 678 2522 681 2678
rect 670 2392 673 2498
rect 646 2362 649 2368
rect 710 2322 713 2748
rect 718 2332 721 2728
rect 514 2318 521 2321
rect 478 1942 481 2028
rect 518 1992 521 2318
rect 790 2301 793 3258
rect 838 3072 841 3098
rect 846 2992 849 3358
rect 942 3312 945 3338
rect 856 3303 858 3307
rect 862 3303 865 3307
rect 870 3303 872 3307
rect 950 3302 953 3308
rect 906 3298 910 3301
rect 958 3292 961 3308
rect 902 3252 905 3258
rect 856 3103 858 3107
rect 862 3103 865 3107
rect 870 3103 872 3107
rect 918 3072 921 3198
rect 966 3162 969 3338
rect 974 3022 977 3418
rect 1142 3402 1145 3648
rect 1150 3552 1153 3558
rect 1022 3352 1025 3358
rect 1070 3322 1073 3358
rect 982 3298 990 3301
rect 982 3122 985 3298
rect 1066 3288 1070 3291
rect 1042 3258 1046 3261
rect 862 2922 865 2948
rect 856 2903 858 2907
rect 862 2903 865 2907
rect 870 2903 872 2907
rect 856 2703 858 2707
rect 862 2703 865 2707
rect 870 2703 872 2707
rect 786 2298 793 2301
rect 806 2292 809 2658
rect 858 2558 862 2561
rect 856 2503 858 2507
rect 862 2503 865 2507
rect 870 2503 872 2507
rect 846 2312 849 2418
rect 856 2303 858 2307
rect 862 2303 865 2307
rect 870 2303 872 2307
rect 782 2122 785 2148
rect 856 2103 858 2107
rect 862 2103 865 2107
rect 870 2103 872 2107
rect 310 1562 313 1678
rect 366 1652 369 1678
rect 344 1603 346 1607
rect 350 1603 353 1607
rect 358 1603 360 1607
rect 430 1552 433 1868
rect 438 1662 441 1748
rect 486 1672 489 1698
rect 494 1692 497 1748
rect 250 1478 254 1481
rect 174 1472 177 1478
rect 222 1092 225 1438
rect 344 1403 346 1407
rect 350 1403 353 1407
rect 358 1403 360 1407
rect 334 1192 337 1208
rect 344 1203 346 1207
rect 350 1203 353 1207
rect 358 1203 360 1207
rect 74 1078 81 1081
rect 78 972 81 1078
rect 344 1003 346 1007
rect 350 1003 353 1007
rect 358 1003 360 1007
rect 366 962 369 1248
rect 374 1102 377 1258
rect 382 1062 385 1428
rect 478 1332 481 1538
rect 486 1382 489 1668
rect 494 1482 497 1688
rect 502 1512 505 1738
rect 534 1732 537 1748
rect 542 1722 545 1848
rect 582 1822 585 2078
rect 594 1918 601 1921
rect 598 1642 601 1918
rect 856 1903 858 1907
rect 862 1903 865 1907
rect 870 1903 872 1907
rect 642 1858 646 1861
rect 694 1742 697 1868
rect 878 1802 881 2958
rect 1006 2932 1009 2948
rect 886 2712 889 2738
rect 902 2572 905 2858
rect 902 2332 905 2358
rect 894 1762 897 2018
rect 910 1912 913 2798
rect 974 2712 977 2748
rect 986 2678 990 2681
rect 998 2592 1001 2678
rect 1006 2362 1009 2858
rect 1058 2678 1062 2681
rect 1078 2652 1081 2948
rect 1086 2668 1094 2671
rect 1086 2642 1089 2668
rect 1118 2582 1121 2738
rect 1126 2662 1129 2688
rect 1126 2612 1129 2638
rect 1070 2462 1073 2548
rect 1034 2438 1038 2441
rect 950 2242 953 2328
rect 1034 2288 1038 2291
rect 958 2242 961 2258
rect 1030 2248 1038 2251
rect 1030 2192 1033 2248
rect 922 2008 929 2011
rect 914 1768 918 1771
rect 534 1432 537 1538
rect 406 1161 409 1168
rect 402 1158 409 1161
rect 414 1161 417 1308
rect 542 1302 545 1378
rect 546 1298 553 1301
rect 414 1158 422 1161
rect 406 972 409 1128
rect 510 962 513 1018
rect 542 892 545 1148
rect 550 1092 553 1298
rect 574 1132 577 1188
rect 594 1068 598 1071
rect 6 882 9 888
rect 558 882 561 1018
rect 546 878 550 881
rect 302 862 305 878
rect 614 842 617 1738
rect 926 1712 929 2008
rect 856 1703 858 1707
rect 862 1703 865 1707
rect 870 1703 872 1707
rect 626 1658 630 1661
rect 646 1542 649 1698
rect 698 1688 702 1691
rect 898 1688 902 1691
rect 686 1678 694 1681
rect 686 1662 689 1678
rect 654 1532 657 1548
rect 726 1541 729 1688
rect 766 1662 769 1668
rect 722 1538 729 1541
rect 714 1488 718 1491
rect 734 1482 737 1518
rect 750 1342 753 1638
rect 854 1612 857 1658
rect 810 1438 814 1441
rect 802 1258 806 1261
rect 710 1072 713 1078
rect 822 1072 825 1238
rect 838 1222 841 1518
rect 846 1492 849 1508
rect 856 1503 858 1507
rect 862 1503 865 1507
rect 870 1503 872 1507
rect 866 1458 870 1461
rect 856 1303 858 1307
rect 862 1303 865 1307
rect 870 1303 872 1307
rect 862 1252 865 1258
rect 926 1232 929 1708
rect 856 1103 858 1107
rect 862 1103 865 1107
rect 870 1103 872 1107
rect 742 1052 745 1068
rect 802 948 806 951
rect 856 903 858 907
rect 862 903 865 907
rect 870 903 872 907
rect 746 888 750 891
rect 734 882 737 888
rect 6 752 9 818
rect 344 803 346 807
rect 350 803 353 807
rect 358 803 360 807
rect 190 652 193 668
rect 38 342 41 498
rect 62 352 65 358
rect 118 162 121 518
rect 230 492 233 748
rect 254 662 257 698
rect 326 642 329 748
rect 434 728 438 731
rect 386 668 393 671
rect 390 652 393 668
rect 338 648 342 651
rect 344 603 346 607
rect 350 603 353 607
rect 358 603 360 607
rect 322 548 326 551
rect 344 403 346 407
rect 350 403 353 407
rect 358 403 360 407
rect 398 392 401 468
rect 334 202 337 338
rect 344 203 346 207
rect 350 203 353 207
rect 358 203 360 207
rect 262 52 265 98
rect 398 62 401 388
rect 502 352 505 778
rect 662 742 665 838
rect 798 752 801 758
rect 654 732 657 738
rect 546 728 550 731
rect 558 692 561 718
rect 534 652 537 658
rect 526 412 529 608
rect 710 532 713 548
rect 554 458 558 461
rect 490 148 494 151
rect 502 12 505 348
rect 514 78 518 81
rect 526 22 529 268
rect 534 148 542 151
rect 534 142 537 148
rect 534 72 537 78
rect 542 72 545 78
rect 558 22 561 458
rect 658 148 662 151
rect 610 138 614 141
rect 758 92 761 368
rect 738 58 742 61
rect 798 22 801 748
rect 856 703 858 707
rect 862 703 865 707
rect 870 703 872 707
rect 806 532 809 538
rect 856 503 858 507
rect 862 503 865 507
rect 870 503 872 507
rect 846 112 849 338
rect 856 303 858 307
rect 862 303 865 307
rect 870 303 872 307
rect 878 272 881 1218
rect 934 1052 937 1618
rect 970 1608 974 1611
rect 946 1548 950 1551
rect 958 1142 961 1418
rect 950 1042 953 1118
rect 934 952 937 958
rect 950 848 958 851
rect 950 632 953 848
rect 982 592 985 1888
rect 998 1592 1001 2118
rect 1046 2102 1049 2458
rect 1058 2378 1065 2381
rect 1062 2222 1065 2378
rect 1070 2362 1073 2368
rect 1134 2292 1137 2768
rect 1174 2702 1177 3458
rect 1182 3362 1185 3368
rect 1182 3322 1185 3328
rect 1190 3302 1193 3538
rect 1198 3352 1201 3468
rect 1254 3352 1257 3358
rect 1274 3348 1278 3351
rect 1198 2942 1201 3348
rect 1258 3288 1262 3291
rect 1210 3068 1214 3071
rect 1218 3048 1222 3051
rect 1230 2891 1233 3058
rect 1322 3048 1326 3051
rect 1230 2888 1238 2891
rect 1294 2832 1297 2948
rect 1334 2792 1337 3608
rect 1368 3603 1370 3607
rect 1374 3603 1377 3607
rect 1382 3603 1384 3607
rect 1358 3552 1361 3598
rect 1368 3403 1370 3407
rect 1374 3403 1377 3407
rect 1382 3403 1384 3407
rect 1370 3338 1374 3341
rect 1350 3332 1353 3338
rect 1422 3322 1425 3658
rect 1506 3648 1510 3651
rect 1626 3648 1630 3651
rect 1466 3348 1470 3351
rect 1458 3328 1462 3331
rect 1410 3318 1414 3321
rect 1368 3203 1370 3207
rect 1374 3203 1377 3207
rect 1382 3203 1384 3207
rect 1368 3003 1370 3007
rect 1374 3003 1377 3007
rect 1382 3003 1384 3007
rect 1406 2892 1409 3098
rect 1478 3002 1481 3548
rect 1538 3438 1542 3441
rect 1510 3132 1513 3148
rect 1518 2992 1521 3328
rect 1526 3132 1529 3238
rect 1368 2803 1370 2807
rect 1374 2803 1377 2807
rect 1382 2803 1384 2807
rect 1390 2612 1393 2848
rect 1368 2603 1370 2607
rect 1374 2603 1377 2607
rect 1382 2603 1384 2607
rect 1310 2452 1313 2528
rect 1318 2452 1321 2518
rect 1334 2512 1337 2528
rect 1368 2403 1370 2407
rect 1374 2403 1377 2407
rect 1382 2403 1384 2407
rect 1394 2368 1398 2371
rect 1102 2232 1105 2258
rect 1090 2128 1094 2131
rect 1082 2118 1086 2121
rect 998 1542 1001 1548
rect 1090 1538 1094 1541
rect 1102 1462 1105 1898
rect 1110 1642 1113 1658
rect 1122 1488 1126 1491
rect 1006 1352 1009 1368
rect 1022 1292 1025 1458
rect 1118 1362 1121 1368
rect 1058 1358 1062 1361
rect 1022 1152 1025 1288
rect 1094 1192 1097 1338
rect 1038 952 1041 958
rect 1046 822 1049 858
rect 1014 702 1017 718
rect 1030 552 1033 738
rect 1074 688 1078 691
rect 1094 602 1097 948
rect 1086 572 1089 598
rect 890 528 894 531
rect 1026 528 1030 531
rect 838 82 841 108
rect 856 103 858 107
rect 862 103 865 107
rect 870 103 872 107
rect 946 78 953 81
rect 950 72 953 78
rect 962 68 966 71
rect 1046 62 1049 68
rect 990 52 993 58
rect 1078 22 1081 418
rect 1102 352 1105 1188
rect 1134 992 1137 2278
rect 1190 2152 1193 2328
rect 1150 1852 1153 1858
rect 1146 1768 1150 1771
rect 1158 1592 1161 1868
rect 1166 1752 1169 2038
rect 1142 1542 1145 1548
rect 1158 1412 1161 1588
rect 1174 1541 1177 1778
rect 1170 1538 1177 1541
rect 1198 1492 1201 2258
rect 1334 2172 1337 2238
rect 1368 2203 1370 2207
rect 1374 2203 1377 2207
rect 1382 2203 1384 2207
rect 1258 2148 1262 2151
rect 1338 2058 1342 2061
rect 1246 2042 1249 2058
rect 1368 2003 1370 2007
rect 1374 2003 1377 2007
rect 1382 2003 1384 2007
rect 1286 1872 1289 1928
rect 1310 1792 1313 1838
rect 1214 1752 1217 1758
rect 1238 1752 1241 1758
rect 1190 1462 1193 1478
rect 1170 1348 1174 1351
rect 1126 862 1129 878
rect 1158 842 1161 908
rect 1182 462 1185 1368
rect 1238 1161 1241 1658
rect 1302 1462 1305 1468
rect 1310 1332 1313 1738
rect 1338 1468 1342 1471
rect 1318 1442 1321 1448
rect 1246 1262 1249 1278
rect 1258 1168 1262 1171
rect 1238 1158 1246 1161
rect 1090 268 1094 271
rect 1102 12 1105 348
rect 1142 342 1145 428
rect 1138 338 1142 341
rect 1150 332 1153 368
rect 1130 78 1134 81
rect 1182 12 1185 458
rect 1214 12 1217 1158
rect 1238 812 1241 1128
rect 1262 872 1265 878
rect 1270 752 1273 1318
rect 1342 1282 1345 1288
rect 1338 1138 1342 1141
rect 1310 852 1313 988
rect 1274 748 1281 751
rect 1222 132 1225 188
rect 1222 62 1225 128
rect 1230 32 1233 558
rect 1242 298 1246 301
rect 1254 262 1257 298
rect 1270 242 1273 268
rect 1278 22 1281 748
rect 1294 672 1297 688
rect 1302 592 1305 688
rect 1318 632 1321 728
rect 1302 522 1305 538
rect 1286 72 1289 308
rect 1294 142 1297 488
rect 1310 152 1313 618
rect 1322 298 1326 301
rect 1322 268 1326 271
rect 1310 12 1313 148
rect 1342 102 1345 468
rect 1350 12 1353 1298
rect 1358 892 1361 1838
rect 1368 1803 1370 1807
rect 1374 1803 1377 1807
rect 1382 1803 1384 1807
rect 1382 1742 1385 1748
rect 1368 1603 1370 1607
rect 1374 1603 1377 1607
rect 1382 1603 1384 1607
rect 1390 1432 1393 1938
rect 1368 1403 1370 1407
rect 1374 1403 1377 1407
rect 1382 1403 1384 1407
rect 1368 1203 1370 1207
rect 1374 1203 1377 1207
rect 1382 1203 1384 1207
rect 1368 1003 1370 1007
rect 1374 1003 1377 1007
rect 1382 1003 1384 1007
rect 1366 942 1369 958
rect 1398 952 1401 2208
rect 1422 2192 1425 2918
rect 1446 2472 1449 2728
rect 1486 2392 1489 2468
rect 1462 2352 1465 2358
rect 1414 2072 1417 2188
rect 1474 2178 1478 2181
rect 1486 2132 1489 2388
rect 1518 2352 1521 2748
rect 1526 2512 1529 2718
rect 1498 2348 1505 2351
rect 1462 2058 1470 2061
rect 1446 1911 1449 1968
rect 1446 1908 1454 1911
rect 1406 1462 1409 1608
rect 1410 1268 1414 1271
rect 1422 952 1425 1728
rect 1454 1702 1457 1828
rect 1462 1402 1465 2058
rect 1494 1882 1497 2148
rect 1502 2142 1505 2348
rect 1510 1822 1513 2268
rect 1494 1732 1497 1748
rect 1494 1322 1497 1528
rect 1518 1462 1521 2348
rect 1462 1132 1465 1138
rect 1458 1088 1465 1091
rect 1462 982 1465 1088
rect 1368 803 1370 807
rect 1374 803 1377 807
rect 1382 803 1384 807
rect 1368 603 1370 607
rect 1374 603 1377 607
rect 1382 603 1384 607
rect 1368 403 1370 407
rect 1374 403 1377 407
rect 1382 403 1384 407
rect 1368 203 1370 207
rect 1374 203 1377 207
rect 1382 203 1384 207
rect 1390 22 1393 948
rect 1410 868 1414 871
rect 1458 748 1462 751
rect 1470 732 1473 918
rect 1478 732 1481 748
rect 1406 562 1409 618
rect 1454 462 1457 608
rect 1494 602 1497 728
rect 1502 712 1505 1158
rect 1510 1012 1513 1228
rect 1518 952 1521 1008
rect 1526 782 1529 2268
rect 1542 2142 1545 2148
rect 1542 2102 1545 2138
rect 1534 1572 1537 2028
rect 1550 1862 1553 2338
rect 1566 2092 1569 3228
rect 1574 2888 1582 2891
rect 1574 2312 1577 2888
rect 1606 2862 1609 3098
rect 1614 3092 1617 3648
rect 1742 3642 1745 3678
rect 1790 3672 1793 3678
rect 1674 3478 1681 3481
rect 1678 3452 1681 3478
rect 1702 3442 1705 3448
rect 1714 3438 1718 3441
rect 1670 3332 1673 3338
rect 1702 3332 1705 3338
rect 1710 3302 1713 3348
rect 1678 3278 1686 3281
rect 1678 3272 1681 3278
rect 1718 3092 1721 3368
rect 1770 3338 1774 3341
rect 1646 2772 1649 2778
rect 1586 2438 1590 2441
rect 1606 2372 1609 2588
rect 1594 2278 1598 2281
rect 1606 2112 1609 2368
rect 1614 2142 1617 2738
rect 1654 2582 1657 2948
rect 1678 2542 1681 2828
rect 1630 2332 1633 2338
rect 1646 2242 1649 2538
rect 1634 2238 1638 2241
rect 1638 2212 1641 2228
rect 1630 2192 1633 2208
rect 1622 2042 1625 2158
rect 1630 2112 1633 2158
rect 1550 1392 1553 1858
rect 1558 1482 1561 1688
rect 1566 1472 1569 2008
rect 1550 1262 1553 1278
rect 1550 992 1553 1118
rect 1542 862 1545 868
rect 1550 862 1553 988
rect 1574 942 1577 968
rect 1514 768 1518 771
rect 1530 768 1534 771
rect 1570 748 1574 751
rect 1502 672 1505 708
rect 1426 338 1430 341
rect 1398 192 1401 258
rect 1442 128 1446 131
rect 1442 58 1446 61
rect 1454 12 1457 458
rect 1478 62 1481 68
rect 1494 12 1497 548
rect 1582 422 1585 1678
rect 1590 792 1593 1938
rect 1614 1902 1617 1958
rect 1622 1892 1625 1998
rect 1606 1752 1609 1818
rect 1598 1292 1601 1668
rect 1622 1652 1625 1868
rect 1598 1202 1601 1288
rect 1606 1262 1609 1318
rect 1614 1012 1617 1348
rect 1614 642 1617 728
rect 1622 722 1625 938
rect 1598 582 1601 608
rect 1614 602 1617 638
rect 1630 552 1633 1688
rect 1638 822 1641 2178
rect 1670 2172 1673 2508
rect 1670 2052 1673 2128
rect 1646 1761 1649 1928
rect 1654 1802 1657 1938
rect 1654 1772 1657 1798
rect 1646 1758 1657 1761
rect 1646 1672 1649 1678
rect 1646 662 1649 1078
rect 1654 832 1657 1758
rect 1662 1632 1665 2048
rect 1670 1842 1673 2038
rect 1678 1852 1681 2538
rect 1686 2152 1689 2158
rect 1694 1922 1697 2258
rect 1702 1842 1705 2528
rect 1710 2402 1713 2948
rect 1718 2712 1721 3058
rect 1710 1962 1713 2258
rect 1678 1732 1681 1838
rect 1670 1282 1673 1668
rect 1686 1562 1689 1638
rect 1678 1542 1681 1548
rect 1686 1322 1689 1558
rect 1662 872 1665 888
rect 1662 672 1665 868
rect 1514 348 1521 351
rect 1502 112 1505 208
rect 1518 202 1521 348
rect 1526 342 1529 348
rect 1606 332 1609 348
rect 1546 268 1550 271
rect 1594 268 1598 271
rect 1526 202 1529 268
rect 1578 138 1582 141
rect 1646 12 1649 658
rect 1654 158 1662 161
rect 1654 152 1657 158
rect 1678 11 1681 1158
rect 1694 1152 1697 1738
rect 1702 1592 1705 1798
rect 1710 1522 1713 1908
rect 1718 1662 1721 2338
rect 1726 2302 1729 2428
rect 1734 2312 1737 2688
rect 1734 2242 1737 2308
rect 1742 2302 1745 3278
rect 1790 3182 1793 3668
rect 1838 3472 1841 3488
rect 1846 3482 1849 3638
rect 1862 3532 1865 3548
rect 1872 3503 1874 3507
rect 1878 3503 1881 3507
rect 1886 3503 1888 3507
rect 1806 3261 1809 3318
rect 1802 3258 1809 3261
rect 1750 2592 1753 3108
rect 1766 2792 1769 2858
rect 1798 2502 1801 2728
rect 1814 2702 1817 3338
rect 1872 3303 1874 3307
rect 1878 3303 1881 3307
rect 1886 3303 1888 3307
rect 1872 3103 1874 3107
rect 1878 3103 1881 3107
rect 1886 3103 1888 3107
rect 1822 3038 1830 3041
rect 1822 2592 1825 3038
rect 1766 2432 1769 2438
rect 1806 2362 1809 2458
rect 1822 2392 1825 2548
rect 1746 2268 1750 2271
rect 1742 2082 1745 2148
rect 1706 1458 1710 1461
rect 1726 1442 1729 2038
rect 1734 2022 1737 2038
rect 1738 1758 1742 1761
rect 1734 1562 1737 1688
rect 1750 1572 1753 2128
rect 1734 1362 1737 1558
rect 1750 1552 1753 1568
rect 1742 1458 1750 1461
rect 1734 1302 1737 1358
rect 1702 1252 1705 1258
rect 1726 772 1729 918
rect 1694 142 1697 188
rect 1678 8 1686 11
rect 1734 11 1737 1048
rect 1742 842 1745 1458
rect 1758 1252 1761 2348
rect 1766 2062 1769 2068
rect 1766 1482 1769 1488
rect 1766 1352 1769 1428
rect 1766 1232 1769 1348
rect 1774 1062 1777 1718
rect 1790 1672 1793 1718
rect 1798 1642 1801 1728
rect 1806 1672 1809 2358
rect 1818 2348 1825 2351
rect 1822 1922 1825 2348
rect 1782 1392 1785 1448
rect 1790 1342 1793 1518
rect 1790 1292 1793 1338
rect 1798 1312 1801 1638
rect 1814 1452 1817 1698
rect 1822 1422 1825 1668
rect 1830 1612 1833 2718
rect 1838 2348 1846 2351
rect 1838 1392 1841 2348
rect 1846 1622 1849 1728
rect 1854 1642 1857 3058
rect 1872 2903 1874 2907
rect 1878 2903 1881 2907
rect 1886 2903 1888 2907
rect 1872 2703 1874 2707
rect 1878 2703 1881 2707
rect 1886 2703 1888 2707
rect 1894 2701 1897 2758
rect 1894 2698 1902 2701
rect 1894 2512 1897 2648
rect 1872 2503 1874 2507
rect 1878 2503 1881 2507
rect 1886 2503 1888 2507
rect 1870 2332 1873 2338
rect 1886 2332 1889 2458
rect 1902 2342 1905 2348
rect 1862 2292 1865 2318
rect 1872 2303 1874 2307
rect 1878 2303 1881 2307
rect 1886 2303 1888 2307
rect 1862 2051 1865 2168
rect 1872 2103 1874 2107
rect 1878 2103 1881 2107
rect 1886 2103 1888 2107
rect 1862 2048 1870 2051
rect 1872 1903 1874 1907
rect 1878 1903 1881 1907
rect 1886 1903 1888 1907
rect 1894 1822 1897 2278
rect 1902 2112 1905 2178
rect 1902 1912 1905 1928
rect 1926 1862 1929 3648
rect 1962 3468 1966 3471
rect 1970 3248 1974 3251
rect 2014 3152 2017 3398
rect 2038 3252 2041 3298
rect 1986 3088 1990 3091
rect 1938 2728 1942 2731
rect 1950 2592 1953 3078
rect 1966 2862 1969 2868
rect 1982 2662 1985 3048
rect 2046 3022 2049 3498
rect 2058 3348 2062 3351
rect 2026 2858 2030 2861
rect 2038 2842 2041 2948
rect 2054 2792 2057 3258
rect 2070 3132 2073 3368
rect 2094 3332 2097 3388
rect 1990 2632 1993 2788
rect 2058 2728 2062 2731
rect 2066 2668 2070 2671
rect 1954 2578 1958 2581
rect 2026 2548 2030 2551
rect 1934 2348 1942 2351
rect 1934 2282 1937 2348
rect 1934 2072 1937 2278
rect 1934 1932 1937 2068
rect 1942 1842 1945 2268
rect 1862 1712 1865 1758
rect 1894 1712 1897 1778
rect 1872 1703 1874 1707
rect 1878 1703 1881 1707
rect 1886 1703 1888 1707
rect 1902 1642 1905 1658
rect 1758 602 1761 858
rect 1782 752 1785 1268
rect 1798 1262 1801 1268
rect 1790 832 1793 1258
rect 1798 962 1801 1118
rect 1806 1072 1809 1368
rect 1814 1242 1817 1338
rect 1822 1272 1825 1328
rect 1846 1312 1849 1598
rect 1862 1502 1865 1528
rect 1872 1503 1874 1507
rect 1878 1503 1881 1507
rect 1886 1503 1888 1507
rect 1842 1268 1846 1271
rect 1846 1132 1849 1158
rect 1798 882 1801 928
rect 1790 112 1793 188
rect 1798 142 1801 148
rect 1806 12 1809 858
rect 1846 722 1849 1128
rect 1862 772 1865 1468
rect 1894 1382 1897 1528
rect 1902 1442 1905 1458
rect 1902 1382 1905 1428
rect 1874 1338 1878 1341
rect 1872 1303 1874 1307
rect 1878 1303 1881 1307
rect 1886 1303 1888 1307
rect 1882 1268 1886 1271
rect 1872 1103 1874 1107
rect 1878 1103 1881 1107
rect 1886 1103 1888 1107
rect 1872 903 1874 907
rect 1878 903 1881 907
rect 1886 903 1888 907
rect 1902 842 1905 1378
rect 1910 1282 1913 1698
rect 1918 1572 1921 1668
rect 1926 1542 1929 1718
rect 1942 1622 1945 1838
rect 1950 1692 1953 2468
rect 1958 1622 1961 2178
rect 1966 1692 1969 2458
rect 1994 2358 2001 2361
rect 1974 1611 1977 2258
rect 1966 1608 1977 1611
rect 1926 1492 1929 1498
rect 1926 1448 1934 1451
rect 1918 1262 1921 1418
rect 1926 1322 1929 1448
rect 1934 1092 1937 1138
rect 1910 862 1913 1088
rect 1930 878 1934 881
rect 1862 672 1865 708
rect 1872 703 1874 707
rect 1878 703 1881 707
rect 1886 703 1888 707
rect 1826 668 1830 671
rect 1872 503 1874 507
rect 1878 503 1881 507
rect 1886 503 1888 507
rect 1898 348 1902 351
rect 1872 303 1874 307
rect 1878 303 1881 307
rect 1886 303 1888 307
rect 1866 128 1870 131
rect 1872 103 1874 107
rect 1878 103 1881 107
rect 1886 103 1888 107
rect 1894 72 1897 98
rect 1918 71 1921 718
rect 1926 622 1929 778
rect 1942 632 1945 1428
rect 1950 812 1953 1528
rect 1958 1432 1961 1558
rect 1966 922 1969 1608
rect 1982 1582 1985 1948
rect 1990 1762 1993 2168
rect 1998 2122 2001 2358
rect 1998 1872 2001 1948
rect 2006 1922 2009 1938
rect 2014 1842 2017 2448
rect 2042 2328 2046 2331
rect 2006 1658 2014 1661
rect 1990 1538 1998 1541
rect 1982 1482 1985 1538
rect 1990 1532 1993 1538
rect 1998 1492 2001 1538
rect 2006 1522 2009 1658
rect 2022 1492 2025 1958
rect 2030 1662 2033 2328
rect 2038 1661 2041 2318
rect 2054 2162 2057 2288
rect 2070 2201 2073 2458
rect 2118 2402 2121 2448
rect 2126 2422 2129 2738
rect 2134 2501 2137 2728
rect 2142 2592 2145 3248
rect 2134 2498 2142 2501
rect 2094 2252 2097 2268
rect 2070 2198 2078 2201
rect 2078 2152 2081 2188
rect 2046 1722 2049 2108
rect 2062 1702 2065 2048
rect 2046 1672 2049 1688
rect 2062 1681 2065 1688
rect 2058 1678 2065 1681
rect 2038 1658 2049 1661
rect 2014 1482 2017 1488
rect 2030 1472 2033 1598
rect 2002 1468 2006 1471
rect 1974 1222 1977 1318
rect 1982 1142 1985 1278
rect 1974 1072 1977 1078
rect 1974 222 1977 1058
rect 1982 992 1985 1138
rect 1990 1112 1993 1128
rect 1998 1112 2001 1438
rect 1990 862 1993 1108
rect 1998 492 2001 1068
rect 2006 612 2009 1458
rect 2030 1222 2033 1468
rect 2038 1342 2041 1518
rect 2046 1452 2049 1658
rect 2062 1542 2065 1548
rect 2058 1528 2062 1531
rect 2030 1132 2033 1188
rect 2030 952 2033 968
rect 2014 412 2017 468
rect 2014 222 2017 408
rect 1994 188 1998 191
rect 1914 68 1921 71
rect 2022 62 2025 478
rect 2030 12 2033 948
rect 2038 831 2041 1158
rect 2054 832 2057 918
rect 2062 902 2065 1418
rect 2038 828 2046 831
rect 2038 622 2041 658
rect 2038 352 2041 568
rect 2038 42 2041 348
rect 2046 32 2049 688
rect 2062 21 2065 768
rect 2070 452 2073 2058
rect 2078 1782 2081 2148
rect 2086 1972 2089 2198
rect 2126 2152 2129 2238
rect 2134 2212 2137 2488
rect 2142 2462 2145 2468
rect 2150 2412 2153 2528
rect 2142 2212 2145 2408
rect 2142 2142 2145 2188
rect 2086 1942 2089 1948
rect 2078 1562 2081 1668
rect 2078 1542 2081 1558
rect 2094 1542 2097 2068
rect 2102 1942 2105 1948
rect 2110 1822 2113 2018
rect 2118 1802 2121 2068
rect 2126 1842 2129 2128
rect 2142 2012 2145 2128
rect 2158 2022 2161 2538
rect 2174 2292 2177 3698
rect 2270 3672 2273 3688
rect 2302 3532 2305 3638
rect 2346 3528 2353 3531
rect 2226 3468 2230 3471
rect 2190 3462 2193 3468
rect 2226 3448 2230 3451
rect 2182 3252 2185 3288
rect 2282 3248 2286 3251
rect 2182 2502 2185 2748
rect 2134 1952 2137 1958
rect 2090 1528 2094 1531
rect 2086 1172 2089 1458
rect 2102 1342 2105 1678
rect 2110 1332 2113 1738
rect 2118 1361 2121 1798
rect 2142 1732 2145 1858
rect 2118 1358 2126 1361
rect 2134 1322 2137 1448
rect 2142 1412 2145 1728
rect 2150 1352 2153 1508
rect 2134 1262 2137 1318
rect 2142 1182 2145 1258
rect 2086 922 2089 998
rect 2078 902 2081 908
rect 2086 722 2089 918
rect 2094 572 2097 928
rect 2102 552 2105 1128
rect 2142 852 2145 878
rect 2118 601 2121 688
rect 2114 598 2121 601
rect 2074 348 2078 351
rect 2094 212 2097 498
rect 2094 82 2097 108
rect 2062 18 2070 21
rect 2102 12 2105 548
rect 2150 262 2153 1278
rect 2158 852 2161 1908
rect 2166 1022 2169 2088
rect 2174 1882 2177 2068
rect 2182 2052 2185 2408
rect 2190 2402 2193 3148
rect 2238 2502 2241 3108
rect 2246 2862 2249 2868
rect 2302 2692 2305 3528
rect 2350 3502 2353 3528
rect 2322 3468 2326 3471
rect 2310 3462 2313 3468
rect 2358 3362 2361 3668
rect 2518 3662 2521 3668
rect 2392 3603 2394 3607
rect 2398 3603 2401 3607
rect 2406 3603 2408 3607
rect 2392 3403 2394 3407
rect 2398 3403 2401 3407
rect 2406 3403 2408 3407
rect 2310 3092 2313 3108
rect 2342 2911 2345 3228
rect 2392 3203 2394 3207
rect 2398 3203 2401 3207
rect 2406 3203 2408 3207
rect 2414 3082 2417 3508
rect 2342 2908 2350 2911
rect 2262 2672 2265 2678
rect 2366 2662 2369 3058
rect 2262 2582 2265 2658
rect 2294 2552 2297 2558
rect 2190 2232 2193 2328
rect 2182 1902 2185 2048
rect 2190 1632 2193 2228
rect 2198 1692 2201 2338
rect 2214 2322 2217 2348
rect 2174 1452 2177 1538
rect 2174 1272 2177 1278
rect 2174 1252 2177 1258
rect 2182 1082 2185 1538
rect 2190 1502 2193 1568
rect 2190 1482 2193 1488
rect 2198 1472 2201 1498
rect 2206 1362 2209 2068
rect 2214 1422 2217 2308
rect 2222 2202 2225 2248
rect 2222 1938 2230 1941
rect 2222 1902 2225 1938
rect 2222 1772 2225 1888
rect 2222 1401 2225 1768
rect 2230 1742 2233 1768
rect 2246 1672 2249 2348
rect 2254 2262 2257 2538
rect 2282 2268 2289 2271
rect 2286 2262 2289 2268
rect 2294 2262 2297 2268
rect 2214 1398 2225 1401
rect 2190 1312 2193 1358
rect 2130 128 2134 131
rect 2150 22 2153 258
rect 2158 62 2161 338
rect 2174 202 2177 938
rect 2214 712 2217 1398
rect 2222 1232 2225 1358
rect 2234 1338 2238 1341
rect 2230 1012 2233 1328
rect 2170 128 2174 131
rect 2182 32 2185 488
rect 2190 12 2193 498
rect 2198 22 2201 568
rect 2222 282 2225 368
rect 2206 132 2209 148
rect 2230 72 2233 488
rect 2246 282 2249 1478
rect 2254 1122 2257 1348
rect 2254 62 2257 548
rect 2262 272 2265 2128
rect 2294 2072 2297 2118
rect 2278 1872 2281 1978
rect 2286 1932 2289 1938
rect 2302 1892 2305 2548
rect 2314 2448 2318 2451
rect 2374 2402 2377 3028
rect 2392 3003 2394 3007
rect 2398 3003 2401 3007
rect 2406 3003 2408 3007
rect 2392 2803 2394 2807
rect 2398 2803 2401 2807
rect 2406 2803 2408 2807
rect 2382 2382 2385 2668
rect 2406 2622 2409 2648
rect 2392 2603 2394 2607
rect 2398 2603 2401 2607
rect 2406 2603 2408 2607
rect 2392 2403 2394 2407
rect 2398 2403 2401 2407
rect 2406 2403 2408 2407
rect 2318 1932 2321 2238
rect 2274 1728 2278 1731
rect 2286 1552 2289 1868
rect 2298 1838 2305 1841
rect 2302 1572 2305 1838
rect 2278 1472 2281 1548
rect 2274 1348 2278 1351
rect 2278 822 2281 1258
rect 2286 912 2289 1438
rect 2310 1252 2313 1428
rect 2294 1072 2297 1158
rect 2302 182 2305 1138
rect 2318 62 2321 1538
rect 2326 462 2329 2128
rect 2350 1852 2353 2338
rect 2358 2222 2361 2268
rect 2366 1902 2369 2278
rect 2392 2203 2394 2207
rect 2398 2203 2401 2207
rect 2406 2203 2408 2207
rect 2392 2003 2394 2007
rect 2398 2003 2401 2007
rect 2406 2003 2408 2007
rect 2386 1918 2390 1921
rect 2430 1892 2433 2248
rect 2392 1803 2394 1807
rect 2398 1803 2401 1807
rect 2406 1803 2408 1807
rect 2350 1732 2353 1748
rect 2392 1603 2394 1607
rect 2398 1603 2401 1607
rect 2406 1603 2408 1607
rect 2366 1322 2369 1538
rect 2392 1403 2394 1407
rect 2398 1403 2401 1407
rect 2406 1403 2408 1407
rect 2386 1328 2390 1331
rect 2374 1292 2377 1328
rect 2382 1282 2385 1318
rect 2334 952 2337 1258
rect 2392 1203 2394 1207
rect 2398 1203 2401 1207
rect 2406 1203 2408 1207
rect 2382 1012 2385 1078
rect 2392 1003 2394 1007
rect 2398 1003 2401 1007
rect 2406 1003 2408 1007
rect 2334 472 2337 938
rect 2342 862 2345 948
rect 2354 868 2358 871
rect 2386 858 2390 861
rect 2392 803 2394 807
rect 2398 803 2401 807
rect 2406 803 2408 807
rect 2370 738 2374 741
rect 2392 603 2394 607
rect 2398 603 2401 607
rect 2406 603 2408 607
rect 2354 468 2358 471
rect 2254 12 2257 58
rect 1734 8 1742 11
rect 2358 11 2361 278
rect 2382 262 2385 498
rect 2414 472 2417 1498
rect 2422 1342 2425 1878
rect 2434 1768 2441 1771
rect 2438 1702 2441 1768
rect 2446 1592 2449 2648
rect 2462 2592 2465 3658
rect 2670 3562 2673 3608
rect 2486 3331 2489 3418
rect 2482 3328 2489 3331
rect 2518 2811 2521 3258
rect 2550 3112 2553 3188
rect 2558 2892 2561 3128
rect 2562 2868 2566 2871
rect 2582 2862 2585 2938
rect 2514 2808 2521 2811
rect 2598 2802 2601 3378
rect 2606 3342 2609 3358
rect 2470 2762 2473 2778
rect 2582 2678 2590 2681
rect 2582 2632 2585 2678
rect 2482 2538 2486 2541
rect 2478 1962 2481 2038
rect 2454 1702 2457 1788
rect 2470 1732 2473 1738
rect 2462 1312 2465 1458
rect 2470 1282 2473 1288
rect 2446 802 2449 988
rect 2466 858 2470 861
rect 2458 738 2462 741
rect 2466 728 2470 731
rect 2426 708 2430 711
rect 2392 403 2394 407
rect 2398 403 2401 407
rect 2406 403 2408 407
rect 2398 332 2401 338
rect 2392 203 2394 207
rect 2398 203 2401 207
rect 2406 203 2408 207
rect 2382 122 2385 138
rect 2354 8 2361 11
rect 2414 12 2417 468
rect 2478 362 2481 1708
rect 2486 1482 2489 2148
rect 2494 1792 2497 2538
rect 2506 2438 2510 2441
rect 2606 2392 2609 3018
rect 2638 2742 2641 2898
rect 2654 2722 2657 3378
rect 2638 2522 2641 2588
rect 2622 2442 2625 2448
rect 2506 2348 2510 2351
rect 2510 1851 2513 2048
rect 2506 1848 2513 1851
rect 2498 1728 2502 1731
rect 2506 1678 2510 1681
rect 2510 1652 2513 1678
rect 2470 328 2478 331
rect 2470 322 2473 328
rect 2494 232 2497 1528
rect 2506 958 2510 961
rect 2518 762 2521 2128
rect 2618 2048 2622 2051
rect 2618 2038 2625 2041
rect 2526 1762 2529 1998
rect 2526 1342 2529 1358
rect 2534 952 2537 1418
rect 2550 1342 2553 1938
rect 2558 1772 2561 2008
rect 2622 1922 2625 2038
rect 2614 1732 2617 1748
rect 2542 972 2545 1328
rect 2558 1262 2561 1668
rect 2566 1562 2569 1628
rect 2586 1318 2590 1321
rect 2562 1258 2566 1261
rect 2598 882 2601 1038
rect 2606 951 2609 1498
rect 2622 1362 2625 1888
rect 2622 952 2625 958
rect 2606 948 2614 951
rect 2618 908 2622 911
rect 2586 868 2590 871
rect 2502 728 2510 731
rect 2502 722 2505 728
rect 2574 632 2577 708
rect 2614 698 2622 701
rect 2614 692 2617 698
rect 2446 72 2449 168
rect 2478 142 2481 148
rect 2526 101 2529 458
rect 2534 132 2537 138
rect 2522 98 2529 101
rect 2498 68 2502 71
rect 2446 62 2449 68
rect 2558 22 2561 448
rect 2630 422 2633 2138
rect 2638 1912 2641 2268
rect 2646 2142 2649 2158
rect 2646 1942 2649 2108
rect 2638 1832 2641 1908
rect 2646 1752 2649 1838
rect 2654 1762 2657 2678
rect 2662 2592 2665 3068
rect 2670 2842 2673 2848
rect 2678 2732 2681 2868
rect 2678 2451 2681 2478
rect 2674 2448 2681 2451
rect 2694 2362 2697 3698
rect 2702 3112 2705 3198
rect 2702 2492 2705 2658
rect 2710 2252 2713 3688
rect 2894 3452 2897 3508
rect 2904 3503 2906 3507
rect 2910 3503 2913 3507
rect 2918 3503 2920 3507
rect 2718 3212 2721 3428
rect 2726 3282 2729 3408
rect 2982 3392 2985 3468
rect 2990 3462 2993 3488
rect 2838 3242 2841 3348
rect 2890 3338 2894 3341
rect 2904 3303 2906 3307
rect 2910 3303 2913 3307
rect 2918 3303 2920 3307
rect 2822 3142 2825 3198
rect 2718 2742 2721 3118
rect 2904 3103 2906 3107
rect 2910 3103 2913 3107
rect 2918 3103 2920 3107
rect 2904 2903 2906 2907
rect 2910 2903 2913 2907
rect 2918 2903 2920 2907
rect 2826 2838 2830 2841
rect 2926 2802 2929 3108
rect 2982 3072 2985 3078
rect 2874 2548 2878 2551
rect 2774 2142 2777 2538
rect 2790 2532 2793 2548
rect 2790 2052 2793 2528
rect 2798 2132 2801 2248
rect 2806 2142 2809 2258
rect 2778 2048 2782 2051
rect 2778 1948 2785 1951
rect 2782 1912 2785 1948
rect 2798 1922 2801 2128
rect 2638 972 2641 1678
rect 2646 1592 2649 1748
rect 2674 1548 2678 1551
rect 2702 1542 2705 1898
rect 2766 1872 2769 1878
rect 2750 1642 2753 1648
rect 2782 1512 2785 1908
rect 2806 1722 2809 2138
rect 2814 2052 2817 2538
rect 2830 2352 2833 2398
rect 2830 2152 2833 2348
rect 2846 2292 2849 2418
rect 2822 2072 2825 2148
rect 2822 2062 2825 2068
rect 2830 1842 2833 2068
rect 2854 2052 2857 2238
rect 2854 1832 2857 1938
rect 2870 1712 2873 2088
rect 2810 1658 2817 1661
rect 2666 1058 2670 1061
rect 2638 872 2641 878
rect 2662 632 2665 728
rect 2674 688 2678 691
rect 2678 432 2681 458
rect 2694 392 2697 1468
rect 2742 1462 2745 1478
rect 2742 1452 2745 1458
rect 2774 1052 2777 1058
rect 2782 952 2785 1458
rect 2790 1242 2793 1268
rect 2706 938 2710 941
rect 2754 928 2761 931
rect 2758 622 2761 928
rect 2814 882 2817 1658
rect 2790 692 2793 748
rect 2814 712 2817 718
rect 2806 652 2809 708
rect 2798 532 2801 578
rect 2766 482 2769 498
rect 2758 382 2761 478
rect 2798 432 2801 528
rect 2854 372 2857 1618
rect 2862 1052 2865 1128
rect 2870 912 2873 1198
rect 2878 522 2881 1748
rect 2886 1152 2889 2348
rect 2894 2312 2897 2728
rect 2904 2703 2906 2707
rect 2910 2703 2913 2707
rect 2918 2703 2920 2707
rect 2970 2658 2974 2661
rect 3014 2602 3017 3148
rect 3026 3068 3030 3071
rect 3022 2812 3025 2848
rect 3030 2732 3033 2998
rect 2904 2503 2906 2507
rect 2910 2503 2913 2507
rect 2918 2503 2920 2507
rect 3038 2502 3041 3288
rect 3046 2962 3049 3008
rect 3054 2692 3057 3138
rect 3062 2762 3065 3328
rect 3070 3272 3073 3288
rect 3086 3242 3089 3298
rect 3094 3151 3097 3518
rect 3090 3148 3097 3151
rect 3126 3081 3129 3578
rect 3186 3348 3193 3351
rect 3190 3252 3193 3348
rect 3122 3078 3129 3081
rect 3198 3042 3201 3168
rect 3210 3058 3214 3061
rect 3126 2772 3129 2958
rect 3138 2858 3142 2861
rect 3198 2852 3201 2938
rect 3210 2778 3214 2781
rect 3222 2702 3225 2958
rect 3234 2928 3238 2931
rect 3198 2552 3201 2558
rect 3246 2512 3249 3088
rect 3258 2858 3262 2861
rect 3286 2492 3289 3688
rect 3366 3312 3369 3658
rect 3416 3603 3418 3607
rect 3422 3603 3425 3607
rect 3430 3603 3432 3607
rect 3538 3408 3545 3411
rect 3416 3403 3418 3407
rect 3422 3403 3425 3407
rect 3430 3403 3432 3407
rect 3542 3302 3545 3408
rect 3630 3402 3633 3548
rect 3928 3503 3930 3507
rect 3934 3503 3937 3507
rect 3942 3503 3944 3507
rect 3354 3298 3361 3301
rect 3342 2742 3345 3178
rect 3358 3102 3361 3298
rect 3366 2992 3369 3138
rect 3382 2922 3385 3018
rect 3382 2682 3385 2848
rect 3390 2752 3393 3108
rect 3398 3012 3401 3258
rect 3416 3203 3418 3207
rect 3422 3203 3425 3207
rect 3430 3203 3432 3207
rect 3406 3002 3409 3148
rect 3416 3003 3418 3007
rect 3422 3003 3425 3007
rect 3430 3003 3432 3007
rect 3406 2762 3409 2958
rect 3430 2942 3433 2948
rect 3438 2932 3441 2948
rect 3416 2803 3418 2807
rect 3422 2803 3425 2807
rect 3430 2803 3432 2807
rect 3390 2742 3393 2748
rect 3446 2692 3449 3068
rect 3462 2922 3465 2928
rect 3470 2692 3473 2938
rect 3486 2742 3489 2988
rect 3578 2958 3582 2961
rect 3582 2882 3585 2958
rect 3614 2822 3617 3028
rect 3558 2722 3561 2738
rect 3598 2732 3601 2758
rect 3526 2652 3529 2658
rect 2986 2438 2993 2441
rect 2990 2432 2993 2438
rect 3138 2358 3142 2361
rect 2904 2303 2906 2307
rect 2910 2303 2913 2307
rect 2918 2303 2920 2307
rect 2904 2103 2906 2107
rect 2910 2103 2913 2107
rect 2918 2103 2920 2107
rect 2934 1932 2937 2138
rect 2974 2062 2977 2208
rect 2946 2018 2950 2021
rect 2934 1922 2937 1928
rect 2942 1922 2945 1928
rect 2904 1903 2906 1907
rect 2910 1903 2913 1907
rect 2918 1903 2920 1907
rect 2926 1882 2929 1908
rect 2894 462 2897 1738
rect 2904 1703 2906 1707
rect 2910 1703 2913 1707
rect 2918 1703 2920 1707
rect 2904 1503 2906 1507
rect 2910 1503 2913 1507
rect 2918 1503 2920 1507
rect 2904 1303 2906 1307
rect 2910 1303 2913 1307
rect 2918 1303 2920 1307
rect 2902 1242 2905 1258
rect 2904 1103 2906 1107
rect 2910 1103 2913 1107
rect 2918 1103 2920 1107
rect 2904 903 2906 907
rect 2910 903 2913 907
rect 2918 903 2920 907
rect 2926 832 2929 1738
rect 2934 1682 2937 1708
rect 2942 1032 2945 1758
rect 2958 1392 2961 1458
rect 2970 1388 2974 1391
rect 2958 1212 2961 1388
rect 2904 703 2906 707
rect 2910 703 2913 707
rect 2918 703 2920 707
rect 2904 503 2906 507
rect 2910 503 2913 507
rect 2918 503 2920 507
rect 2904 303 2906 307
rect 2910 303 2913 307
rect 2918 303 2920 307
rect 2762 278 2766 281
rect 2622 222 2625 238
rect 2850 158 2854 161
rect 2734 142 2737 158
rect 2858 138 2862 141
rect 2830 82 2833 128
rect 2904 103 2906 107
rect 2910 103 2913 107
rect 2918 103 2920 107
rect 2786 78 2790 81
rect 2750 42 2753 78
rect 2814 72 2817 78
rect 2926 22 2929 798
rect 2934 602 2937 628
rect 2942 602 2945 678
rect 2950 542 2953 648
rect 2966 642 2969 1188
rect 2982 1052 2985 2138
rect 2990 1692 2993 2158
rect 3034 2148 3038 2151
rect 3062 2062 3065 2088
rect 3002 1948 3006 1951
rect 2998 1362 3001 1928
rect 3014 1672 3017 1838
rect 3022 1552 3025 1948
rect 3078 1892 3081 2298
rect 3142 2152 3145 2258
rect 3106 2138 3110 2141
rect 3086 1922 3089 1938
rect 3078 1862 3081 1888
rect 3174 1882 3177 2218
rect 3222 2052 3225 2068
rect 3186 2038 3190 2041
rect 3218 2038 3222 2041
rect 3246 2012 3249 2468
rect 3326 2432 3329 2628
rect 3416 2603 3418 2607
rect 3422 2603 3425 2607
rect 3430 2603 3432 2607
rect 3590 2592 3593 2688
rect 3614 2672 3617 2818
rect 3622 2752 3625 2958
rect 3538 2548 3542 2551
rect 3638 2542 3641 2548
rect 3342 2392 3345 2508
rect 3534 2452 3537 2468
rect 3416 2403 3418 2407
rect 3422 2403 3425 2407
rect 3430 2403 3432 2407
rect 3342 2362 3345 2388
rect 3266 2358 3270 2361
rect 3534 2292 3537 2448
rect 3586 2268 3590 2271
rect 3416 2203 3418 2207
rect 3422 2203 3425 2207
rect 3430 2203 3432 2207
rect 3322 2148 3326 2151
rect 3270 2142 3273 2148
rect 3406 2072 3409 2078
rect 3294 1902 3297 2058
rect 3416 2003 3418 2007
rect 3422 2003 3425 2007
rect 3430 2003 3432 2007
rect 3438 2002 3441 2168
rect 3346 1938 3350 1941
rect 3034 1538 3038 1541
rect 2998 1342 3001 1358
rect 3078 1262 3081 1268
rect 3002 1258 3006 1261
rect 3094 1202 3097 1738
rect 3110 1002 3113 1848
rect 3158 1422 3161 1848
rect 3186 1558 3193 1561
rect 3190 1522 3193 1558
rect 3290 1478 3294 1481
rect 3310 1392 3313 1918
rect 3326 1442 3329 1848
rect 3334 1532 3337 1748
rect 3382 1542 3385 1548
rect 3206 1352 3209 1378
rect 3374 1322 3377 1428
rect 3306 1268 3310 1271
rect 3390 1212 3393 1978
rect 3406 1772 3409 1808
rect 3416 1803 3418 1807
rect 3422 1803 3425 1807
rect 3430 1803 3432 1807
rect 3462 1762 3465 2118
rect 3490 2068 3494 2071
rect 3474 1658 3478 1661
rect 3416 1603 3418 1607
rect 3422 1603 3425 1607
rect 3430 1603 3432 1607
rect 3502 1522 3505 2258
rect 3510 1952 3513 2108
rect 3534 1942 3537 2178
rect 3598 2162 3601 2318
rect 3678 2312 3681 2558
rect 3574 1972 3577 2158
rect 3598 2152 3601 2158
rect 3630 2072 3633 2198
rect 3522 1548 3526 1551
rect 3502 1442 3505 1518
rect 3510 1482 3513 1488
rect 3416 1403 3418 1407
rect 3422 1403 3425 1407
rect 3430 1403 3432 1407
rect 3402 1258 3409 1261
rect 3406 1112 3409 1258
rect 3416 1203 3418 1207
rect 3422 1203 3425 1207
rect 3430 1203 3432 1207
rect 3462 1132 3465 1428
rect 3534 1362 3537 1938
rect 3582 1922 3585 1938
rect 3694 1932 3697 2658
rect 3710 2591 3713 3448
rect 3774 3438 3782 3441
rect 3718 2942 3721 2948
rect 3726 2722 3729 3138
rect 3734 2902 3737 2938
rect 3750 2792 3753 2798
rect 3706 2588 3713 2591
rect 3590 1922 3593 1928
rect 3702 1862 3705 2528
rect 3750 2522 3753 2748
rect 3714 2088 3718 2091
rect 3710 1772 3713 1918
rect 3522 1348 3526 1351
rect 3542 1342 3545 1348
rect 3494 1252 3497 1328
rect 3498 1248 3505 1251
rect 3502 1122 3505 1248
rect 3038 881 3041 888
rect 3026 878 3041 881
rect 3118 872 3121 878
rect 3054 742 3057 758
rect 3102 742 3105 748
rect 3166 682 3169 688
rect 3214 672 3217 1068
rect 3416 1003 3418 1007
rect 3422 1003 3425 1007
rect 3430 1003 3432 1007
rect 3326 862 3329 898
rect 3470 862 3473 948
rect 3482 868 3486 871
rect 3326 732 3329 858
rect 3416 803 3418 807
rect 3422 803 3425 807
rect 3430 803 3432 807
rect 3254 722 3257 728
rect 2934 362 2937 498
rect 3214 472 3217 668
rect 3326 662 3329 728
rect 3416 603 3418 607
rect 3422 603 3425 607
rect 3430 603 3432 607
rect 3346 598 3353 601
rect 3350 482 3353 598
rect 3246 458 3254 461
rect 2954 158 2958 161
rect 2942 72 2945 78
rect 2974 12 2977 388
rect 2986 138 2990 141
rect 3006 11 3009 458
rect 3078 242 3081 258
rect 3082 128 3086 131
rect 3070 91 3073 128
rect 3066 88 3073 91
rect 3094 12 3097 348
rect 3106 338 3110 341
rect 3102 172 3105 338
rect 3170 238 3174 241
rect 3150 152 3153 168
rect 3150 42 3153 68
rect 3182 22 3185 368
rect 3246 292 3249 458
rect 3438 422 3441 538
rect 3470 452 3473 538
rect 3416 403 3418 407
rect 3422 403 3425 407
rect 3430 403 3432 407
rect 3294 282 3297 338
rect 3290 278 3294 281
rect 3234 258 3238 261
rect 3270 102 3273 118
rect 3254 98 3262 101
rect 3254 62 3257 98
rect 3334 12 3337 358
rect 3366 332 3369 388
rect 3438 352 3441 418
rect 3342 71 3345 128
rect 3350 112 3353 128
rect 3350 82 3353 88
rect 3358 72 3361 78
rect 3366 72 3369 328
rect 3478 302 3481 318
rect 3374 252 3377 258
rect 3470 252 3473 298
rect 3416 203 3418 207
rect 3422 203 3425 207
rect 3430 203 3432 207
rect 3438 202 3441 218
rect 3394 128 3398 131
rect 3342 68 3350 71
rect 3414 62 3417 68
rect 3510 12 3513 748
rect 3522 738 3526 741
rect 3550 682 3553 1748
rect 3562 1658 3566 1661
rect 3558 1638 3566 1641
rect 3558 1302 3561 1638
rect 3678 1608 3686 1611
rect 3678 1342 3681 1608
rect 3694 1572 3697 1608
rect 3726 1522 3729 1538
rect 3702 1222 3705 1448
rect 3734 1072 3737 1118
rect 3742 822 3745 1938
rect 3766 882 3769 3348
rect 3774 3132 3777 3438
rect 3846 3292 3849 3358
rect 3928 3303 3930 3307
rect 3934 3303 3937 3307
rect 3942 3303 3944 3307
rect 3950 3192 3953 3398
rect 3846 3062 3849 3068
rect 3870 3062 3873 3148
rect 3928 3103 3930 3107
rect 3934 3103 3937 3107
rect 3942 3103 3944 3107
rect 3910 3072 3913 3098
rect 3974 3051 3977 3698
rect 3974 3048 3982 3051
rect 3928 2903 3930 2907
rect 3934 2903 3937 2907
rect 3942 2903 3944 2907
rect 3874 2748 3878 2751
rect 3962 2748 3966 2751
rect 3890 2738 3894 2741
rect 3928 2703 3930 2707
rect 3934 2703 3937 2707
rect 3942 2703 3944 2707
rect 3950 2512 3953 2528
rect 3928 2503 3930 2507
rect 3934 2503 3937 2507
rect 3942 2503 3944 2507
rect 3774 2292 3777 2308
rect 3928 2303 3930 2307
rect 3934 2303 3937 2307
rect 3942 2303 3944 2307
rect 3910 2132 3913 2148
rect 3826 2128 3830 2131
rect 3928 2103 3930 2107
rect 3934 2103 3937 2107
rect 3942 2103 3944 2107
rect 3870 1892 3873 1948
rect 3818 1688 3822 1691
rect 3894 1482 3897 1968
rect 3928 1903 3930 1907
rect 3934 1903 3937 1907
rect 3942 1903 3944 1907
rect 3928 1703 3930 1707
rect 3934 1703 3937 1707
rect 3942 1703 3944 1707
rect 3928 1503 3930 1507
rect 3934 1503 3937 1507
rect 3942 1503 3944 1507
rect 3790 1442 3793 1448
rect 3918 1282 3921 1468
rect 3928 1303 3930 1307
rect 3934 1303 3937 1307
rect 3942 1303 3944 1307
rect 3950 1292 3953 1658
rect 3958 1462 3961 1708
rect 3966 1182 3969 1698
rect 3974 1552 3977 3048
rect 3998 2632 4001 3698
rect 4078 3622 4081 3698
rect 4086 3482 4089 3648
rect 4110 3361 4113 3548
rect 4106 3358 4113 3361
rect 4110 3032 4113 3258
rect 4214 2922 4217 3698
rect 4238 3552 4241 3688
rect 4270 3132 4273 3258
rect 4278 3052 4281 3348
rect 4022 2558 4030 2561
rect 4022 2502 4025 2558
rect 3982 2372 3985 2468
rect 4014 2252 4017 2408
rect 4038 2212 4041 2308
rect 4054 2072 4057 2328
rect 3982 2062 3985 2068
rect 4054 1822 4057 2068
rect 4070 1972 4073 2828
rect 4294 2752 4297 3688
rect 4302 3172 4305 3538
rect 4366 3462 4369 3468
rect 4334 3452 4337 3458
rect 4374 2862 4377 3698
rect 5238 3698 5246 3701
rect 4440 3603 4442 3607
rect 4446 3603 4449 3607
rect 4454 3603 4456 3607
rect 4482 3478 4486 3481
rect 4494 3462 4497 3548
rect 4570 3478 4574 3481
rect 4610 3468 4614 3471
rect 4386 3458 4390 3461
rect 4440 3403 4442 3407
rect 4446 3403 4449 3407
rect 4454 3403 4456 3407
rect 4650 3398 4657 3401
rect 4554 3318 4561 3321
rect 4558 3232 4561 3318
rect 4440 3203 4442 3207
rect 4446 3203 4449 3207
rect 4454 3203 4456 3207
rect 4654 3092 4657 3398
rect 4670 3292 4673 3458
rect 4718 3438 4726 3441
rect 4682 3358 4686 3361
rect 4718 3272 4721 3438
rect 4734 3242 4737 3348
rect 4742 3262 4745 3518
rect 4886 3462 4889 3528
rect 4952 3503 4954 3507
rect 4958 3503 4961 3507
rect 4966 3503 4968 3507
rect 4886 3342 4889 3458
rect 5014 3392 5017 3478
rect 5002 3358 5009 3361
rect 5006 3342 5009 3358
rect 5014 3352 5017 3388
rect 5022 3352 5025 3358
rect 4870 3182 4873 3288
rect 4890 3278 4894 3281
rect 4910 3192 4913 3338
rect 4952 3303 4954 3307
rect 4958 3303 4961 3307
rect 4966 3303 4968 3307
rect 4950 3282 4953 3288
rect 4922 3268 4926 3271
rect 4870 3161 4873 3178
rect 4870 3158 4878 3161
rect 4942 3092 4945 3278
rect 4958 3272 4961 3278
rect 4952 3103 4954 3107
rect 4958 3103 4961 3107
rect 4966 3103 4968 3107
rect 4440 3003 4442 3007
rect 4446 3003 4449 3007
rect 4454 3003 4456 3007
rect 4952 2903 4954 2907
rect 4958 2903 4961 2907
rect 4966 2903 4968 2907
rect 4882 2828 4886 2831
rect 4440 2803 4442 2807
rect 4446 2803 4449 2807
rect 4454 2803 4456 2807
rect 4294 2722 4297 2748
rect 4502 2742 4505 2748
rect 4546 2738 4550 2741
rect 4440 2603 4442 2607
rect 4446 2603 4449 2607
rect 4454 2603 4456 2607
rect 4678 2582 4681 2698
rect 4710 2561 4713 2708
rect 4734 2641 4737 2698
rect 4734 2638 4742 2641
rect 4710 2558 4718 2561
rect 4834 2548 4838 2551
rect 4110 2262 4113 2268
rect 3974 1462 3977 1498
rect 4014 1192 4017 1548
rect 4102 1172 4105 1748
rect 4126 1692 4129 2548
rect 4190 2432 4193 2498
rect 4246 2362 4249 2538
rect 4506 2468 4513 2471
rect 4322 2388 4329 2391
rect 4290 2238 4294 2241
rect 4142 1902 4145 2108
rect 4158 1872 4161 2218
rect 4242 2058 4249 2061
rect 4178 1938 4182 1941
rect 4158 1542 4161 1868
rect 4246 1812 4249 2058
rect 4302 1862 4305 1868
rect 4198 1372 4201 1458
rect 4198 1262 4201 1368
rect 4214 1292 4217 1548
rect 4254 1492 4257 1818
rect 4326 1442 4329 2388
rect 4382 2242 4385 2268
rect 4390 2232 4393 2258
rect 4342 1512 4345 2058
rect 4350 1862 4353 1868
rect 4350 1692 4353 1758
rect 4358 1752 4361 1888
rect 4366 1742 4369 1758
rect 4374 1542 4377 2078
rect 4398 2022 4401 2448
rect 4440 2403 4442 2407
rect 4446 2403 4449 2407
rect 4454 2403 4456 2407
rect 4440 2203 4442 2207
rect 4446 2203 4449 2207
rect 4454 2203 4456 2207
rect 4406 1832 4409 2058
rect 4440 2003 4442 2007
rect 4446 2003 4449 2007
rect 4454 2003 4456 2007
rect 4430 1612 4433 1988
rect 4440 1803 4442 1807
rect 4446 1803 4449 1807
rect 4454 1803 4456 1807
rect 4440 1603 4442 1607
rect 4446 1603 4449 1607
rect 4454 1603 4456 1607
rect 4478 1582 4481 2108
rect 4494 2072 4497 2088
rect 4510 2032 4513 2468
rect 4526 2112 4529 2548
rect 4734 2532 4737 2548
rect 4574 2242 4577 2258
rect 4526 1732 4529 1778
rect 4478 1552 4481 1578
rect 4542 1532 4545 1538
rect 4442 1528 4446 1531
rect 4440 1403 4442 1407
rect 4446 1403 4449 1407
rect 4454 1403 4456 1407
rect 4294 1262 4297 1348
rect 4398 1342 4401 1348
rect 4506 1278 4510 1281
rect 4270 1172 4273 1218
rect 4440 1203 4442 1207
rect 4446 1203 4449 1207
rect 4454 1203 4456 1207
rect 4102 1152 4105 1168
rect 4238 1162 4241 1168
rect 3928 1103 3930 1107
rect 3934 1103 3937 1107
rect 3942 1103 3944 1107
rect 3950 1082 3953 1098
rect 3928 903 3930 907
rect 3934 903 3937 907
rect 3942 903 3944 907
rect 3582 732 3585 738
rect 3550 462 3553 468
rect 3558 22 3561 638
rect 3618 568 3622 571
rect 3678 462 3681 468
rect 3650 458 3654 461
rect 3606 322 3609 338
rect 3590 172 3593 308
rect 3574 72 3577 78
rect 3622 72 3625 108
rect 3610 68 3614 71
rect 3650 58 3654 61
rect 3718 22 3721 788
rect 4022 742 4025 1078
rect 4238 992 4241 1158
rect 4440 1003 4442 1007
rect 4446 1003 4449 1007
rect 4454 1003 4456 1007
rect 4222 932 4225 948
rect 4390 942 4393 968
rect 4170 928 4174 931
rect 4126 812 4129 908
rect 4440 803 4442 807
rect 4446 803 4449 807
rect 4454 803 4456 807
rect 4198 752 4201 768
rect 3928 703 3930 707
rect 3934 703 3937 707
rect 3942 703 3944 707
rect 3958 662 3961 668
rect 3962 568 3966 571
rect 3762 468 3766 471
rect 3838 462 3841 528
rect 3928 503 3930 507
rect 3934 503 3937 507
rect 3942 503 3944 507
rect 3734 292 3737 328
rect 3794 278 3798 281
rect 3854 92 3857 168
rect 3918 102 3921 408
rect 3928 303 3930 307
rect 3934 303 3937 307
rect 3942 303 3944 307
rect 3928 103 3930 107
rect 3934 103 3937 107
rect 3942 103 3944 107
rect 3982 92 3985 558
rect 3998 272 4001 738
rect 4034 658 4038 661
rect 4022 302 4025 648
rect 4054 432 4057 528
rect 4078 388 4086 391
rect 4078 302 4081 388
rect 4102 192 4105 328
rect 3006 8 3014 11
rect 4046 11 4049 138
rect 4094 22 4097 158
rect 4102 102 4105 178
rect 4142 122 4145 308
rect 4174 252 4177 568
rect 4198 12 4201 748
rect 4262 692 4265 748
rect 4550 702 4553 2068
rect 4606 1742 4609 1848
rect 4582 1482 4585 1688
rect 4614 1542 4617 2508
rect 4798 2342 4801 2348
rect 4630 2282 4633 2288
rect 4682 2278 4686 2281
rect 4630 1902 4633 2028
rect 4710 1942 4713 2338
rect 4738 2278 4742 2281
rect 4722 2258 4726 2261
rect 4718 2062 4721 2068
rect 4686 1908 4694 1911
rect 4630 1352 4633 1898
rect 4638 1762 4641 1858
rect 4686 1682 4689 1908
rect 4638 1432 4641 1528
rect 4662 1252 4665 1468
rect 4702 1322 4705 1908
rect 4710 1522 4713 1938
rect 4738 1928 4745 1931
rect 4742 1322 4745 1928
rect 4750 1751 4753 1778
rect 4750 1748 4758 1751
rect 4578 1248 4585 1251
rect 4582 1102 4585 1248
rect 4738 1148 4742 1151
rect 4622 842 4625 1098
rect 4742 1062 4745 1088
rect 4262 672 4265 678
rect 4314 648 4318 651
rect 4440 603 4442 607
rect 4446 603 4449 607
rect 4454 603 4456 607
rect 4226 288 4230 291
rect 4262 92 4265 498
rect 4440 403 4442 407
rect 4446 403 4449 407
rect 4454 403 4456 407
rect 4334 282 4337 288
rect 4342 162 4345 378
rect 4440 203 4442 207
rect 4446 203 4449 207
rect 4454 203 4456 207
rect 4046 8 4054 11
rect 4422 11 4425 158
rect 4486 22 4489 688
rect 4574 672 4577 818
rect 4766 802 4769 2068
rect 4798 2052 4801 2268
rect 4798 1862 4801 2048
rect 4822 1872 4825 2388
rect 4830 2341 4833 2358
rect 4830 2338 4838 2341
rect 4790 1342 4793 1518
rect 4854 1391 4857 1548
rect 4854 1388 4862 1391
rect 4878 1222 4881 2668
rect 4894 1872 4897 2298
rect 4902 2122 4905 2738
rect 4952 2703 4954 2707
rect 4958 2703 4961 2707
rect 4966 2703 4968 2707
rect 4952 2503 4954 2507
rect 4958 2503 4961 2507
rect 4966 2503 4968 2507
rect 4910 2262 4913 2278
rect 4942 1991 4945 2328
rect 4952 2303 4954 2307
rect 4958 2303 4961 2307
rect 4966 2303 4968 2307
rect 4958 2142 4961 2198
rect 4952 2103 4954 2107
rect 4958 2103 4961 2107
rect 4966 2103 4968 2107
rect 4938 1988 4945 1991
rect 4982 2092 4985 2508
rect 5006 2252 5009 2338
rect 4952 1903 4954 1907
rect 4958 1903 4961 1907
rect 4966 1903 4968 1907
rect 4886 1122 4889 1848
rect 4902 1262 4905 1348
rect 4910 1062 4913 1868
rect 4982 1752 4985 2088
rect 5014 1872 5017 2528
rect 5022 1872 5025 2728
rect 4952 1703 4954 1707
rect 4958 1703 4961 1707
rect 4966 1703 4968 1707
rect 4918 1662 4921 1668
rect 4606 752 4609 758
rect 4674 748 4678 751
rect 4942 722 4945 1578
rect 4952 1503 4954 1507
rect 4958 1503 4961 1507
rect 4966 1503 4968 1507
rect 4974 1471 4977 1598
rect 4974 1468 4982 1471
rect 4952 1303 4954 1307
rect 4958 1303 4961 1307
rect 4966 1303 4968 1307
rect 4952 1103 4954 1107
rect 4958 1103 4961 1107
rect 4966 1103 4968 1107
rect 5006 1092 5009 1858
rect 5014 1652 5017 1868
rect 5030 1672 5033 1938
rect 5030 1352 5033 1458
rect 5022 1062 5025 1288
rect 5030 1012 5033 1348
rect 5046 1241 5049 1538
rect 5054 1252 5057 3028
rect 5102 2732 5105 2748
rect 5106 2638 5110 2641
rect 5086 2442 5089 2478
rect 5062 2152 5065 2368
rect 5082 2348 5086 2351
rect 5070 1761 5073 1768
rect 5066 1758 5073 1761
rect 5066 1268 5073 1271
rect 5042 1238 5049 1241
rect 5070 1242 5073 1268
rect 4952 903 4954 907
rect 4958 903 4961 907
rect 4966 903 4968 907
rect 5054 872 5057 1228
rect 5078 1062 5081 1618
rect 4952 703 4954 707
rect 4958 703 4961 707
rect 4966 703 4968 707
rect 5054 542 5057 868
rect 5094 762 5097 2548
rect 5126 1992 5129 2448
rect 5126 862 5129 1868
rect 5134 1482 5137 2768
rect 5142 2632 5145 2638
rect 5150 2292 5153 2658
rect 5142 682 5145 2218
rect 5150 1982 5153 2288
rect 5150 1882 5153 1978
rect 5150 1672 5153 1698
rect 5158 1361 5161 2318
rect 5166 2022 5169 2538
rect 5174 2032 5177 3658
rect 5238 3652 5241 3698
rect 5306 3648 5310 3651
rect 5182 3222 5185 3348
rect 5182 1962 5185 2218
rect 5190 1962 5193 3548
rect 5198 2412 5201 2418
rect 5206 2202 5209 3528
rect 5214 2352 5217 3338
rect 5198 2162 5201 2168
rect 5150 1358 5161 1361
rect 5166 1512 5169 1738
rect 5174 1712 5177 1848
rect 5150 772 5153 1358
rect 5158 1222 5161 1348
rect 5166 742 5169 1508
rect 5174 932 5177 1648
rect 5182 1522 5185 1948
rect 5190 1482 5193 1878
rect 5198 1782 5201 1958
rect 5206 1942 5209 2198
rect 5206 1832 5209 1938
rect 5198 1672 5201 1768
rect 5206 1542 5209 1828
rect 5214 1752 5217 2348
rect 5214 1682 5217 1748
rect 5190 672 5193 1408
rect 5206 972 5209 1538
rect 5198 952 5201 958
rect 5206 752 5209 788
rect 5214 622 5217 1678
rect 5222 1212 5225 2928
rect 5230 1661 5233 3048
rect 5238 2262 5241 2948
rect 5238 2112 5241 2248
rect 5238 2042 5241 2098
rect 5246 1981 5249 3288
rect 5254 3172 5257 3368
rect 5238 1978 5249 1981
rect 5238 1752 5241 1978
rect 5238 1692 5241 1748
rect 5246 1712 5249 1968
rect 5254 1872 5257 3158
rect 5262 2651 5265 3618
rect 5282 3548 5286 3551
rect 5270 3452 5273 3458
rect 5270 2992 5273 3438
rect 5278 3432 5281 3438
rect 5278 3072 5281 3228
rect 5270 2702 5273 2938
rect 5262 2648 5270 2651
rect 5238 1672 5241 1678
rect 5230 1658 5241 1661
rect 5230 942 5233 1298
rect 5238 1282 5241 1658
rect 5246 1292 5249 1698
rect 5246 1272 5249 1278
rect 5238 962 5241 1258
rect 5246 872 5249 878
rect 5254 692 5257 1868
rect 5254 552 5257 558
rect 4952 503 4954 507
rect 4958 503 4961 507
rect 4966 503 4968 507
rect 5070 472 5073 478
rect 4866 468 4870 471
rect 5062 462 5065 468
rect 4938 458 4942 461
rect 4614 362 4617 408
rect 5262 372 5265 2638
rect 5270 542 5273 2648
rect 5278 2512 5281 3048
rect 4952 303 4954 307
rect 4958 303 4961 307
rect 4966 303 4968 307
rect 4558 91 4561 258
rect 5206 152 5209 298
rect 4952 103 4954 107
rect 4958 103 4961 107
rect 4966 103 4968 107
rect 4554 88 4561 91
rect 4422 8 4430 11
rect 5246 11 5249 138
rect 5262 52 5265 368
rect 5270 362 5273 528
rect 5278 342 5281 2508
rect 5286 2472 5289 3258
rect 5294 3192 5297 3468
rect 5294 2672 5297 3178
rect 5302 3072 5305 3358
rect 5302 2692 5305 3058
rect 5302 2672 5305 2678
rect 5298 2658 5305 2661
rect 5302 2632 5305 2658
rect 5294 2572 5297 2628
rect 5294 2522 5297 2558
rect 5302 2542 5305 2578
rect 5286 1722 5289 2468
rect 5278 252 5281 338
rect 5286 192 5289 1718
rect 5294 72 5297 2508
rect 5302 2152 5305 2528
rect 5310 2282 5313 3558
rect 5310 2152 5313 2258
rect 5302 1522 5305 2128
rect 5310 2052 5313 2138
rect 5358 2132 5361 3568
rect 5310 1662 5313 1668
rect 5302 882 5305 1488
rect 5310 1462 5313 1488
rect 5310 1152 5313 1158
rect 5310 1082 5313 1088
rect 5310 952 5313 958
rect 5306 858 5310 861
rect 5302 152 5305 538
rect 5310 322 5313 838
rect 5302 82 5305 88
rect 5242 8 5249 11
rect 344 3 346 7
rect 350 3 353 7
rect 358 3 360 7
rect 1368 3 1370 7
rect 1374 3 1377 7
rect 1382 3 1384 7
rect 2392 3 2394 7
rect 2398 3 2401 7
rect 2406 3 2408 7
rect 3416 3 3418 7
rect 3422 3 3425 7
rect 3430 3 3432 7
rect 4440 3 4442 7
rect 4446 3 4449 7
rect 4454 3 4456 7
<< m5contact >>
rect 858 3703 862 3707
rect 865 3703 866 3707
rect 866 3703 869 3707
rect 1874 3703 1878 3707
rect 1881 3703 1882 3707
rect 1882 3703 1885 3707
rect 2906 3703 2910 3707
rect 2913 3703 2914 3707
rect 2914 3703 2917 3707
rect 3930 3703 3934 3707
rect 3937 3703 3938 3707
rect 3938 3703 3941 3707
rect 4954 3703 4958 3707
rect 4961 3703 4962 3707
rect 4962 3703 4965 3707
rect 942 3668 946 3672
rect 966 3668 970 3672
rect 1206 3668 1210 3672
rect 1358 3668 1362 3672
rect 1790 3678 1794 3682
rect 1974 3678 1978 3682
rect 346 3603 350 3607
rect 353 3603 354 3607
rect 354 3603 357 3607
rect 346 3403 350 3407
rect 353 3403 354 3407
rect 354 3403 357 3407
rect 346 3203 350 3207
rect 353 3203 354 3207
rect 354 3203 357 3207
rect 526 3368 530 3372
rect 582 3368 586 3372
rect 346 3003 350 3007
rect 353 3003 354 3007
rect 354 3003 357 3007
rect 346 2803 350 2807
rect 353 2803 354 2807
rect 354 2803 357 2807
rect 22 2608 26 2612
rect 110 2598 114 2602
rect 142 2538 146 2542
rect 346 2603 350 2607
rect 353 2603 354 2607
rect 354 2603 357 2607
rect 566 3138 570 3142
rect 638 3128 642 3132
rect 198 2538 202 2542
rect 1094 3548 1098 3552
rect 858 3503 862 3507
rect 865 3503 866 3507
rect 866 3503 869 3507
rect 814 3288 818 3292
rect 662 2738 666 2742
rect 22 2198 26 2202
rect 54 2068 58 2072
rect 102 2128 106 2132
rect 190 2288 194 2292
rect 346 2403 350 2407
rect 353 2403 354 2407
rect 354 2403 357 2407
rect 118 2208 122 2212
rect 346 2203 350 2207
rect 353 2203 354 2207
rect 354 2203 357 2207
rect 366 2118 370 2122
rect 302 2068 306 2072
rect 346 2003 350 2007
rect 353 2003 354 2007
rect 354 2003 357 2007
rect 346 1803 350 1807
rect 353 1803 354 1807
rect 354 1803 357 1807
rect 102 1558 106 1562
rect 174 1558 178 1562
rect 630 2578 634 2582
rect 662 2558 666 2562
rect 646 2368 650 2372
rect 710 2318 714 2322
rect 494 2158 498 2162
rect 838 3068 842 3072
rect 942 3338 946 3342
rect 858 3303 862 3307
rect 865 3303 866 3307
rect 866 3303 869 3307
rect 902 3298 906 3302
rect 950 3298 954 3302
rect 958 3288 962 3292
rect 902 3258 906 3262
rect 858 3103 862 3107
rect 865 3103 866 3107
rect 866 3103 869 3107
rect 1150 3548 1154 3552
rect 1022 3348 1026 3352
rect 1070 3288 1074 3292
rect 1046 3258 1050 3262
rect 862 2918 866 2922
rect 858 2903 862 2907
rect 865 2903 866 2907
rect 866 2903 869 2907
rect 858 2703 862 2707
rect 865 2703 866 2707
rect 866 2703 869 2707
rect 854 2558 858 2562
rect 858 2503 862 2507
rect 865 2503 866 2507
rect 866 2503 869 2507
rect 858 2303 862 2307
rect 865 2303 866 2307
rect 866 2303 869 2307
rect 858 2103 862 2107
rect 865 2103 866 2107
rect 866 2103 869 2107
rect 346 1603 350 1607
rect 353 1603 354 1607
rect 354 1603 357 1607
rect 534 1748 538 1752
rect 174 1478 178 1482
rect 254 1478 258 1482
rect 346 1403 350 1407
rect 353 1403 354 1407
rect 354 1403 357 1407
rect 346 1203 350 1207
rect 353 1203 354 1207
rect 354 1203 357 1207
rect 346 1003 350 1007
rect 353 1003 354 1007
rect 354 1003 357 1007
rect 858 1903 862 1907
rect 865 1903 866 1907
rect 866 1903 869 1907
rect 646 1858 650 1862
rect 902 2358 906 2362
rect 894 2018 898 2022
rect 990 2678 994 2682
rect 1054 2678 1058 2682
rect 1078 2648 1082 2652
rect 1086 2638 1090 2642
rect 1126 2638 1130 2642
rect 1030 2438 1034 2442
rect 1030 2288 1034 2292
rect 958 2238 962 2242
rect 1030 2188 1034 2192
rect 918 1768 922 1772
rect 406 1168 410 1172
rect 590 1068 594 1072
rect 6 888 10 892
rect 542 878 546 882
rect 858 1703 862 1707
rect 865 1703 866 1707
rect 866 1703 869 1707
rect 630 1658 634 1662
rect 694 1688 698 1692
rect 894 1688 898 1692
rect 686 1658 690 1662
rect 766 1658 770 1662
rect 718 1488 722 1492
rect 854 1608 858 1612
rect 814 1438 818 1442
rect 806 1258 810 1262
rect 858 1503 862 1507
rect 865 1503 866 1507
rect 866 1503 869 1507
rect 870 1458 874 1462
rect 858 1303 862 1307
rect 865 1303 866 1307
rect 866 1303 869 1307
rect 862 1258 866 1262
rect 858 1103 862 1107
rect 865 1103 866 1107
rect 866 1103 869 1107
rect 710 1068 714 1072
rect 806 948 810 952
rect 858 903 862 907
rect 865 903 866 907
rect 866 903 869 907
rect 742 888 746 892
rect 6 818 10 822
rect 346 803 350 807
rect 353 803 354 807
rect 354 803 357 807
rect 502 778 506 782
rect 190 648 194 652
rect 62 358 66 362
rect 254 658 258 662
rect 438 728 442 732
rect 334 648 338 652
rect 390 648 394 652
rect 346 603 350 607
rect 353 603 354 607
rect 354 603 357 607
rect 326 548 330 552
rect 346 403 350 407
rect 353 403 354 407
rect 354 403 357 407
rect 334 338 338 342
rect 346 203 350 207
rect 353 203 354 207
rect 354 203 357 207
rect 798 758 802 762
rect 542 728 546 732
rect 654 728 658 732
rect 558 688 562 692
rect 534 658 538 662
rect 710 528 714 532
rect 558 458 562 462
rect 486 148 490 152
rect 518 78 522 82
rect 534 138 538 142
rect 542 78 546 82
rect 534 68 538 72
rect 654 148 658 152
rect 606 138 610 142
rect 742 58 746 62
rect 858 703 862 707
rect 865 703 866 707
rect 866 703 869 707
rect 806 538 810 542
rect 858 503 862 507
rect 865 503 866 507
rect 866 503 869 507
rect 858 303 862 307
rect 865 303 866 307
rect 866 303 869 307
rect 966 1608 970 1612
rect 942 1548 946 1552
rect 934 958 938 962
rect 1070 2358 1074 2362
rect 1182 3358 1186 3362
rect 1182 3328 1186 3332
rect 1254 3358 1258 3362
rect 1270 3348 1274 3352
rect 1254 3288 1258 3292
rect 1206 3068 1210 3072
rect 1222 3048 1226 3052
rect 1318 3048 1322 3052
rect 1370 3603 1374 3607
rect 1377 3603 1378 3607
rect 1378 3603 1381 3607
rect 1370 3403 1374 3407
rect 1377 3403 1378 3407
rect 1378 3403 1381 3407
rect 1366 3338 1370 3342
rect 1350 3328 1354 3332
rect 1510 3648 1514 3652
rect 1622 3648 1626 3652
rect 1470 3348 1474 3352
rect 1462 3328 1466 3332
rect 1414 3318 1418 3322
rect 1370 3203 1374 3207
rect 1377 3203 1378 3207
rect 1378 3203 1381 3207
rect 1370 3003 1374 3007
rect 1377 3003 1378 3007
rect 1378 3003 1381 3007
rect 1542 3438 1546 3442
rect 1422 2918 1426 2922
rect 1370 2803 1374 2807
rect 1377 2803 1378 2807
rect 1378 2803 1381 2807
rect 1370 2603 1374 2607
rect 1377 2603 1378 2607
rect 1378 2603 1381 2607
rect 1370 2403 1374 2407
rect 1377 2403 1378 2407
rect 1378 2403 1381 2407
rect 1390 2368 1394 2372
rect 1102 2228 1106 2232
rect 1094 2128 1098 2132
rect 1078 2118 1082 2122
rect 998 1538 1002 1542
rect 1086 1538 1090 1542
rect 1118 1488 1122 1492
rect 1062 1358 1066 1362
rect 1118 1358 1122 1362
rect 1038 958 1042 962
rect 1046 858 1050 862
rect 1078 688 1082 692
rect 894 528 898 532
rect 1030 528 1034 532
rect 858 103 862 107
rect 865 103 866 107
rect 866 103 869 107
rect 950 68 954 72
rect 966 68 970 72
rect 1046 68 1050 72
rect 990 58 994 62
rect 1150 1858 1154 1862
rect 1142 1768 1146 1772
rect 1142 1548 1146 1552
rect 1370 2203 1374 2207
rect 1377 2203 1378 2207
rect 1378 2203 1381 2207
rect 1334 2168 1338 2172
rect 1262 2148 1266 2152
rect 1342 2058 1346 2062
rect 1246 2038 1250 2042
rect 1370 2003 1374 2007
rect 1377 2003 1378 2007
rect 1378 2003 1381 2007
rect 1286 1868 1290 1872
rect 1310 1788 1314 1792
rect 1214 1758 1218 1762
rect 1238 1748 1242 1752
rect 1198 1488 1202 1492
rect 1190 1478 1194 1482
rect 1174 1348 1178 1352
rect 1302 1468 1306 1472
rect 1334 1468 1338 1472
rect 1318 1438 1322 1442
rect 1246 1278 1250 1282
rect 1262 1168 1266 1172
rect 1094 268 1098 272
rect 1134 338 1138 342
rect 1150 328 1154 332
rect 1134 78 1138 82
rect 1262 868 1266 872
rect 1342 1288 1346 1292
rect 1334 1138 1338 1142
rect 1222 58 1226 62
rect 1238 298 1242 302
rect 1294 668 1298 672
rect 1318 298 1322 302
rect 1318 268 1322 272
rect 1370 1803 1374 1807
rect 1377 1803 1378 1807
rect 1378 1803 1381 1807
rect 1382 1738 1386 1742
rect 1370 1603 1374 1607
rect 1377 1603 1378 1607
rect 1378 1603 1381 1607
rect 1370 1403 1374 1407
rect 1377 1403 1378 1407
rect 1378 1403 1381 1407
rect 1370 1203 1374 1207
rect 1377 1203 1378 1207
rect 1378 1203 1381 1207
rect 1370 1003 1374 1007
rect 1377 1003 1378 1007
rect 1378 1003 1381 1007
rect 1462 2358 1466 2362
rect 1470 2178 1474 2182
rect 1526 2718 1530 2722
rect 1446 1968 1450 1972
rect 1406 1458 1410 1462
rect 1414 1268 1418 1272
rect 1518 2348 1522 2352
rect 1494 1728 1498 1732
rect 1462 1138 1466 1142
rect 1398 948 1402 952
rect 1366 938 1370 942
rect 1370 803 1374 807
rect 1377 803 1378 807
rect 1378 803 1381 807
rect 1370 603 1374 607
rect 1377 603 1378 607
rect 1378 603 1381 607
rect 1370 403 1374 407
rect 1377 403 1378 407
rect 1378 403 1381 407
rect 1370 203 1374 207
rect 1377 203 1378 207
rect 1378 203 1381 207
rect 1406 868 1410 872
rect 1462 748 1466 752
rect 1406 618 1410 622
rect 1542 2138 1546 2142
rect 1702 3448 1706 3452
rect 1718 3438 1722 3442
rect 1670 3338 1674 3342
rect 1702 3328 1706 3332
rect 1774 3338 1778 3342
rect 1646 2768 1650 2772
rect 1614 2738 1618 2742
rect 1582 2438 1586 2442
rect 1598 2278 1602 2282
rect 1678 2828 1682 2832
rect 1630 2328 1634 2332
rect 1630 2238 1634 2242
rect 1630 2158 1634 2162
rect 1558 1688 1562 1692
rect 1542 858 1546 862
rect 1526 778 1530 782
rect 1518 768 1522 772
rect 1526 768 1530 772
rect 1566 748 1570 752
rect 1422 338 1426 342
rect 1398 188 1402 192
rect 1446 128 1450 132
rect 1446 58 1450 62
rect 1478 68 1482 72
rect 1622 1868 1626 1872
rect 1606 1318 1610 1322
rect 1590 788 1594 792
rect 1670 2048 1674 2052
rect 1646 1678 1650 1682
rect 1638 818 1642 822
rect 1694 2258 1698 2262
rect 1686 2148 1690 2152
rect 1726 2428 1730 2432
rect 1710 1958 1714 1962
rect 1678 1838 1682 1842
rect 1702 1838 1706 1842
rect 1678 1548 1682 1552
rect 1630 548 1634 552
rect 1526 338 1530 342
rect 1550 268 1554 272
rect 1590 268 1594 272
rect 1582 138 1586 142
rect 1654 148 1658 152
rect 1926 3648 1930 3652
rect 1874 3503 1878 3507
rect 1881 3503 1882 3507
rect 1882 3503 1885 3507
rect 1838 3468 1842 3472
rect 1806 3318 1810 3322
rect 1874 3303 1878 3307
rect 1881 3303 1882 3307
rect 1882 3303 1885 3307
rect 1874 3103 1878 3107
rect 1881 3103 1882 3107
rect 1882 3103 1885 3107
rect 1822 2588 1826 2592
rect 1766 2438 1770 2442
rect 1806 2358 1810 2362
rect 1742 2268 1746 2272
rect 1734 2038 1738 2042
rect 1710 1518 1714 1522
rect 1710 1458 1714 1462
rect 1734 1758 1738 1762
rect 1750 1568 1754 1572
rect 1726 1438 1730 1442
rect 1702 1248 1706 1252
rect 1694 1148 1698 1152
rect 1694 138 1698 142
rect 1766 2058 1770 2062
rect 1790 1718 1794 1722
rect 1766 1478 1770 1482
rect 1798 1638 1802 1642
rect 1790 1518 1794 1522
rect 1782 1388 1786 1392
rect 1874 2903 1878 2907
rect 1881 2903 1882 2907
rect 1882 2903 1885 2907
rect 1894 2758 1898 2762
rect 1874 2703 1878 2707
rect 1881 2703 1882 2707
rect 1882 2703 1885 2707
rect 1894 2648 1898 2652
rect 1874 2503 1878 2507
rect 1881 2503 1882 2507
rect 1882 2503 1885 2507
rect 1870 2338 1874 2342
rect 1902 2338 1906 2342
rect 1862 2318 1866 2322
rect 1874 2303 1878 2307
rect 1881 2303 1882 2307
rect 1882 2303 1885 2307
rect 1874 2103 1878 2107
rect 1881 2103 1882 2107
rect 1882 2103 1885 2107
rect 1874 1903 1878 1907
rect 1881 1903 1882 1907
rect 1882 1903 1885 1907
rect 1902 2178 1906 2182
rect 1902 1908 1906 1912
rect 1958 3468 1962 3472
rect 1974 3248 1978 3252
rect 1990 3088 1994 3092
rect 1942 2728 1946 2732
rect 1966 2868 1970 2872
rect 2054 3348 2058 3352
rect 2030 2858 2034 2862
rect 1990 2788 1994 2792
rect 2054 2728 2058 2732
rect 2062 2668 2066 2672
rect 1950 2578 1954 2582
rect 2030 2548 2034 2552
rect 1934 2278 1938 2282
rect 1934 1928 1938 1932
rect 1874 1703 1878 1707
rect 1881 1703 1882 1707
rect 1882 1703 1885 1707
rect 1838 1388 1842 1392
rect 1790 1288 1794 1292
rect 1798 1268 1802 1272
rect 1822 1328 1826 1332
rect 1862 1528 1866 1532
rect 1874 1503 1878 1507
rect 1881 1503 1882 1507
rect 1882 1503 1885 1507
rect 1846 1268 1850 1272
rect 1798 958 1802 962
rect 1798 878 1802 882
rect 1782 748 1786 752
rect 1798 148 1802 152
rect 1902 1458 1906 1462
rect 1902 1378 1906 1382
rect 1878 1338 1882 1342
rect 1874 1303 1878 1307
rect 1881 1303 1882 1307
rect 1882 1303 1885 1307
rect 1878 1268 1882 1272
rect 1874 1103 1878 1107
rect 1881 1103 1882 1107
rect 1882 1103 1885 1107
rect 1874 903 1878 907
rect 1881 903 1882 907
rect 1882 903 1885 907
rect 1942 1618 1946 1622
rect 1990 2168 1994 2172
rect 1926 1538 1930 1542
rect 1926 1498 1930 1502
rect 1934 1088 1938 1092
rect 1934 878 1938 882
rect 1862 768 1866 772
rect 1874 703 1878 707
rect 1881 703 1882 707
rect 1882 703 1885 707
rect 1822 668 1826 672
rect 1874 503 1878 507
rect 1881 503 1882 507
rect 1882 503 1885 507
rect 1902 348 1906 352
rect 1874 303 1878 307
rect 1881 303 1882 307
rect 1882 303 1885 307
rect 1862 128 1866 132
rect 1874 103 1878 107
rect 1881 103 1882 107
rect 1882 103 1885 107
rect 1894 68 1898 72
rect 1958 1428 1962 1432
rect 2006 1918 2010 1922
rect 2038 2328 2042 2332
rect 2022 1958 2026 1962
rect 1982 1578 1986 1582
rect 1990 1528 1994 1532
rect 2118 2448 2122 2452
rect 2134 2488 2138 2492
rect 2094 2248 2098 2252
rect 2078 2188 2082 2192
rect 2062 2048 2066 2052
rect 2046 1718 2050 1722
rect 2062 1688 2066 1692
rect 2046 1668 2050 1672
rect 1998 1488 2002 1492
rect 2014 1478 2018 1482
rect 2006 1468 2010 1472
rect 1998 1438 2002 1442
rect 1974 1068 1978 1072
rect 1982 988 1986 992
rect 2062 1548 2066 1552
rect 2062 1528 2066 1532
rect 2062 1418 2066 1422
rect 2038 1338 2042 1342
rect 2030 1218 2034 1222
rect 2030 968 2034 972
rect 1974 218 1978 222
rect 1990 188 1994 192
rect 2038 618 2042 622
rect 2142 2458 2146 2462
rect 2086 1968 2090 1972
rect 2086 1948 2090 1952
rect 2078 1558 2082 1562
rect 2102 1948 2106 1952
rect 2270 3668 2274 3672
rect 2518 3668 2522 3672
rect 2230 3468 2234 3472
rect 2190 3458 2194 3462
rect 2230 3448 2234 3452
rect 2278 3248 2282 3252
rect 2134 1948 2138 1952
rect 2094 1538 2098 1542
rect 2086 1528 2090 1532
rect 2142 1728 2146 1732
rect 2142 1258 2146 1262
rect 2078 908 2082 912
rect 2070 348 2074 352
rect 2094 78 2098 82
rect 2246 2858 2250 2862
rect 2318 3468 2322 3472
rect 2310 3458 2314 3462
rect 2394 3603 2398 3607
rect 2401 3603 2402 3607
rect 2402 3603 2405 3607
rect 2394 3403 2398 3407
rect 2401 3403 2402 3407
rect 2402 3403 2405 3407
rect 2310 3088 2314 3092
rect 2394 3203 2398 3207
rect 2401 3203 2402 3207
rect 2402 3203 2405 3207
rect 2262 2668 2266 2672
rect 2262 2658 2266 2662
rect 2294 2558 2298 2562
rect 2190 2228 2194 2232
rect 2198 1688 2202 1692
rect 2174 1448 2178 1452
rect 2174 1268 2178 1272
rect 2174 1248 2178 1252
rect 2190 1478 2194 1482
rect 2198 1468 2202 1472
rect 2222 2248 2226 2252
rect 2222 1888 2226 1892
rect 2294 2268 2298 2272
rect 2286 2258 2290 2262
rect 2182 1078 2186 1082
rect 2134 128 2138 132
rect 2238 1338 2242 1342
rect 2166 128 2170 132
rect 2286 1938 2290 1942
rect 2318 2448 2322 2452
rect 2394 3003 2398 3007
rect 2401 3003 2402 3007
rect 2402 3003 2405 3007
rect 2394 2803 2398 2807
rect 2401 2803 2402 2807
rect 2402 2803 2405 2807
rect 2406 2648 2410 2652
rect 2394 2603 2398 2607
rect 2401 2603 2402 2607
rect 2402 2603 2405 2607
rect 2394 2403 2398 2407
rect 2401 2403 2402 2407
rect 2402 2403 2405 2407
rect 2278 1728 2282 1732
rect 2318 1538 2322 1542
rect 2286 1438 2290 1442
rect 2270 1348 2274 1352
rect 2302 178 2306 182
rect 2358 2218 2362 2222
rect 2394 2203 2398 2207
rect 2401 2203 2402 2207
rect 2402 2203 2405 2207
rect 2394 2003 2398 2007
rect 2401 2003 2402 2007
rect 2402 2003 2405 2007
rect 2382 1918 2386 1922
rect 2394 1803 2398 1807
rect 2401 1803 2402 1807
rect 2402 1803 2405 1807
rect 2350 1728 2354 1732
rect 2394 1603 2398 1607
rect 2401 1603 2402 1607
rect 2402 1603 2405 1607
rect 2394 1403 2398 1407
rect 2401 1403 2402 1407
rect 2402 1403 2405 1407
rect 2382 1328 2386 1332
rect 2374 1288 2378 1292
rect 2382 1278 2386 1282
rect 2394 1203 2398 1207
rect 2401 1203 2402 1207
rect 2402 1203 2405 1207
rect 2394 1003 2398 1007
rect 2401 1003 2402 1007
rect 2402 1003 2405 1007
rect 2334 948 2338 952
rect 2358 868 2362 872
rect 2390 858 2394 862
rect 2394 803 2398 807
rect 2401 803 2402 807
rect 2402 803 2405 807
rect 2374 738 2378 742
rect 2394 603 2398 607
rect 2401 603 2402 607
rect 2402 603 2405 607
rect 2358 468 2362 472
rect 2326 458 2330 462
rect 2558 2868 2562 2872
rect 2606 3338 2610 3342
rect 2486 2538 2490 2542
rect 2454 1788 2458 1792
rect 2470 1728 2474 1732
rect 2470 1278 2474 1282
rect 2446 988 2450 992
rect 2462 858 2466 862
rect 2462 738 2466 742
rect 2462 728 2466 732
rect 2422 708 2426 712
rect 2394 403 2398 407
rect 2401 403 2402 407
rect 2402 403 2405 407
rect 2398 328 2402 332
rect 2394 203 2398 207
rect 2401 203 2402 207
rect 2402 203 2405 207
rect 2382 118 2386 122
rect 2502 2438 2506 2442
rect 2638 2588 2642 2592
rect 2622 2448 2626 2452
rect 2502 2348 2506 2352
rect 2494 1728 2498 1732
rect 2510 1678 2514 1682
rect 2494 1528 2498 1532
rect 2478 358 2482 362
rect 2470 318 2474 322
rect 2502 958 2506 962
rect 2614 2048 2618 2052
rect 2614 2038 2618 2042
rect 2526 1358 2530 1362
rect 2614 1748 2618 1752
rect 2566 1558 2570 1562
rect 2582 1318 2586 1322
rect 2566 1258 2570 1262
rect 2622 958 2626 962
rect 2614 908 2618 912
rect 2582 868 2586 872
rect 2518 758 2522 762
rect 2502 718 2506 722
rect 2574 708 2578 712
rect 2614 688 2618 692
rect 2446 168 2450 172
rect 2478 148 2482 152
rect 2534 128 2538 132
rect 2502 68 2506 72
rect 2446 58 2450 62
rect 2646 2158 2650 2162
rect 2670 2838 2674 2842
rect 2702 2488 2706 2492
rect 2906 3503 2910 3507
rect 2913 3503 2914 3507
rect 2914 3503 2917 3507
rect 2894 3338 2898 3342
rect 2906 3303 2910 3307
rect 2913 3303 2914 3307
rect 2914 3303 2917 3307
rect 2906 3103 2910 3107
rect 2913 3103 2914 3107
rect 2914 3103 2917 3107
rect 2906 2903 2910 2907
rect 2913 2903 2914 2907
rect 2914 2903 2917 2907
rect 2830 2838 2834 2842
rect 2982 3068 2986 3072
rect 2894 2728 2898 2732
rect 2790 2548 2794 2552
rect 2878 2548 2882 2552
rect 2806 2138 2810 2142
rect 2774 2048 2778 2052
rect 2782 1908 2786 1912
rect 2670 1548 2674 1552
rect 2766 1878 2770 1882
rect 2750 1638 2754 1642
rect 2886 2348 2890 2352
rect 2822 2068 2826 2072
rect 2694 1468 2698 1472
rect 2670 1058 2674 1062
rect 2638 968 2642 972
rect 2638 878 2642 882
rect 2662 728 2666 732
rect 2670 688 2674 692
rect 2742 1458 2746 1462
rect 2774 1058 2778 1062
rect 2782 948 2786 952
rect 2702 938 2706 942
rect 2814 878 2818 882
rect 2814 718 2818 722
rect 2806 648 2810 652
rect 2906 2703 2910 2707
rect 2913 2703 2914 2707
rect 2914 2703 2917 2707
rect 2966 2658 2970 2662
rect 3022 3068 3026 3072
rect 2906 2503 2910 2507
rect 2913 2503 2914 2507
rect 2914 2503 2917 2507
rect 3046 2958 3050 2962
rect 3206 3058 3210 3062
rect 3142 2858 3146 2862
rect 3206 2778 3210 2782
rect 3062 2758 3066 2762
rect 3230 2928 3234 2932
rect 3198 2558 3202 2562
rect 3254 2858 3258 2862
rect 3418 3603 3422 3607
rect 3425 3603 3426 3607
rect 3426 3603 3429 3607
rect 3418 3403 3422 3407
rect 3425 3403 3426 3407
rect 3426 3403 3429 3407
rect 3930 3503 3934 3507
rect 3937 3503 3938 3507
rect 3938 3503 3941 3507
rect 3630 3398 3634 3402
rect 3418 3203 3422 3207
rect 3425 3203 3426 3207
rect 3426 3203 3429 3207
rect 3418 3003 3422 3007
rect 3425 3003 3426 3007
rect 3426 3003 3429 3007
rect 3430 2938 3434 2942
rect 3418 2803 3422 2807
rect 3425 2803 3426 2807
rect 3426 2803 3429 2807
rect 3390 2738 3394 2742
rect 3462 2928 3466 2932
rect 3574 2958 3578 2962
rect 3526 2648 3530 2652
rect 2990 2428 2994 2432
rect 3142 2358 3146 2362
rect 2906 2303 2910 2307
rect 2913 2303 2914 2307
rect 2914 2303 2917 2307
rect 2906 2103 2910 2107
rect 2913 2103 2914 2107
rect 2914 2103 2917 2107
rect 2942 2018 2946 2022
rect 2942 1928 2946 1932
rect 2934 1918 2938 1922
rect 2906 1903 2910 1907
rect 2913 1903 2914 1907
rect 2914 1903 2917 1907
rect 2926 1878 2930 1882
rect 2906 1703 2910 1707
rect 2913 1703 2914 1707
rect 2914 1703 2917 1707
rect 2906 1503 2910 1507
rect 2913 1503 2914 1507
rect 2914 1503 2917 1507
rect 2906 1303 2910 1307
rect 2913 1303 2914 1307
rect 2914 1303 2917 1307
rect 2902 1258 2906 1262
rect 2906 1103 2910 1107
rect 2913 1103 2914 1107
rect 2914 1103 2917 1107
rect 2906 903 2910 907
rect 2913 903 2914 907
rect 2914 903 2917 907
rect 2934 1678 2938 1682
rect 2966 1388 2970 1392
rect 2906 703 2910 707
rect 2913 703 2914 707
rect 2914 703 2917 707
rect 2906 503 2910 507
rect 2913 503 2914 507
rect 2914 503 2917 507
rect 2906 303 2910 307
rect 2913 303 2914 307
rect 2914 303 2917 307
rect 2766 278 2770 282
rect 2854 158 2858 162
rect 2734 138 2738 142
rect 2862 138 2866 142
rect 2906 103 2910 107
rect 2913 103 2914 107
rect 2914 103 2917 107
rect 2782 78 2786 82
rect 2814 78 2818 82
rect 2830 78 2834 82
rect 3038 2148 3042 2152
rect 3062 2058 3066 2062
rect 3006 1948 3010 1952
rect 3014 1668 3018 1672
rect 3110 2138 3114 2142
rect 3086 1938 3090 1942
rect 3190 2038 3194 2042
rect 3214 2038 3218 2042
rect 3418 2603 3422 2607
rect 3425 2603 3426 2607
rect 3426 2603 3429 2607
rect 3534 2548 3538 2552
rect 3638 2538 3642 2542
rect 3418 2403 3422 2407
rect 3425 2403 3426 2407
rect 3426 2403 3429 2407
rect 3262 2358 3266 2362
rect 3590 2268 3594 2272
rect 3418 2203 3422 2207
rect 3425 2203 3426 2207
rect 3426 2203 3429 2207
rect 3318 2148 3322 2152
rect 3270 2138 3274 2142
rect 3406 2068 3410 2072
rect 3418 2003 3422 2007
rect 3425 2003 3426 2007
rect 3426 2003 3429 2007
rect 3342 1938 3346 1942
rect 3038 1538 3042 1542
rect 2998 1358 3002 1362
rect 3006 1258 3010 1262
rect 3078 1258 3082 1262
rect 3286 1478 3290 1482
rect 3158 1418 3162 1422
rect 3382 1548 3386 1552
rect 3326 1438 3330 1442
rect 3374 1428 3378 1432
rect 3206 1378 3210 1382
rect 3302 1268 3306 1272
rect 3418 1803 3422 1807
rect 3425 1803 3426 1807
rect 3426 1803 3429 1807
rect 3406 1768 3410 1772
rect 3494 2068 3498 2072
rect 3478 1658 3482 1662
rect 3418 1603 3422 1607
rect 3425 1603 3426 1607
rect 3426 1603 3429 1607
rect 3510 1948 3514 1952
rect 3598 2158 3602 2162
rect 3582 1938 3586 1942
rect 3518 1548 3522 1552
rect 3502 1518 3506 1522
rect 3510 1478 3514 1482
rect 3418 1403 3422 1407
rect 3425 1403 3426 1407
rect 3426 1403 3429 1407
rect 3418 1203 3422 1207
rect 3425 1203 3426 1207
rect 3426 1203 3429 1207
rect 3718 2948 3722 2952
rect 3750 2788 3754 2792
rect 3694 1928 3698 1932
rect 3590 1918 3594 1922
rect 3718 2088 3722 2092
rect 3526 1348 3530 1352
rect 3542 1338 3546 1342
rect 3118 868 3122 872
rect 3102 738 3106 742
rect 3166 678 3170 682
rect 3418 1003 3422 1007
rect 3425 1003 3426 1007
rect 3426 1003 3429 1007
rect 3478 868 3482 872
rect 3418 803 3422 807
rect 3425 803 3426 807
rect 3426 803 3429 807
rect 3254 728 3258 732
rect 3418 603 3422 607
rect 3425 603 3426 607
rect 3426 603 3429 607
rect 3214 468 3218 472
rect 2958 158 2962 162
rect 2942 78 2946 82
rect 2982 138 2986 142
rect 3078 238 3082 242
rect 3078 128 3082 132
rect 3110 338 3114 342
rect 3166 238 3170 242
rect 3150 148 3154 152
rect 3150 68 3154 72
rect 3418 403 3422 407
rect 3425 403 3426 407
rect 3426 403 3429 407
rect 3286 278 3290 282
rect 3238 258 3242 262
rect 3270 118 3274 122
rect 3366 328 3370 332
rect 3342 128 3346 132
rect 3350 108 3354 112
rect 3350 88 3354 92
rect 3478 318 3482 322
rect 3374 258 3378 262
rect 3438 218 3442 222
rect 3418 203 3422 207
rect 3425 203 3426 207
rect 3426 203 3429 207
rect 3390 128 3394 132
rect 3358 68 3362 72
rect 3414 58 3418 62
rect 3518 738 3522 742
rect 3558 1658 3562 1662
rect 3694 1568 3698 1572
rect 3726 1538 3730 1542
rect 3950 3398 3954 3402
rect 3930 3303 3934 3307
rect 3937 3303 3938 3307
rect 3938 3303 3941 3307
rect 3930 3103 3934 3107
rect 3937 3103 3938 3107
rect 3938 3103 3941 3107
rect 3846 3058 3850 3062
rect 3930 2903 3934 2907
rect 3937 2903 3938 2907
rect 3938 2903 3941 2907
rect 3878 2748 3882 2752
rect 3958 2748 3962 2752
rect 3886 2738 3890 2742
rect 3930 2703 3934 2707
rect 3937 2703 3938 2707
rect 3938 2703 3941 2707
rect 3930 2503 3934 2507
rect 3937 2503 3938 2507
rect 3938 2503 3941 2507
rect 3930 2303 3934 2307
rect 3937 2303 3938 2307
rect 3938 2303 3941 2307
rect 3830 2128 3834 2132
rect 3910 2128 3914 2132
rect 3930 2103 3934 2107
rect 3937 2103 3938 2107
rect 3938 2103 3941 2107
rect 3870 1888 3874 1892
rect 3814 1688 3818 1692
rect 3930 1903 3934 1907
rect 3937 1903 3938 1907
rect 3938 1903 3941 1907
rect 3930 1703 3934 1707
rect 3937 1703 3938 1707
rect 3938 1703 3941 1707
rect 3930 1503 3934 1507
rect 3937 1503 3938 1507
rect 3938 1503 3941 1507
rect 3790 1448 3794 1452
rect 3930 1303 3934 1307
rect 3937 1303 3938 1307
rect 3938 1303 3941 1307
rect 3950 1288 3954 1292
rect 3982 2068 3986 2072
rect 4366 3468 4370 3472
rect 4334 3458 4338 3462
rect 4442 3603 4446 3607
rect 4449 3603 4450 3607
rect 4450 3603 4453 3607
rect 4486 3478 4490 3482
rect 4566 3478 4570 3482
rect 4606 3468 4610 3472
rect 4382 3458 4386 3462
rect 4442 3403 4446 3407
rect 4449 3403 4450 3407
rect 4450 3403 4453 3407
rect 4442 3203 4446 3207
rect 4449 3203 4450 3207
rect 4450 3203 4453 3207
rect 4678 3358 4682 3362
rect 4954 3503 4958 3507
rect 4961 3503 4962 3507
rect 4962 3503 4965 3507
rect 5022 3358 5026 3362
rect 4894 3278 4898 3282
rect 4954 3303 4958 3307
rect 4961 3303 4962 3307
rect 4962 3303 4965 3307
rect 4950 3278 4954 3282
rect 4926 3268 4930 3272
rect 4958 3268 4962 3272
rect 4954 3103 4958 3107
rect 4961 3103 4962 3107
rect 4962 3103 4965 3107
rect 4442 3003 4446 3007
rect 4449 3003 4450 3007
rect 4450 3003 4453 3007
rect 4954 2903 4958 2907
rect 4961 2903 4962 2907
rect 4962 2903 4965 2907
rect 4878 2828 4882 2832
rect 4442 2803 4446 2807
rect 4449 2803 4450 2807
rect 4450 2803 4453 2807
rect 4502 2738 4506 2742
rect 4542 2738 4546 2742
rect 4294 2718 4298 2722
rect 4442 2603 4446 2607
rect 4449 2603 4450 2607
rect 4450 2603 4453 2607
rect 4734 2548 4738 2552
rect 4830 2548 4834 2552
rect 4110 2268 4114 2272
rect 3974 1458 3978 1462
rect 4294 2238 4298 2242
rect 4174 1938 4178 1942
rect 4302 1858 4306 1862
rect 4390 2258 4394 2262
rect 4350 1868 4354 1872
rect 4442 2403 4446 2407
rect 4449 2403 4450 2407
rect 4450 2403 4453 2407
rect 4442 2203 4446 2207
rect 4449 2203 4450 2207
rect 4450 2203 4453 2207
rect 4442 2003 4446 2007
rect 4449 2003 4450 2007
rect 4450 2003 4453 2007
rect 4442 1803 4446 1807
rect 4449 1803 4450 1807
rect 4450 1803 4453 1807
rect 4442 1603 4446 1607
rect 4449 1603 4450 1607
rect 4450 1603 4453 1607
rect 4494 2088 4498 2092
rect 4574 2238 4578 2242
rect 4446 1528 4450 1532
rect 4542 1528 4546 1532
rect 4442 1403 4446 1407
rect 4449 1403 4450 1407
rect 4450 1403 4453 1407
rect 4398 1348 4402 1352
rect 4502 1278 4506 1282
rect 4270 1218 4274 1222
rect 4442 1203 4446 1207
rect 4449 1203 4450 1207
rect 4450 1203 4453 1207
rect 3930 1103 3934 1107
rect 3937 1103 3938 1107
rect 3938 1103 3941 1107
rect 3950 1078 3954 1082
rect 3930 903 3934 907
rect 3937 903 3938 907
rect 3938 903 3941 907
rect 3582 728 3586 732
rect 3550 678 3554 682
rect 3550 468 3554 472
rect 3622 568 3626 572
rect 3654 458 3658 462
rect 3678 458 3682 462
rect 3606 338 3610 342
rect 3590 168 3594 172
rect 3622 108 3626 112
rect 3574 78 3578 82
rect 3606 68 3610 72
rect 3646 58 3650 62
rect 4442 1003 4446 1007
rect 4449 1003 4450 1007
rect 4450 1003 4453 1007
rect 4174 928 4178 932
rect 4222 928 4226 932
rect 4442 803 4446 807
rect 4449 803 4450 807
rect 4450 803 4453 807
rect 4198 768 4202 772
rect 4262 748 4266 752
rect 3930 703 3934 707
rect 3937 703 3938 707
rect 3938 703 3941 707
rect 3958 658 3962 662
rect 3958 568 3962 572
rect 3766 468 3770 472
rect 3930 503 3934 507
rect 3937 503 3938 507
rect 3938 503 3941 507
rect 3734 288 3738 292
rect 3798 278 3802 282
rect 3930 303 3934 307
rect 3937 303 3938 307
rect 3938 303 3941 307
rect 3930 103 3934 107
rect 3937 103 3938 107
rect 3938 103 3941 107
rect 4038 658 4042 662
rect 4102 178 4106 182
rect 4798 2348 4802 2352
rect 4630 2278 4634 2282
rect 4686 2278 4690 2282
rect 4742 2278 4746 2282
rect 4718 2258 4722 2262
rect 4718 2058 4722 2062
rect 4734 1148 4738 1152
rect 4742 1088 4746 1092
rect 4262 678 4266 682
rect 4310 648 4314 652
rect 4442 603 4446 607
rect 4449 603 4450 607
rect 4450 603 4453 607
rect 4222 288 4226 292
rect 4442 403 4446 407
rect 4449 403 4450 407
rect 4450 403 4453 407
rect 4334 278 4338 282
rect 4442 203 4446 207
rect 4449 203 4450 207
rect 4450 203 4453 207
rect 4954 2703 4958 2707
rect 4961 2703 4962 2707
rect 4962 2703 4965 2707
rect 4954 2503 4958 2507
rect 4961 2503 4962 2507
rect 4962 2503 4965 2507
rect 4910 2278 4914 2282
rect 4954 2303 4958 2307
rect 4961 2303 4962 2307
rect 4962 2303 4965 2307
rect 4954 2103 4958 2107
rect 4961 2103 4962 2107
rect 4962 2103 4965 2107
rect 4954 1903 4958 1907
rect 4961 1903 4962 1907
rect 4962 1903 4965 1907
rect 4954 1703 4958 1707
rect 4961 1703 4962 1707
rect 4962 1703 4965 1707
rect 4918 1668 4922 1672
rect 4918 1658 4922 1662
rect 4942 1578 4946 1582
rect 4606 748 4610 752
rect 4670 748 4674 752
rect 4954 1503 4958 1507
rect 4961 1503 4962 1507
rect 4962 1503 4965 1507
rect 4954 1303 4958 1307
rect 4961 1303 4962 1307
rect 4962 1303 4965 1307
rect 4954 1103 4958 1107
rect 4961 1103 4962 1107
rect 4962 1103 4965 1107
rect 5102 2728 5106 2732
rect 5110 2638 5114 2642
rect 5086 2348 5090 2352
rect 5070 1768 5074 1772
rect 5078 1618 5082 1622
rect 4954 903 4958 907
rect 4961 903 4962 907
rect 4962 903 4965 907
rect 4954 703 4958 707
rect 4961 703 4962 707
rect 4962 703 4965 707
rect 5142 2638 5146 2642
rect 5142 2218 5146 2222
rect 5302 3648 5306 3652
rect 5198 2408 5202 2412
rect 5198 2168 5202 2172
rect 5182 1958 5186 1962
rect 5198 1958 5202 1962
rect 5198 958 5202 962
rect 5206 788 5210 792
rect 5238 2258 5242 2262
rect 5238 2108 5242 2112
rect 5238 2098 5242 2102
rect 5254 3168 5258 3172
rect 5278 3548 5282 3552
rect 5270 3448 5274 3452
rect 5278 3428 5282 3432
rect 5278 3068 5282 3072
rect 5278 3048 5282 3052
rect 5270 2988 5274 2992
rect 5262 2638 5266 2642
rect 5238 1678 5242 1682
rect 5246 1288 5250 1292
rect 5246 1268 5250 1272
rect 5246 878 5250 882
rect 5254 558 5258 562
rect 4954 503 4958 507
rect 4961 503 4962 507
rect 4962 503 4965 507
rect 4862 468 4866 472
rect 5070 468 5074 472
rect 4942 458 4946 462
rect 5062 458 5066 462
rect 5270 528 5274 532
rect 4954 303 4958 307
rect 4961 303 4962 307
rect 4962 303 4965 307
rect 4954 103 4958 107
rect 4961 103 4962 107
rect 4962 103 4965 107
rect 5302 3068 5306 3072
rect 5302 2668 5306 2672
rect 5302 2628 5306 2632
rect 5302 2578 5306 2582
rect 5294 2568 5298 2572
rect 5294 2518 5298 2522
rect 5310 2258 5314 2262
rect 5310 2148 5314 2152
rect 5310 2138 5314 2142
rect 5310 1668 5314 1672
rect 5310 1488 5314 1492
rect 5310 1148 5314 1152
rect 5310 1088 5314 1092
rect 5310 958 5314 962
rect 5310 858 5314 862
rect 5310 838 5314 842
rect 5302 88 5306 92
rect 346 3 350 7
rect 353 3 354 7
rect 354 3 357 7
rect 1370 3 1374 7
rect 1377 3 1378 7
rect 1378 3 1381 7
rect 2394 3 2398 7
rect 2401 3 2402 7
rect 2402 3 2405 7
rect 3418 3 3422 7
rect 3425 3 3426 7
rect 3426 3 3429 7
rect 4442 3 4446 7
rect 4449 3 4450 7
rect 4450 3 4453 7
<< metal5 >>
rect 862 3703 865 3707
rect 862 3702 866 3703
rect 1878 3703 1881 3707
rect 1878 3702 1882 3703
rect 2910 3703 2913 3707
rect 2910 3702 2914 3703
rect 3934 3703 3937 3707
rect 3934 3702 3938 3703
rect 4958 3703 4961 3707
rect 4958 3702 4962 3703
rect 1794 3678 1974 3681
rect 946 3668 966 3671
rect 1210 3668 1358 3671
rect 2274 3668 2518 3671
rect 1514 3648 1622 3651
rect 1930 3648 5302 3651
rect 350 3603 353 3607
rect 350 3602 354 3603
rect 1374 3603 1377 3607
rect 1374 3602 1378 3603
rect 2398 3603 2401 3607
rect 2398 3602 2402 3603
rect 3422 3603 3425 3607
rect 3422 3602 3426 3603
rect 4446 3603 4449 3607
rect 4446 3602 4450 3603
rect 1098 3548 1150 3551
rect 5235 3548 5278 3551
rect 862 3503 865 3507
rect 862 3502 866 3503
rect 1878 3503 1881 3507
rect 1878 3502 1882 3503
rect 2910 3503 2913 3507
rect 2910 3502 2914 3503
rect 3934 3503 3937 3507
rect 3934 3502 3938 3503
rect 4958 3503 4961 3507
rect 4958 3502 4962 3503
rect 4490 3478 4566 3481
rect 1842 3468 1958 3471
rect 2234 3468 2318 3471
rect 4370 3468 4606 3471
rect 2194 3458 2310 3461
rect 4338 3458 4382 3461
rect 5267 3458 5273 3461
rect 5270 3452 5273 3458
rect 1706 3448 2230 3451
rect 1546 3438 1718 3441
rect 5278 3432 5281 3437
rect 350 3403 353 3407
rect 350 3402 354 3403
rect 1374 3403 1377 3407
rect 1374 3402 1378 3403
rect 2398 3403 2401 3407
rect 2398 3402 2402 3403
rect 3422 3403 3425 3407
rect 3422 3402 3426 3403
rect 4446 3403 4449 3407
rect 4446 3402 4450 3403
rect 3634 3398 3950 3401
rect 530 3368 582 3371
rect 1186 3358 1254 3361
rect 4682 3358 5022 3361
rect 1026 3348 1270 3351
rect 1474 3348 2054 3351
rect 946 3338 1366 3341
rect 1674 3338 1774 3341
rect 2610 3338 2894 3341
rect 1186 3328 1350 3331
rect 1466 3328 1702 3331
rect 1418 3318 1806 3321
rect 862 3303 865 3307
rect 862 3302 866 3303
rect 1878 3303 1881 3307
rect 1878 3302 1882 3303
rect 2910 3303 2913 3307
rect 2910 3302 2914 3303
rect 3934 3303 3937 3307
rect 3934 3302 3938 3303
rect 4958 3303 4961 3307
rect 4958 3302 4962 3303
rect 906 3298 950 3301
rect 818 3288 958 3291
rect 1074 3288 1254 3291
rect 4898 3278 4950 3281
rect 4930 3268 4958 3271
rect 906 3258 1046 3261
rect 1978 3248 2278 3251
rect 350 3203 353 3207
rect 350 3202 354 3203
rect 1374 3203 1377 3207
rect 1374 3202 1378 3203
rect 2398 3203 2401 3207
rect 2398 3202 2402 3203
rect 3422 3203 3425 3207
rect 3422 3202 3426 3203
rect 4446 3203 4449 3207
rect 4446 3202 4450 3203
rect 5251 3168 5254 3171
rect 570 3138 641 3141
rect 638 3132 641 3138
rect 862 3103 865 3107
rect 862 3102 866 3103
rect 1878 3103 1881 3107
rect 1878 3102 1882 3103
rect 2910 3103 2913 3107
rect 2910 3102 2914 3103
rect 3934 3103 3937 3107
rect 3934 3102 3938 3103
rect 4958 3103 4961 3107
rect 4958 3102 4962 3103
rect 1994 3088 2310 3091
rect 842 3068 1206 3071
rect 2986 3068 3022 3071
rect 5282 3068 5293 3071
rect 5306 3068 5309 3071
rect 3210 3058 3846 3061
rect 5278 3052 5281 3057
rect 1226 3048 1318 3051
rect 350 3003 353 3007
rect 350 3002 354 3003
rect 1374 3003 1377 3007
rect 1374 3002 1378 3003
rect 2398 3003 2401 3007
rect 2398 3002 2402 3003
rect 3422 3003 3425 3007
rect 3422 3002 3426 3003
rect 4446 3003 4449 3007
rect 4446 3002 4450 3003
rect 5274 2988 5277 2991
rect 3050 2958 3574 2961
rect 3718 2941 3721 2948
rect 3434 2938 3721 2941
rect 3234 2928 3462 2931
rect 866 2918 1422 2921
rect 862 2903 865 2907
rect 862 2902 866 2903
rect 1878 2903 1881 2907
rect 1878 2902 1882 2903
rect 2910 2903 2913 2907
rect 2910 2902 2914 2903
rect 3934 2903 3937 2907
rect 3934 2902 3938 2903
rect 4958 2903 4961 2907
rect 4958 2902 4962 2903
rect 1970 2868 2558 2871
rect 2034 2858 2246 2861
rect 3146 2858 3254 2861
rect 2674 2838 2830 2841
rect 1682 2828 4878 2831
rect 350 2803 353 2807
rect 350 2802 354 2803
rect 1374 2803 1377 2807
rect 1374 2802 1378 2803
rect 2398 2803 2401 2807
rect 2398 2802 2402 2803
rect 3422 2803 3425 2807
rect 3422 2802 3426 2803
rect 4446 2803 4449 2807
rect 4446 2802 4450 2803
rect 1994 2788 3750 2791
rect 1646 2778 3206 2781
rect 1646 2772 1649 2778
rect 1898 2758 3062 2761
rect 3882 2748 3958 2751
rect 666 2738 1614 2741
rect 3394 2738 3886 2741
rect 4506 2738 4542 2741
rect 1946 2728 2054 2731
rect 2898 2728 5102 2731
rect 1530 2718 4294 2721
rect 862 2703 865 2707
rect 862 2702 866 2703
rect 1878 2703 1881 2707
rect 1878 2702 1882 2703
rect 2910 2703 2913 2707
rect 2910 2702 2914 2703
rect 3934 2703 3937 2707
rect 3934 2702 3938 2703
rect 4958 2703 4961 2707
rect 4958 2702 4962 2703
rect 994 2678 1054 2681
rect 5299 2678 5305 2681
rect 5302 2672 5305 2678
rect 2066 2668 2262 2671
rect 2266 2658 2966 2661
rect 1082 2648 1894 2651
rect 2410 2648 3526 2651
rect 1090 2638 1126 2641
rect 5114 2638 5142 2641
rect 5266 2638 5277 2641
rect 5283 2628 5302 2631
rect 22 2601 25 2608
rect 350 2603 353 2607
rect 350 2602 354 2603
rect 1374 2603 1377 2607
rect 1374 2602 1378 2603
rect 2398 2603 2401 2607
rect 2398 2602 2402 2603
rect 3422 2603 3425 2607
rect 3422 2602 3426 2603
rect 4446 2603 4449 2607
rect 4446 2602 4450 2603
rect 22 2598 110 2601
rect 1826 2588 2638 2591
rect 634 2578 1950 2581
rect 5306 2578 5309 2581
rect 5298 2568 5309 2571
rect 666 2558 854 2561
rect 2298 2558 3198 2561
rect 2034 2548 2790 2551
rect 2882 2548 3534 2551
rect 4738 2548 4830 2551
rect 146 2538 198 2541
rect 2490 2538 3638 2541
rect 5298 2518 5357 2521
rect 862 2503 865 2507
rect 862 2502 866 2503
rect 1878 2503 1881 2507
rect 1878 2502 1882 2503
rect 2910 2503 2913 2507
rect 2910 2502 2914 2503
rect 3934 2503 3937 2507
rect 3934 2502 3938 2503
rect 4958 2503 4961 2507
rect 4958 2502 4962 2503
rect 2138 2488 2702 2491
rect 2142 2462 2145 2467
rect 2122 2448 2318 2451
rect 2622 2443 2625 2448
rect 1034 2438 1582 2441
rect 1770 2438 2502 2441
rect 1730 2428 2990 2431
rect 5202 2408 5213 2411
rect 350 2403 353 2407
rect 350 2402 354 2403
rect 1374 2403 1377 2407
rect 1374 2402 1378 2403
rect 2398 2403 2401 2407
rect 2398 2402 2402 2403
rect 3422 2403 3425 2407
rect 3422 2402 3426 2403
rect 4446 2403 4449 2407
rect 4446 2402 4450 2403
rect 650 2368 1390 2371
rect 906 2358 1070 2361
rect 1466 2358 1806 2361
rect 3146 2358 3262 2361
rect 1522 2348 2502 2351
rect 2506 2348 2886 2351
rect 4802 2348 5086 2351
rect 1874 2338 1902 2341
rect 1634 2328 2038 2331
rect 714 2318 1862 2321
rect 862 2303 865 2307
rect 862 2302 866 2303
rect 1878 2303 1881 2307
rect 1878 2302 1882 2303
rect 2910 2303 2913 2307
rect 2910 2302 2914 2303
rect 3934 2303 3937 2307
rect 3934 2302 3938 2303
rect 4958 2303 4961 2307
rect 4958 2302 4962 2303
rect 194 2288 1030 2291
rect 1602 2278 1934 2281
rect 4634 2278 4686 2281
rect 4746 2278 4910 2281
rect 1746 2268 2294 2271
rect 3594 2268 4110 2271
rect 1698 2258 2286 2261
rect 4394 2258 4718 2261
rect 5242 2258 5310 2261
rect 2098 2248 2222 2251
rect 962 2238 1630 2241
rect 4298 2238 4574 2241
rect 1106 2228 2190 2231
rect 2362 2218 5142 2221
rect 22 2208 118 2211
rect 22 2202 25 2208
rect 350 2203 353 2207
rect 350 2202 354 2203
rect 1374 2203 1377 2207
rect 1374 2202 1378 2203
rect 2398 2203 2401 2207
rect 2398 2202 2402 2203
rect 3422 2203 3425 2207
rect 3422 2202 3426 2203
rect 4446 2203 4449 2207
rect 4446 2202 4450 2203
rect 1034 2188 2078 2191
rect 1474 2178 1902 2181
rect 1338 2168 1990 2171
rect 5202 2168 5213 2171
rect 498 2158 1630 2161
rect 2650 2158 3598 2161
rect 1266 2148 1686 2151
rect 3042 2148 3318 2151
rect 5219 2148 5310 2151
rect 1546 2138 2806 2141
rect 3114 2138 3270 2141
rect 5283 2138 5310 2141
rect 106 2128 1094 2131
rect 3834 2128 3910 2131
rect 5235 2128 5277 2131
rect 370 2118 1078 2121
rect 862 2103 865 2107
rect 862 2102 866 2103
rect 1878 2103 1881 2107
rect 1878 2102 1882 2103
rect 2910 2103 2913 2107
rect 2910 2102 2914 2103
rect 3934 2103 3937 2107
rect 3934 2102 3938 2103
rect 5235 2108 5238 2111
rect 4958 2103 4961 2107
rect 4958 2102 4962 2103
rect 5242 2098 5277 2101
rect 3722 2088 4494 2091
rect 58 2068 302 2071
rect 3410 2068 3494 2071
rect 3986 2068 4721 2071
rect 1346 2058 1766 2061
rect 2822 2061 2825 2068
rect 4718 2062 4721 2068
rect 2822 2058 3062 2061
rect 1674 2048 2062 2051
rect 2618 2048 2774 2051
rect 1250 2038 1734 2041
rect 2618 2038 2621 2041
rect 3194 2038 3214 2041
rect 898 2018 2942 2021
rect 350 2003 353 2007
rect 350 2002 354 2003
rect 1374 2003 1377 2007
rect 1374 2002 1378 2003
rect 2398 2003 2401 2007
rect 2398 2002 2402 2003
rect 3422 2003 3425 2007
rect 3422 2002 3426 2003
rect 4446 2003 4449 2007
rect 4446 2002 4450 2003
rect 1450 1968 2086 1971
rect 1714 1958 2022 1961
rect 5186 1958 5198 1961
rect 2106 1948 2134 1951
rect 3010 1948 3510 1951
rect 2086 1941 2089 1948
rect 2086 1938 2286 1941
rect 3090 1938 3342 1941
rect 3586 1938 4174 1941
rect 1938 1928 2942 1931
rect 2946 1928 3694 1931
rect 2010 1918 2382 1921
rect 2938 1918 3590 1921
rect 1906 1908 2782 1911
rect 862 1903 865 1907
rect 862 1902 866 1903
rect 1878 1903 1881 1907
rect 1878 1902 1882 1903
rect 2910 1903 2913 1907
rect 2910 1902 2914 1903
rect 3934 1903 3937 1907
rect 3934 1902 3938 1903
rect 4958 1903 4961 1907
rect 4958 1902 4962 1903
rect 2226 1888 3870 1891
rect 2770 1878 2926 1881
rect 1290 1868 1622 1871
rect 650 1858 1150 1861
rect 4350 1861 4353 1868
rect 4306 1858 4353 1861
rect 1682 1838 1702 1841
rect 350 1803 353 1807
rect 350 1802 354 1803
rect 1374 1803 1377 1807
rect 1374 1802 1378 1803
rect 2398 1803 2401 1807
rect 2398 1802 2402 1803
rect 3422 1803 3425 1807
rect 3422 1802 3426 1803
rect 4446 1803 4449 1807
rect 4446 1802 4450 1803
rect 1314 1788 2454 1791
rect 922 1768 1142 1771
rect 3410 1768 5070 1771
rect 1218 1758 1734 1761
rect 538 1748 1238 1751
rect 1382 1748 2614 1751
rect 1382 1742 1385 1748
rect 1498 1728 2142 1731
rect 2282 1728 2350 1731
rect 2474 1728 2494 1731
rect 1794 1718 2046 1721
rect 862 1703 865 1707
rect 862 1702 866 1703
rect 1878 1703 1881 1707
rect 1878 1702 1882 1703
rect 2910 1703 2913 1707
rect 2910 1702 2914 1703
rect 3934 1703 3937 1707
rect 3934 1702 3938 1703
rect 4958 1703 4961 1707
rect 4958 1702 4962 1703
rect 698 1688 894 1691
rect 1562 1688 2062 1691
rect 2066 1688 2198 1691
rect 2202 1688 3814 1691
rect 2514 1678 2934 1681
rect 1646 1671 1649 1678
rect 5235 1678 5238 1681
rect 1646 1668 2046 1671
rect 3018 1668 4918 1671
rect 634 1658 686 1661
rect 690 1658 766 1661
rect 3482 1658 3558 1661
rect 5310 1661 5313 1668
rect 4922 1658 5313 1661
rect 1802 1638 2750 1641
rect 1946 1618 5078 1621
rect 858 1608 966 1611
rect 350 1603 353 1607
rect 350 1602 354 1603
rect 1374 1603 1377 1607
rect 1374 1602 1378 1603
rect 2398 1603 2401 1607
rect 2398 1602 2402 1603
rect 3422 1603 3425 1607
rect 3422 1602 3426 1603
rect 4446 1603 4449 1607
rect 4446 1602 4450 1603
rect 1986 1578 4942 1581
rect 1754 1568 3694 1571
rect 106 1558 174 1561
rect 2082 1558 2566 1561
rect 946 1548 1142 1551
rect 2066 1548 2670 1551
rect 3386 1548 3518 1551
rect 1002 1538 1086 1541
rect 1678 1541 1681 1548
rect 1678 1538 1926 1541
rect 2098 1538 2318 1541
rect 3042 1538 3726 1541
rect 1866 1528 1990 1531
rect 2066 1528 2086 1531
rect 2090 1528 2494 1531
rect 4450 1528 4542 1531
rect 1714 1518 1790 1521
rect 1794 1518 3502 1521
rect 862 1503 865 1507
rect 862 1502 866 1503
rect 1878 1503 1881 1507
rect 1878 1502 1882 1503
rect 2910 1503 2913 1507
rect 2910 1502 2914 1503
rect 3934 1503 3937 1507
rect 3934 1502 3938 1503
rect 4958 1503 4961 1507
rect 4958 1502 4962 1503
rect 722 1488 1118 1491
rect 1926 1491 1929 1498
rect 1202 1488 1929 1491
rect 2002 1488 5310 1491
rect 178 1478 254 1481
rect 1194 1478 1766 1481
rect 2018 1478 2190 1481
rect 3290 1478 3510 1481
rect 1306 1468 1334 1471
rect 2010 1468 2198 1471
rect 2202 1468 2694 1471
rect 874 1458 1406 1461
rect 1714 1458 1902 1461
rect 2746 1458 3974 1461
rect 2178 1448 3790 1451
rect 818 1438 1318 1441
rect 1730 1438 1998 1441
rect 2290 1438 3326 1441
rect 1962 1428 3374 1431
rect 2066 1418 3158 1421
rect 350 1403 353 1407
rect 350 1402 354 1403
rect 1374 1403 1377 1407
rect 1374 1402 1378 1403
rect 2398 1403 2401 1407
rect 2398 1402 2402 1403
rect 3422 1403 3425 1407
rect 3422 1402 3426 1403
rect 4446 1403 4449 1407
rect 4446 1402 4450 1403
rect 1786 1388 1838 1391
rect 1842 1388 2966 1391
rect 1906 1378 3206 1381
rect 1066 1358 1118 1361
rect 2530 1358 2998 1361
rect 1178 1348 2270 1351
rect 3530 1348 4398 1351
rect 1882 1338 2038 1341
rect 2242 1338 3542 1341
rect 1826 1328 2382 1331
rect 1610 1318 2582 1321
rect 862 1303 865 1307
rect 862 1302 866 1303
rect 1878 1303 1881 1307
rect 1878 1302 1882 1303
rect 2910 1303 2913 1307
rect 2910 1302 2914 1303
rect 3934 1303 3937 1307
rect 3934 1302 3938 1303
rect 4958 1303 4961 1307
rect 4958 1302 4962 1303
rect 1346 1288 1790 1291
rect 2378 1288 3950 1291
rect 5250 1288 5277 1291
rect 1250 1278 2382 1281
rect 2474 1278 4502 1281
rect 5219 1278 5249 1281
rect 1418 1268 1798 1271
rect 1850 1268 1878 1271
rect 5246 1272 5249 1278
rect 2178 1268 3302 1271
rect 2142 1262 2145 1267
rect 810 1258 862 1261
rect 2570 1258 2902 1261
rect 3010 1258 3078 1261
rect 1706 1248 2174 1251
rect 2034 1218 4270 1221
rect 350 1203 353 1207
rect 350 1202 354 1203
rect 1374 1203 1377 1207
rect 1374 1202 1378 1203
rect 2398 1203 2401 1207
rect 2398 1202 2402 1203
rect 3422 1203 3425 1207
rect 3422 1202 3426 1203
rect 4446 1203 4449 1207
rect 4446 1202 4450 1203
rect 410 1168 1262 1171
rect 1698 1148 4734 1151
rect 4738 1148 5310 1151
rect 1338 1138 1462 1141
rect 862 1103 865 1107
rect 862 1102 866 1103
rect 1878 1103 1881 1107
rect 1878 1102 1882 1103
rect 2910 1103 2913 1107
rect 2910 1102 2914 1103
rect 3934 1103 3937 1107
rect 3934 1102 3938 1103
rect 4958 1103 4961 1107
rect 4958 1102 4962 1103
rect 1938 1088 4742 1091
rect 4746 1088 5310 1091
rect 1974 1078 2182 1081
rect 2186 1078 3950 1081
rect 1974 1072 1977 1078
rect 594 1068 710 1071
rect 2674 1058 2774 1061
rect 350 1003 353 1007
rect 350 1002 354 1003
rect 1374 1003 1377 1007
rect 1374 1002 1378 1003
rect 2398 1003 2401 1007
rect 2398 1002 2402 1003
rect 3422 1003 3425 1007
rect 3422 1002 3426 1003
rect 4446 1003 4449 1007
rect 4446 1002 4450 1003
rect 1986 988 2446 991
rect 2034 968 2638 971
rect 938 958 1038 961
rect 1802 958 2502 961
rect 810 948 1398 951
rect 2622 951 2625 958
rect 2338 948 2625 951
rect 5198 951 5201 958
rect 5310 951 5313 958
rect 2786 948 5313 951
rect 1370 938 2702 941
rect 4178 928 4222 931
rect 2082 908 2614 911
rect 862 903 865 907
rect 862 902 866 903
rect 1878 903 1881 907
rect 1878 902 1882 903
rect 2910 903 2913 907
rect 2910 902 2914 903
rect 3934 903 3937 907
rect 3934 902 3938 903
rect 4958 903 4961 907
rect 4958 902 4962 903
rect 10 888 742 891
rect 546 878 1798 881
rect 1938 878 2638 881
rect 2642 878 2814 881
rect 5246 873 5249 878
rect 1266 868 1406 871
rect 2362 868 2582 871
rect 3122 868 3478 871
rect 1050 858 1542 861
rect 2394 858 2462 861
rect 5314 858 5357 861
rect 5310 842 5313 847
rect 10 818 1638 821
rect 350 803 353 807
rect 350 802 354 803
rect 1374 803 1377 807
rect 1374 802 1378 803
rect 2398 803 2401 807
rect 2398 802 2402 803
rect 3422 803 3425 807
rect 3422 802 3426 803
rect 4446 803 4449 807
rect 4446 802 4450 803
rect 1594 788 5206 791
rect 506 778 1526 781
rect 1510 768 1518 771
rect 1522 768 1526 771
rect 1866 768 4198 771
rect 802 758 2518 761
rect 1466 748 1566 751
rect 1786 748 4262 751
rect 4610 748 4670 751
rect 2378 738 2462 741
rect 3106 738 3518 741
rect 442 728 542 731
rect 546 728 654 731
rect 2466 728 2662 731
rect 3258 728 3582 731
rect 2506 718 2814 721
rect 2426 708 2574 711
rect 862 703 865 707
rect 862 702 866 703
rect 1878 703 1881 707
rect 1878 702 1882 703
rect 2910 703 2913 707
rect 2910 702 2914 703
rect 3934 703 3937 707
rect 3934 702 3938 703
rect 4958 703 4961 707
rect 4958 702 4962 703
rect 562 688 1078 691
rect 2618 688 2670 691
rect 3170 678 3550 681
rect 3554 678 4262 681
rect 1298 668 1822 671
rect 258 658 534 661
rect 3962 658 4038 661
rect 194 648 334 651
rect 338 648 390 651
rect 2810 648 4310 651
rect 1410 618 2038 621
rect 350 603 353 607
rect 350 602 354 603
rect 1374 603 1377 607
rect 1374 602 1378 603
rect 2398 603 2401 607
rect 2398 602 2402 603
rect 3422 603 3425 607
rect 3422 602 3426 603
rect 4446 603 4449 607
rect 4446 602 4450 603
rect 3626 568 3958 571
rect 5258 558 5277 561
rect 330 548 1630 551
rect 806 531 809 538
rect 714 528 809 531
rect 898 528 1030 531
rect 5267 528 5270 531
rect 862 503 865 507
rect 862 502 866 503
rect 1878 503 1881 507
rect 1878 502 1882 503
rect 2910 503 2913 507
rect 2910 502 2914 503
rect 3934 503 3937 507
rect 3934 502 3938 503
rect 4958 503 4961 507
rect 4958 502 4962 503
rect 2362 468 3214 471
rect 3554 468 3766 471
rect 4866 468 5070 471
rect 562 458 2326 461
rect 3658 458 3678 461
rect 4946 458 5062 461
rect 350 403 353 407
rect 350 402 354 403
rect 1374 403 1377 407
rect 1374 402 1378 403
rect 2398 403 2401 407
rect 2398 402 2402 403
rect 3422 403 3425 407
rect 3422 402 3426 403
rect 4446 403 4449 407
rect 4446 402 4450 403
rect 66 358 2478 361
rect 1906 348 2070 351
rect 338 338 1134 341
rect 1426 338 1526 341
rect 3114 338 3606 341
rect 1154 328 2398 331
rect 2402 328 3366 331
rect 2474 318 3478 321
rect 862 303 865 307
rect 862 302 866 303
rect 1878 303 1881 307
rect 1878 302 1882 303
rect 2910 303 2913 307
rect 2910 302 2914 303
rect 3934 303 3937 307
rect 3934 302 3938 303
rect 4958 303 4961 307
rect 4958 302 4962 303
rect 1242 298 1318 301
rect 3738 288 4222 291
rect 2770 278 3286 281
rect 3802 278 4334 281
rect 1098 268 1318 271
rect 1554 268 1590 271
rect 3242 258 3374 261
rect 3082 238 3166 241
rect 1978 218 3438 221
rect 350 203 353 207
rect 350 202 354 203
rect 1374 203 1377 207
rect 1374 202 1378 203
rect 2398 203 2401 207
rect 2398 202 2402 203
rect 3422 203 3425 207
rect 3422 202 3426 203
rect 4446 203 4449 207
rect 4446 202 4450 203
rect 1402 188 1990 191
rect 2306 178 4102 181
rect 2450 168 3590 171
rect 2858 158 2958 161
rect 490 148 654 151
rect 1658 148 1798 151
rect 2482 148 3150 151
rect 538 138 606 141
rect 1586 138 1694 141
rect 2738 138 2862 141
rect 2866 138 2982 141
rect 1450 128 1862 131
rect 2138 128 2166 131
rect 2538 128 3078 131
rect 3346 128 3390 131
rect 2386 118 3270 121
rect 3354 108 3622 111
rect 862 103 865 107
rect 862 102 866 103
rect 1878 103 1881 107
rect 1878 102 1882 103
rect 2910 103 2913 107
rect 2910 102 2914 103
rect 3934 103 3937 107
rect 3934 102 3938 103
rect 4958 103 4961 107
rect 4958 102 4962 103
rect 522 78 542 81
rect 1138 78 2094 81
rect 2786 78 2814 81
rect 2834 78 2942 81
rect 3350 81 3353 88
rect 3350 78 3574 81
rect 5302 81 5305 88
rect 5299 78 5305 81
rect 538 68 950 71
rect 970 68 1046 71
rect 1482 68 1894 71
rect 2506 68 3150 71
rect 3362 68 3606 71
rect 746 58 990 61
rect 1226 58 1446 61
rect 1450 58 2446 61
rect 3418 58 3646 61
rect 350 3 353 7
rect 350 2 354 3
rect 1374 3 1377 7
rect 1374 2 1378 3
rect 2398 3 2401 7
rect 2398 2 2402 3
rect 3422 3 3425 7
rect 3422 2 3426 3
rect 4446 3 4449 7
rect 4446 2 4450 3
<< m6contact >>
rect 856 3707 862 3708
rect 866 3707 872 3708
rect 856 3703 858 3707
rect 858 3703 862 3707
rect 866 3703 869 3707
rect 869 3703 872 3707
rect 856 3702 862 3703
rect 866 3702 872 3703
rect 1872 3707 1878 3708
rect 1882 3707 1888 3708
rect 1872 3703 1874 3707
rect 1874 3703 1878 3707
rect 1882 3703 1885 3707
rect 1885 3703 1888 3707
rect 1872 3702 1878 3703
rect 1882 3702 1888 3703
rect 2904 3707 2910 3708
rect 2914 3707 2920 3708
rect 2904 3703 2906 3707
rect 2906 3703 2910 3707
rect 2914 3703 2917 3707
rect 2917 3703 2920 3707
rect 2904 3702 2910 3703
rect 2914 3702 2920 3703
rect 3928 3707 3934 3708
rect 3938 3707 3944 3708
rect 3928 3703 3930 3707
rect 3930 3703 3934 3707
rect 3938 3703 3941 3707
rect 3941 3703 3944 3707
rect 3928 3702 3934 3703
rect 3938 3702 3944 3703
rect 4952 3707 4958 3708
rect 4962 3707 4968 3708
rect 4952 3703 4954 3707
rect 4954 3703 4958 3707
rect 4962 3703 4965 3707
rect 4965 3703 4968 3707
rect 4952 3702 4958 3703
rect 4962 3702 4968 3703
rect 344 3607 350 3608
rect 354 3607 360 3608
rect 344 3603 346 3607
rect 346 3603 350 3607
rect 354 3603 357 3607
rect 357 3603 360 3607
rect 344 3602 350 3603
rect 354 3602 360 3603
rect 1368 3607 1374 3608
rect 1378 3607 1384 3608
rect 1368 3603 1370 3607
rect 1370 3603 1374 3607
rect 1378 3603 1381 3607
rect 1381 3603 1384 3607
rect 1368 3602 1374 3603
rect 1378 3602 1384 3603
rect 2392 3607 2398 3608
rect 2402 3607 2408 3608
rect 2392 3603 2394 3607
rect 2394 3603 2398 3607
rect 2402 3603 2405 3607
rect 2405 3603 2408 3607
rect 2392 3602 2398 3603
rect 2402 3602 2408 3603
rect 3416 3607 3422 3608
rect 3426 3607 3432 3608
rect 3416 3603 3418 3607
rect 3418 3603 3422 3607
rect 3426 3603 3429 3607
rect 3429 3603 3432 3607
rect 3416 3602 3422 3603
rect 3426 3602 3432 3603
rect 4440 3607 4446 3608
rect 4450 3607 4456 3608
rect 4440 3603 4442 3607
rect 4442 3603 4446 3607
rect 4450 3603 4453 3607
rect 4453 3603 4456 3607
rect 4440 3602 4446 3603
rect 4450 3602 4456 3603
rect 5229 3547 5235 3553
rect 856 3507 862 3508
rect 866 3507 872 3508
rect 856 3503 858 3507
rect 858 3503 862 3507
rect 866 3503 869 3507
rect 869 3503 872 3507
rect 856 3502 862 3503
rect 866 3502 872 3503
rect 1872 3507 1878 3508
rect 1882 3507 1888 3508
rect 1872 3503 1874 3507
rect 1874 3503 1878 3507
rect 1882 3503 1885 3507
rect 1885 3503 1888 3507
rect 1872 3502 1878 3503
rect 1882 3502 1888 3503
rect 2904 3507 2910 3508
rect 2914 3507 2920 3508
rect 2904 3503 2906 3507
rect 2906 3503 2910 3507
rect 2914 3503 2917 3507
rect 2917 3503 2920 3507
rect 2904 3502 2910 3503
rect 2914 3502 2920 3503
rect 3928 3507 3934 3508
rect 3938 3507 3944 3508
rect 3928 3503 3930 3507
rect 3930 3503 3934 3507
rect 3938 3503 3941 3507
rect 3941 3503 3944 3507
rect 3928 3502 3934 3503
rect 3938 3502 3944 3503
rect 4952 3507 4958 3508
rect 4962 3507 4968 3508
rect 4952 3503 4954 3507
rect 4954 3503 4958 3507
rect 4962 3503 4965 3507
rect 4965 3503 4968 3507
rect 4952 3502 4958 3503
rect 4962 3502 4968 3503
rect 5261 3457 5267 3463
rect 5277 3437 5283 3443
rect 344 3407 350 3408
rect 354 3407 360 3408
rect 344 3403 346 3407
rect 346 3403 350 3407
rect 354 3403 357 3407
rect 357 3403 360 3407
rect 344 3402 350 3403
rect 354 3402 360 3403
rect 1368 3407 1374 3408
rect 1378 3407 1384 3408
rect 1368 3403 1370 3407
rect 1370 3403 1374 3407
rect 1378 3403 1381 3407
rect 1381 3403 1384 3407
rect 1368 3402 1374 3403
rect 1378 3402 1384 3403
rect 2392 3407 2398 3408
rect 2402 3407 2408 3408
rect 2392 3403 2394 3407
rect 2394 3403 2398 3407
rect 2402 3403 2405 3407
rect 2405 3403 2408 3407
rect 2392 3402 2398 3403
rect 2402 3402 2408 3403
rect 3416 3407 3422 3408
rect 3426 3407 3432 3408
rect 3416 3403 3418 3407
rect 3418 3403 3422 3407
rect 3426 3403 3429 3407
rect 3429 3403 3432 3407
rect 3416 3402 3422 3403
rect 3426 3402 3432 3403
rect 4440 3407 4446 3408
rect 4450 3407 4456 3408
rect 4440 3403 4442 3407
rect 4442 3403 4446 3407
rect 4450 3403 4453 3407
rect 4453 3403 4456 3407
rect 4440 3402 4446 3403
rect 4450 3402 4456 3403
rect 856 3307 862 3308
rect 866 3307 872 3308
rect 856 3303 858 3307
rect 858 3303 862 3307
rect 866 3303 869 3307
rect 869 3303 872 3307
rect 856 3302 862 3303
rect 866 3302 872 3303
rect 1872 3307 1878 3308
rect 1882 3307 1888 3308
rect 1872 3303 1874 3307
rect 1874 3303 1878 3307
rect 1882 3303 1885 3307
rect 1885 3303 1888 3307
rect 1872 3302 1878 3303
rect 1882 3302 1888 3303
rect 2904 3307 2910 3308
rect 2914 3307 2920 3308
rect 2904 3303 2906 3307
rect 2906 3303 2910 3307
rect 2914 3303 2917 3307
rect 2917 3303 2920 3307
rect 2904 3302 2910 3303
rect 2914 3302 2920 3303
rect 3928 3307 3934 3308
rect 3938 3307 3944 3308
rect 3928 3303 3930 3307
rect 3930 3303 3934 3307
rect 3938 3303 3941 3307
rect 3941 3303 3944 3307
rect 3928 3302 3934 3303
rect 3938 3302 3944 3303
rect 4952 3307 4958 3308
rect 4962 3307 4968 3308
rect 4952 3303 4954 3307
rect 4954 3303 4958 3307
rect 4962 3303 4965 3307
rect 4965 3303 4968 3307
rect 4952 3302 4958 3303
rect 4962 3302 4968 3303
rect 344 3207 350 3208
rect 354 3207 360 3208
rect 344 3203 346 3207
rect 346 3203 350 3207
rect 354 3203 357 3207
rect 357 3203 360 3207
rect 344 3202 350 3203
rect 354 3202 360 3203
rect 1368 3207 1374 3208
rect 1378 3207 1384 3208
rect 1368 3203 1370 3207
rect 1370 3203 1374 3207
rect 1378 3203 1381 3207
rect 1381 3203 1384 3207
rect 1368 3202 1374 3203
rect 1378 3202 1384 3203
rect 2392 3207 2398 3208
rect 2402 3207 2408 3208
rect 2392 3203 2394 3207
rect 2394 3203 2398 3207
rect 2402 3203 2405 3207
rect 2405 3203 2408 3207
rect 2392 3202 2398 3203
rect 2402 3202 2408 3203
rect 3416 3207 3422 3208
rect 3426 3207 3432 3208
rect 3416 3203 3418 3207
rect 3418 3203 3422 3207
rect 3426 3203 3429 3207
rect 3429 3203 3432 3207
rect 3416 3202 3422 3203
rect 3426 3202 3432 3203
rect 4440 3207 4446 3208
rect 4450 3207 4456 3208
rect 4440 3203 4442 3207
rect 4442 3203 4446 3207
rect 4450 3203 4453 3207
rect 4453 3203 4456 3207
rect 4440 3202 4446 3203
rect 4450 3202 4456 3203
rect 5245 3167 5251 3173
rect 856 3107 862 3108
rect 866 3107 872 3108
rect 856 3103 858 3107
rect 858 3103 862 3107
rect 866 3103 869 3107
rect 869 3103 872 3107
rect 856 3102 862 3103
rect 866 3102 872 3103
rect 1872 3107 1878 3108
rect 1882 3107 1888 3108
rect 1872 3103 1874 3107
rect 1874 3103 1878 3107
rect 1882 3103 1885 3107
rect 1885 3103 1888 3107
rect 1872 3102 1878 3103
rect 1882 3102 1888 3103
rect 2904 3107 2910 3108
rect 2914 3107 2920 3108
rect 2904 3103 2906 3107
rect 2906 3103 2910 3107
rect 2914 3103 2917 3107
rect 2917 3103 2920 3107
rect 2904 3102 2910 3103
rect 2914 3102 2920 3103
rect 3928 3107 3934 3108
rect 3938 3107 3944 3108
rect 3928 3103 3930 3107
rect 3930 3103 3934 3107
rect 3938 3103 3941 3107
rect 3941 3103 3944 3107
rect 3928 3102 3934 3103
rect 3938 3102 3944 3103
rect 4952 3107 4958 3108
rect 4962 3107 4968 3108
rect 4952 3103 4954 3107
rect 4954 3103 4958 3107
rect 4962 3103 4965 3107
rect 4965 3103 4968 3107
rect 4952 3102 4958 3103
rect 4962 3102 4968 3103
rect 5293 3067 5299 3073
rect 5309 3067 5315 3073
rect 5277 3057 5283 3063
rect 344 3007 350 3008
rect 354 3007 360 3008
rect 344 3003 346 3007
rect 346 3003 350 3007
rect 354 3003 357 3007
rect 357 3003 360 3007
rect 344 3002 350 3003
rect 354 3002 360 3003
rect 1368 3007 1374 3008
rect 1378 3007 1384 3008
rect 1368 3003 1370 3007
rect 1370 3003 1374 3007
rect 1378 3003 1381 3007
rect 1381 3003 1384 3007
rect 1368 3002 1374 3003
rect 1378 3002 1384 3003
rect 2392 3007 2398 3008
rect 2402 3007 2408 3008
rect 2392 3003 2394 3007
rect 2394 3003 2398 3007
rect 2402 3003 2405 3007
rect 2405 3003 2408 3007
rect 2392 3002 2398 3003
rect 2402 3002 2408 3003
rect 3416 3007 3422 3008
rect 3426 3007 3432 3008
rect 3416 3003 3418 3007
rect 3418 3003 3422 3007
rect 3426 3003 3429 3007
rect 3429 3003 3432 3007
rect 3416 3002 3422 3003
rect 3426 3002 3432 3003
rect 4440 3007 4446 3008
rect 4450 3007 4456 3008
rect 4440 3003 4442 3007
rect 4442 3003 4446 3007
rect 4450 3003 4453 3007
rect 4453 3003 4456 3007
rect 4440 3002 4446 3003
rect 4450 3002 4456 3003
rect 5277 2987 5283 2993
rect 856 2907 862 2908
rect 866 2907 872 2908
rect 856 2903 858 2907
rect 858 2903 862 2907
rect 866 2903 869 2907
rect 869 2903 872 2907
rect 856 2902 862 2903
rect 866 2902 872 2903
rect 1872 2907 1878 2908
rect 1882 2907 1888 2908
rect 1872 2903 1874 2907
rect 1874 2903 1878 2907
rect 1882 2903 1885 2907
rect 1885 2903 1888 2907
rect 1872 2902 1878 2903
rect 1882 2902 1888 2903
rect 2904 2907 2910 2908
rect 2914 2907 2920 2908
rect 2904 2903 2906 2907
rect 2906 2903 2910 2907
rect 2914 2903 2917 2907
rect 2917 2903 2920 2907
rect 2904 2902 2910 2903
rect 2914 2902 2920 2903
rect 3928 2907 3934 2908
rect 3938 2907 3944 2908
rect 3928 2903 3930 2907
rect 3930 2903 3934 2907
rect 3938 2903 3941 2907
rect 3941 2903 3944 2907
rect 3928 2902 3934 2903
rect 3938 2902 3944 2903
rect 4952 2907 4958 2908
rect 4962 2907 4968 2908
rect 4952 2903 4954 2907
rect 4954 2903 4958 2907
rect 4962 2903 4965 2907
rect 4965 2903 4968 2907
rect 4952 2902 4958 2903
rect 4962 2902 4968 2903
rect 344 2807 350 2808
rect 354 2807 360 2808
rect 344 2803 346 2807
rect 346 2803 350 2807
rect 354 2803 357 2807
rect 357 2803 360 2807
rect 344 2802 350 2803
rect 354 2802 360 2803
rect 1368 2807 1374 2808
rect 1378 2807 1384 2808
rect 1368 2803 1370 2807
rect 1370 2803 1374 2807
rect 1378 2803 1381 2807
rect 1381 2803 1384 2807
rect 1368 2802 1374 2803
rect 1378 2802 1384 2803
rect 2392 2807 2398 2808
rect 2402 2807 2408 2808
rect 2392 2803 2394 2807
rect 2394 2803 2398 2807
rect 2402 2803 2405 2807
rect 2405 2803 2408 2807
rect 2392 2802 2398 2803
rect 2402 2802 2408 2803
rect 3416 2807 3422 2808
rect 3426 2807 3432 2808
rect 3416 2803 3418 2807
rect 3418 2803 3422 2807
rect 3426 2803 3429 2807
rect 3429 2803 3432 2807
rect 3416 2802 3422 2803
rect 3426 2802 3432 2803
rect 4440 2807 4446 2808
rect 4450 2807 4456 2808
rect 4440 2803 4442 2807
rect 4442 2803 4446 2807
rect 4450 2803 4453 2807
rect 4453 2803 4456 2807
rect 4440 2802 4446 2803
rect 4450 2802 4456 2803
rect 856 2707 862 2708
rect 866 2707 872 2708
rect 856 2703 858 2707
rect 858 2703 862 2707
rect 866 2703 869 2707
rect 869 2703 872 2707
rect 856 2702 862 2703
rect 866 2702 872 2703
rect 1872 2707 1878 2708
rect 1882 2707 1888 2708
rect 1872 2703 1874 2707
rect 1874 2703 1878 2707
rect 1882 2703 1885 2707
rect 1885 2703 1888 2707
rect 1872 2702 1878 2703
rect 1882 2702 1888 2703
rect 2904 2707 2910 2708
rect 2914 2707 2920 2708
rect 2904 2703 2906 2707
rect 2906 2703 2910 2707
rect 2914 2703 2917 2707
rect 2917 2703 2920 2707
rect 2904 2702 2910 2703
rect 2914 2702 2920 2703
rect 3928 2707 3934 2708
rect 3938 2707 3944 2708
rect 3928 2703 3930 2707
rect 3930 2703 3934 2707
rect 3938 2703 3941 2707
rect 3941 2703 3944 2707
rect 3928 2702 3934 2703
rect 3938 2702 3944 2703
rect 4952 2707 4958 2708
rect 4962 2707 4968 2708
rect 4952 2703 4954 2707
rect 4954 2703 4958 2707
rect 4962 2703 4965 2707
rect 4965 2703 4968 2707
rect 4952 2702 4958 2703
rect 4962 2702 4968 2703
rect 5293 2677 5299 2683
rect 5277 2637 5283 2643
rect 5277 2627 5283 2633
rect 344 2607 350 2608
rect 354 2607 360 2608
rect 344 2603 346 2607
rect 346 2603 350 2607
rect 354 2603 357 2607
rect 357 2603 360 2607
rect 344 2602 350 2603
rect 354 2602 360 2603
rect 1368 2607 1374 2608
rect 1378 2607 1384 2608
rect 1368 2603 1370 2607
rect 1370 2603 1374 2607
rect 1378 2603 1381 2607
rect 1381 2603 1384 2607
rect 1368 2602 1374 2603
rect 1378 2602 1384 2603
rect 2392 2607 2398 2608
rect 2402 2607 2408 2608
rect 2392 2603 2394 2607
rect 2394 2603 2398 2607
rect 2402 2603 2405 2607
rect 2405 2603 2408 2607
rect 2392 2602 2398 2603
rect 2402 2602 2408 2603
rect 3416 2607 3422 2608
rect 3426 2607 3432 2608
rect 3416 2603 3418 2607
rect 3418 2603 3422 2607
rect 3426 2603 3429 2607
rect 3429 2603 3432 2607
rect 3416 2602 3422 2603
rect 3426 2602 3432 2603
rect 4440 2607 4446 2608
rect 4450 2607 4456 2608
rect 4440 2603 4442 2607
rect 4442 2603 4446 2607
rect 4450 2603 4453 2607
rect 4453 2603 4456 2607
rect 4440 2602 4446 2603
rect 4450 2602 4456 2603
rect 5309 2577 5315 2583
rect 5309 2567 5315 2573
rect 5357 2517 5363 2523
rect 856 2507 862 2508
rect 866 2507 872 2508
rect 856 2503 858 2507
rect 858 2503 862 2507
rect 866 2503 869 2507
rect 869 2503 872 2507
rect 856 2502 862 2503
rect 866 2502 872 2503
rect 1872 2507 1878 2508
rect 1882 2507 1888 2508
rect 1872 2503 1874 2507
rect 1874 2503 1878 2507
rect 1882 2503 1885 2507
rect 1885 2503 1888 2507
rect 1872 2502 1878 2503
rect 1882 2502 1888 2503
rect 2904 2507 2910 2508
rect 2914 2507 2920 2508
rect 2904 2503 2906 2507
rect 2906 2503 2910 2507
rect 2914 2503 2917 2507
rect 2917 2503 2920 2507
rect 2904 2502 2910 2503
rect 2914 2502 2920 2503
rect 3928 2507 3934 2508
rect 3938 2507 3944 2508
rect 3928 2503 3930 2507
rect 3930 2503 3934 2507
rect 3938 2503 3941 2507
rect 3941 2503 3944 2507
rect 3928 2502 3934 2503
rect 3938 2502 3944 2503
rect 4952 2507 4958 2508
rect 4962 2507 4968 2508
rect 4952 2503 4954 2507
rect 4954 2503 4958 2507
rect 4962 2503 4965 2507
rect 4965 2503 4968 2507
rect 4952 2502 4958 2503
rect 4962 2502 4968 2503
rect 2141 2467 2147 2473
rect 2621 2437 2627 2443
rect 344 2407 350 2408
rect 354 2407 360 2408
rect 344 2403 346 2407
rect 346 2403 350 2407
rect 354 2403 357 2407
rect 357 2403 360 2407
rect 344 2402 350 2403
rect 354 2402 360 2403
rect 1368 2407 1374 2408
rect 1378 2407 1384 2408
rect 1368 2403 1370 2407
rect 1370 2403 1374 2407
rect 1378 2403 1381 2407
rect 1381 2403 1384 2407
rect 1368 2402 1374 2403
rect 1378 2402 1384 2403
rect 2392 2407 2398 2408
rect 2402 2407 2408 2408
rect 2392 2403 2394 2407
rect 2394 2403 2398 2407
rect 2402 2403 2405 2407
rect 2405 2403 2408 2407
rect 2392 2402 2398 2403
rect 2402 2402 2408 2403
rect 3416 2407 3422 2408
rect 3426 2407 3432 2408
rect 3416 2403 3418 2407
rect 3418 2403 3422 2407
rect 3426 2403 3429 2407
rect 3429 2403 3432 2407
rect 3416 2402 3422 2403
rect 3426 2402 3432 2403
rect 4440 2407 4446 2408
rect 4450 2407 4456 2408
rect 5213 2407 5219 2413
rect 4440 2403 4442 2407
rect 4442 2403 4446 2407
rect 4450 2403 4453 2407
rect 4453 2403 4456 2407
rect 4440 2402 4446 2403
rect 4450 2402 4456 2403
rect 856 2307 862 2308
rect 866 2307 872 2308
rect 856 2303 858 2307
rect 858 2303 862 2307
rect 866 2303 869 2307
rect 869 2303 872 2307
rect 856 2302 862 2303
rect 866 2302 872 2303
rect 1872 2307 1878 2308
rect 1882 2307 1888 2308
rect 1872 2303 1874 2307
rect 1874 2303 1878 2307
rect 1882 2303 1885 2307
rect 1885 2303 1888 2307
rect 1872 2302 1878 2303
rect 1882 2302 1888 2303
rect 2904 2307 2910 2308
rect 2914 2307 2920 2308
rect 2904 2303 2906 2307
rect 2906 2303 2910 2307
rect 2914 2303 2917 2307
rect 2917 2303 2920 2307
rect 2904 2302 2910 2303
rect 2914 2302 2920 2303
rect 3928 2307 3934 2308
rect 3938 2307 3944 2308
rect 3928 2303 3930 2307
rect 3930 2303 3934 2307
rect 3938 2303 3941 2307
rect 3941 2303 3944 2307
rect 3928 2302 3934 2303
rect 3938 2302 3944 2303
rect 4952 2307 4958 2308
rect 4962 2307 4968 2308
rect 4952 2303 4954 2307
rect 4954 2303 4958 2307
rect 4962 2303 4965 2307
rect 4965 2303 4968 2307
rect 4952 2302 4958 2303
rect 4962 2302 4968 2303
rect 344 2207 350 2208
rect 354 2207 360 2208
rect 344 2203 346 2207
rect 346 2203 350 2207
rect 354 2203 357 2207
rect 357 2203 360 2207
rect 344 2202 350 2203
rect 354 2202 360 2203
rect 1368 2207 1374 2208
rect 1378 2207 1384 2208
rect 1368 2203 1370 2207
rect 1370 2203 1374 2207
rect 1378 2203 1381 2207
rect 1381 2203 1384 2207
rect 1368 2202 1374 2203
rect 1378 2202 1384 2203
rect 2392 2207 2398 2208
rect 2402 2207 2408 2208
rect 2392 2203 2394 2207
rect 2394 2203 2398 2207
rect 2402 2203 2405 2207
rect 2405 2203 2408 2207
rect 2392 2202 2398 2203
rect 2402 2202 2408 2203
rect 3416 2207 3422 2208
rect 3426 2207 3432 2208
rect 3416 2203 3418 2207
rect 3418 2203 3422 2207
rect 3426 2203 3429 2207
rect 3429 2203 3432 2207
rect 3416 2202 3422 2203
rect 3426 2202 3432 2203
rect 4440 2207 4446 2208
rect 4450 2207 4456 2208
rect 4440 2203 4442 2207
rect 4442 2203 4446 2207
rect 4450 2203 4453 2207
rect 4453 2203 4456 2207
rect 4440 2202 4446 2203
rect 4450 2202 4456 2203
rect 5213 2167 5219 2173
rect 5213 2147 5219 2153
rect 5277 2137 5283 2143
rect 5229 2127 5235 2133
rect 5277 2127 5283 2133
rect 856 2107 862 2108
rect 866 2107 872 2108
rect 856 2103 858 2107
rect 858 2103 862 2107
rect 866 2103 869 2107
rect 869 2103 872 2107
rect 856 2102 862 2103
rect 866 2102 872 2103
rect 1872 2107 1878 2108
rect 1882 2107 1888 2108
rect 1872 2103 1874 2107
rect 1874 2103 1878 2107
rect 1882 2103 1885 2107
rect 1885 2103 1888 2107
rect 1872 2102 1878 2103
rect 1882 2102 1888 2103
rect 2904 2107 2910 2108
rect 2914 2107 2920 2108
rect 2904 2103 2906 2107
rect 2906 2103 2910 2107
rect 2914 2103 2917 2107
rect 2917 2103 2920 2107
rect 2904 2102 2910 2103
rect 2914 2102 2920 2103
rect 3928 2107 3934 2108
rect 3938 2107 3944 2108
rect 3928 2103 3930 2107
rect 3930 2103 3934 2107
rect 3938 2103 3941 2107
rect 3941 2103 3944 2107
rect 3928 2102 3934 2103
rect 3938 2102 3944 2103
rect 4952 2107 4958 2108
rect 4962 2107 4968 2108
rect 5229 2107 5235 2113
rect 4952 2103 4954 2107
rect 4954 2103 4958 2107
rect 4962 2103 4965 2107
rect 4965 2103 4968 2107
rect 4952 2102 4958 2103
rect 4962 2102 4968 2103
rect 5277 2097 5283 2103
rect 2621 2037 2627 2043
rect 344 2007 350 2008
rect 354 2007 360 2008
rect 344 2003 346 2007
rect 346 2003 350 2007
rect 354 2003 357 2007
rect 357 2003 360 2007
rect 344 2002 350 2003
rect 354 2002 360 2003
rect 1368 2007 1374 2008
rect 1378 2007 1384 2008
rect 1368 2003 1370 2007
rect 1370 2003 1374 2007
rect 1378 2003 1381 2007
rect 1381 2003 1384 2007
rect 1368 2002 1374 2003
rect 1378 2002 1384 2003
rect 2392 2007 2398 2008
rect 2402 2007 2408 2008
rect 2392 2003 2394 2007
rect 2394 2003 2398 2007
rect 2402 2003 2405 2007
rect 2405 2003 2408 2007
rect 2392 2002 2398 2003
rect 2402 2002 2408 2003
rect 3416 2007 3422 2008
rect 3426 2007 3432 2008
rect 3416 2003 3418 2007
rect 3418 2003 3422 2007
rect 3426 2003 3429 2007
rect 3429 2003 3432 2007
rect 3416 2002 3422 2003
rect 3426 2002 3432 2003
rect 4440 2007 4446 2008
rect 4450 2007 4456 2008
rect 4440 2003 4442 2007
rect 4442 2003 4446 2007
rect 4450 2003 4453 2007
rect 4453 2003 4456 2007
rect 4440 2002 4446 2003
rect 4450 2002 4456 2003
rect 856 1907 862 1908
rect 866 1907 872 1908
rect 856 1903 858 1907
rect 858 1903 862 1907
rect 866 1903 869 1907
rect 869 1903 872 1907
rect 856 1902 862 1903
rect 866 1902 872 1903
rect 1872 1907 1878 1908
rect 1882 1907 1888 1908
rect 1872 1903 1874 1907
rect 1874 1903 1878 1907
rect 1882 1903 1885 1907
rect 1885 1903 1888 1907
rect 1872 1902 1878 1903
rect 1882 1902 1888 1903
rect 2904 1907 2910 1908
rect 2914 1907 2920 1908
rect 2904 1903 2906 1907
rect 2906 1903 2910 1907
rect 2914 1903 2917 1907
rect 2917 1903 2920 1907
rect 2904 1902 2910 1903
rect 2914 1902 2920 1903
rect 3928 1907 3934 1908
rect 3938 1907 3944 1908
rect 3928 1903 3930 1907
rect 3930 1903 3934 1907
rect 3938 1903 3941 1907
rect 3941 1903 3944 1907
rect 3928 1902 3934 1903
rect 3938 1902 3944 1903
rect 4952 1907 4958 1908
rect 4962 1907 4968 1908
rect 4952 1903 4954 1907
rect 4954 1903 4958 1907
rect 4962 1903 4965 1907
rect 4965 1903 4968 1907
rect 4952 1902 4958 1903
rect 4962 1902 4968 1903
rect 344 1807 350 1808
rect 354 1807 360 1808
rect 344 1803 346 1807
rect 346 1803 350 1807
rect 354 1803 357 1807
rect 357 1803 360 1807
rect 344 1802 350 1803
rect 354 1802 360 1803
rect 1368 1807 1374 1808
rect 1378 1807 1384 1808
rect 1368 1803 1370 1807
rect 1370 1803 1374 1807
rect 1378 1803 1381 1807
rect 1381 1803 1384 1807
rect 1368 1802 1374 1803
rect 1378 1802 1384 1803
rect 2392 1807 2398 1808
rect 2402 1807 2408 1808
rect 2392 1803 2394 1807
rect 2394 1803 2398 1807
rect 2402 1803 2405 1807
rect 2405 1803 2408 1807
rect 2392 1802 2398 1803
rect 2402 1802 2408 1803
rect 3416 1807 3422 1808
rect 3426 1807 3432 1808
rect 3416 1803 3418 1807
rect 3418 1803 3422 1807
rect 3426 1803 3429 1807
rect 3429 1803 3432 1807
rect 3416 1802 3422 1803
rect 3426 1802 3432 1803
rect 4440 1807 4446 1808
rect 4450 1807 4456 1808
rect 4440 1803 4442 1807
rect 4442 1803 4446 1807
rect 4450 1803 4453 1807
rect 4453 1803 4456 1807
rect 4440 1802 4446 1803
rect 4450 1802 4456 1803
rect 856 1707 862 1708
rect 866 1707 872 1708
rect 856 1703 858 1707
rect 858 1703 862 1707
rect 866 1703 869 1707
rect 869 1703 872 1707
rect 856 1702 862 1703
rect 866 1702 872 1703
rect 1872 1707 1878 1708
rect 1882 1707 1888 1708
rect 1872 1703 1874 1707
rect 1874 1703 1878 1707
rect 1882 1703 1885 1707
rect 1885 1703 1888 1707
rect 1872 1702 1878 1703
rect 1882 1702 1888 1703
rect 2904 1707 2910 1708
rect 2914 1707 2920 1708
rect 2904 1703 2906 1707
rect 2906 1703 2910 1707
rect 2914 1703 2917 1707
rect 2917 1703 2920 1707
rect 2904 1702 2910 1703
rect 2914 1702 2920 1703
rect 3928 1707 3934 1708
rect 3938 1707 3944 1708
rect 3928 1703 3930 1707
rect 3930 1703 3934 1707
rect 3938 1703 3941 1707
rect 3941 1703 3944 1707
rect 3928 1702 3934 1703
rect 3938 1702 3944 1703
rect 4952 1707 4958 1708
rect 4962 1707 4968 1708
rect 4952 1703 4954 1707
rect 4954 1703 4958 1707
rect 4962 1703 4965 1707
rect 4965 1703 4968 1707
rect 4952 1702 4958 1703
rect 4962 1702 4968 1703
rect 5229 1677 5235 1683
rect 344 1607 350 1608
rect 354 1607 360 1608
rect 344 1603 346 1607
rect 346 1603 350 1607
rect 354 1603 357 1607
rect 357 1603 360 1607
rect 344 1602 350 1603
rect 354 1602 360 1603
rect 1368 1607 1374 1608
rect 1378 1607 1384 1608
rect 1368 1603 1370 1607
rect 1370 1603 1374 1607
rect 1378 1603 1381 1607
rect 1381 1603 1384 1607
rect 1368 1602 1374 1603
rect 1378 1602 1384 1603
rect 2392 1607 2398 1608
rect 2402 1607 2408 1608
rect 2392 1603 2394 1607
rect 2394 1603 2398 1607
rect 2402 1603 2405 1607
rect 2405 1603 2408 1607
rect 2392 1602 2398 1603
rect 2402 1602 2408 1603
rect 3416 1607 3422 1608
rect 3426 1607 3432 1608
rect 3416 1603 3418 1607
rect 3418 1603 3422 1607
rect 3426 1603 3429 1607
rect 3429 1603 3432 1607
rect 3416 1602 3422 1603
rect 3426 1602 3432 1603
rect 4440 1607 4446 1608
rect 4450 1607 4456 1608
rect 4440 1603 4442 1607
rect 4442 1603 4446 1607
rect 4450 1603 4453 1607
rect 4453 1603 4456 1607
rect 4440 1602 4446 1603
rect 4450 1602 4456 1603
rect 856 1507 862 1508
rect 866 1507 872 1508
rect 856 1503 858 1507
rect 858 1503 862 1507
rect 866 1503 869 1507
rect 869 1503 872 1507
rect 856 1502 862 1503
rect 866 1502 872 1503
rect 1872 1507 1878 1508
rect 1882 1507 1888 1508
rect 1872 1503 1874 1507
rect 1874 1503 1878 1507
rect 1882 1503 1885 1507
rect 1885 1503 1888 1507
rect 1872 1502 1878 1503
rect 1882 1502 1888 1503
rect 2904 1507 2910 1508
rect 2914 1507 2920 1508
rect 2904 1503 2906 1507
rect 2906 1503 2910 1507
rect 2914 1503 2917 1507
rect 2917 1503 2920 1507
rect 2904 1502 2910 1503
rect 2914 1502 2920 1503
rect 3928 1507 3934 1508
rect 3938 1507 3944 1508
rect 3928 1503 3930 1507
rect 3930 1503 3934 1507
rect 3938 1503 3941 1507
rect 3941 1503 3944 1507
rect 3928 1502 3934 1503
rect 3938 1502 3944 1503
rect 4952 1507 4958 1508
rect 4962 1507 4968 1508
rect 4952 1503 4954 1507
rect 4954 1503 4958 1507
rect 4962 1503 4965 1507
rect 4965 1503 4968 1507
rect 4952 1502 4958 1503
rect 4962 1502 4968 1503
rect 344 1407 350 1408
rect 354 1407 360 1408
rect 344 1403 346 1407
rect 346 1403 350 1407
rect 354 1403 357 1407
rect 357 1403 360 1407
rect 344 1402 350 1403
rect 354 1402 360 1403
rect 1368 1407 1374 1408
rect 1378 1407 1384 1408
rect 1368 1403 1370 1407
rect 1370 1403 1374 1407
rect 1378 1403 1381 1407
rect 1381 1403 1384 1407
rect 1368 1402 1374 1403
rect 1378 1402 1384 1403
rect 2392 1407 2398 1408
rect 2402 1407 2408 1408
rect 2392 1403 2394 1407
rect 2394 1403 2398 1407
rect 2402 1403 2405 1407
rect 2405 1403 2408 1407
rect 2392 1402 2398 1403
rect 2402 1402 2408 1403
rect 3416 1407 3422 1408
rect 3426 1407 3432 1408
rect 3416 1403 3418 1407
rect 3418 1403 3422 1407
rect 3426 1403 3429 1407
rect 3429 1403 3432 1407
rect 3416 1402 3422 1403
rect 3426 1402 3432 1403
rect 4440 1407 4446 1408
rect 4450 1407 4456 1408
rect 4440 1403 4442 1407
rect 4442 1403 4446 1407
rect 4450 1403 4453 1407
rect 4453 1403 4456 1407
rect 4440 1402 4446 1403
rect 4450 1402 4456 1403
rect 856 1307 862 1308
rect 866 1307 872 1308
rect 856 1303 858 1307
rect 858 1303 862 1307
rect 866 1303 869 1307
rect 869 1303 872 1307
rect 856 1302 862 1303
rect 866 1302 872 1303
rect 1872 1307 1878 1308
rect 1882 1307 1888 1308
rect 1872 1303 1874 1307
rect 1874 1303 1878 1307
rect 1882 1303 1885 1307
rect 1885 1303 1888 1307
rect 1872 1302 1878 1303
rect 1882 1302 1888 1303
rect 2904 1307 2910 1308
rect 2914 1307 2920 1308
rect 2904 1303 2906 1307
rect 2906 1303 2910 1307
rect 2914 1303 2917 1307
rect 2917 1303 2920 1307
rect 2904 1302 2910 1303
rect 2914 1302 2920 1303
rect 3928 1307 3934 1308
rect 3938 1307 3944 1308
rect 3928 1303 3930 1307
rect 3930 1303 3934 1307
rect 3938 1303 3941 1307
rect 3941 1303 3944 1307
rect 3928 1302 3934 1303
rect 3938 1302 3944 1303
rect 4952 1307 4958 1308
rect 4962 1307 4968 1308
rect 4952 1303 4954 1307
rect 4954 1303 4958 1307
rect 4962 1303 4965 1307
rect 4965 1303 4968 1307
rect 4952 1302 4958 1303
rect 4962 1302 4968 1303
rect 5277 1287 5283 1293
rect 5213 1277 5219 1283
rect 2141 1267 2147 1273
rect 344 1207 350 1208
rect 354 1207 360 1208
rect 344 1203 346 1207
rect 346 1203 350 1207
rect 354 1203 357 1207
rect 357 1203 360 1207
rect 344 1202 350 1203
rect 354 1202 360 1203
rect 1368 1207 1374 1208
rect 1378 1207 1384 1208
rect 1368 1203 1370 1207
rect 1370 1203 1374 1207
rect 1378 1203 1381 1207
rect 1381 1203 1384 1207
rect 1368 1202 1374 1203
rect 1378 1202 1384 1203
rect 2392 1207 2398 1208
rect 2402 1207 2408 1208
rect 2392 1203 2394 1207
rect 2394 1203 2398 1207
rect 2402 1203 2405 1207
rect 2405 1203 2408 1207
rect 2392 1202 2398 1203
rect 2402 1202 2408 1203
rect 3416 1207 3422 1208
rect 3426 1207 3432 1208
rect 3416 1203 3418 1207
rect 3418 1203 3422 1207
rect 3426 1203 3429 1207
rect 3429 1203 3432 1207
rect 3416 1202 3422 1203
rect 3426 1202 3432 1203
rect 4440 1207 4446 1208
rect 4450 1207 4456 1208
rect 4440 1203 4442 1207
rect 4442 1203 4446 1207
rect 4450 1203 4453 1207
rect 4453 1203 4456 1207
rect 4440 1202 4446 1203
rect 4450 1202 4456 1203
rect 856 1107 862 1108
rect 866 1107 872 1108
rect 856 1103 858 1107
rect 858 1103 862 1107
rect 866 1103 869 1107
rect 869 1103 872 1107
rect 856 1102 862 1103
rect 866 1102 872 1103
rect 1872 1107 1878 1108
rect 1882 1107 1888 1108
rect 1872 1103 1874 1107
rect 1874 1103 1878 1107
rect 1882 1103 1885 1107
rect 1885 1103 1888 1107
rect 1872 1102 1878 1103
rect 1882 1102 1888 1103
rect 2904 1107 2910 1108
rect 2914 1107 2920 1108
rect 2904 1103 2906 1107
rect 2906 1103 2910 1107
rect 2914 1103 2917 1107
rect 2917 1103 2920 1107
rect 2904 1102 2910 1103
rect 2914 1102 2920 1103
rect 3928 1107 3934 1108
rect 3938 1107 3944 1108
rect 3928 1103 3930 1107
rect 3930 1103 3934 1107
rect 3938 1103 3941 1107
rect 3941 1103 3944 1107
rect 3928 1102 3934 1103
rect 3938 1102 3944 1103
rect 4952 1107 4958 1108
rect 4962 1107 4968 1108
rect 4952 1103 4954 1107
rect 4954 1103 4958 1107
rect 4962 1103 4965 1107
rect 4965 1103 4968 1107
rect 4952 1102 4958 1103
rect 4962 1102 4968 1103
rect 344 1007 350 1008
rect 354 1007 360 1008
rect 344 1003 346 1007
rect 346 1003 350 1007
rect 354 1003 357 1007
rect 357 1003 360 1007
rect 344 1002 350 1003
rect 354 1002 360 1003
rect 1368 1007 1374 1008
rect 1378 1007 1384 1008
rect 1368 1003 1370 1007
rect 1370 1003 1374 1007
rect 1378 1003 1381 1007
rect 1381 1003 1384 1007
rect 1368 1002 1374 1003
rect 1378 1002 1384 1003
rect 2392 1007 2398 1008
rect 2402 1007 2408 1008
rect 2392 1003 2394 1007
rect 2394 1003 2398 1007
rect 2402 1003 2405 1007
rect 2405 1003 2408 1007
rect 2392 1002 2398 1003
rect 2402 1002 2408 1003
rect 3416 1007 3422 1008
rect 3426 1007 3432 1008
rect 3416 1003 3418 1007
rect 3418 1003 3422 1007
rect 3426 1003 3429 1007
rect 3429 1003 3432 1007
rect 3416 1002 3422 1003
rect 3426 1002 3432 1003
rect 4440 1007 4446 1008
rect 4450 1007 4456 1008
rect 4440 1003 4442 1007
rect 4442 1003 4446 1007
rect 4450 1003 4453 1007
rect 4453 1003 4456 1007
rect 4440 1002 4446 1003
rect 4450 1002 4456 1003
rect 856 907 862 908
rect 866 907 872 908
rect 856 903 858 907
rect 858 903 862 907
rect 866 903 869 907
rect 869 903 872 907
rect 856 902 862 903
rect 866 902 872 903
rect 1872 907 1878 908
rect 1882 907 1888 908
rect 1872 903 1874 907
rect 1874 903 1878 907
rect 1882 903 1885 907
rect 1885 903 1888 907
rect 1872 902 1878 903
rect 1882 902 1888 903
rect 2904 907 2910 908
rect 2914 907 2920 908
rect 2904 903 2906 907
rect 2906 903 2910 907
rect 2914 903 2917 907
rect 2917 903 2920 907
rect 2904 902 2910 903
rect 2914 902 2920 903
rect 3928 907 3934 908
rect 3938 907 3944 908
rect 3928 903 3930 907
rect 3930 903 3934 907
rect 3938 903 3941 907
rect 3941 903 3944 907
rect 3928 902 3934 903
rect 3938 902 3944 903
rect 4952 907 4958 908
rect 4962 907 4968 908
rect 4952 903 4954 907
rect 4954 903 4958 907
rect 4962 903 4965 907
rect 4965 903 4968 907
rect 4952 902 4958 903
rect 4962 902 4968 903
rect 5245 867 5251 873
rect 5357 857 5363 863
rect 5309 847 5315 853
rect 344 807 350 808
rect 354 807 360 808
rect 344 803 346 807
rect 346 803 350 807
rect 354 803 357 807
rect 357 803 360 807
rect 344 802 350 803
rect 354 802 360 803
rect 1368 807 1374 808
rect 1378 807 1384 808
rect 1368 803 1370 807
rect 1370 803 1374 807
rect 1378 803 1381 807
rect 1381 803 1384 807
rect 1368 802 1374 803
rect 1378 802 1384 803
rect 2392 807 2398 808
rect 2402 807 2408 808
rect 2392 803 2394 807
rect 2394 803 2398 807
rect 2402 803 2405 807
rect 2405 803 2408 807
rect 2392 802 2398 803
rect 2402 802 2408 803
rect 3416 807 3422 808
rect 3426 807 3432 808
rect 3416 803 3418 807
rect 3418 803 3422 807
rect 3426 803 3429 807
rect 3429 803 3432 807
rect 3416 802 3422 803
rect 3426 802 3432 803
rect 4440 807 4446 808
rect 4450 807 4456 808
rect 4440 803 4442 807
rect 4442 803 4446 807
rect 4450 803 4453 807
rect 4453 803 4456 807
rect 4440 802 4446 803
rect 4450 802 4456 803
rect 856 707 862 708
rect 866 707 872 708
rect 856 703 858 707
rect 858 703 862 707
rect 866 703 869 707
rect 869 703 872 707
rect 856 702 862 703
rect 866 702 872 703
rect 1872 707 1878 708
rect 1882 707 1888 708
rect 1872 703 1874 707
rect 1874 703 1878 707
rect 1882 703 1885 707
rect 1885 703 1888 707
rect 1872 702 1878 703
rect 1882 702 1888 703
rect 2904 707 2910 708
rect 2914 707 2920 708
rect 2904 703 2906 707
rect 2906 703 2910 707
rect 2914 703 2917 707
rect 2917 703 2920 707
rect 2904 702 2910 703
rect 2914 702 2920 703
rect 3928 707 3934 708
rect 3938 707 3944 708
rect 3928 703 3930 707
rect 3930 703 3934 707
rect 3938 703 3941 707
rect 3941 703 3944 707
rect 3928 702 3934 703
rect 3938 702 3944 703
rect 4952 707 4958 708
rect 4962 707 4968 708
rect 4952 703 4954 707
rect 4954 703 4958 707
rect 4962 703 4965 707
rect 4965 703 4968 707
rect 4952 702 4958 703
rect 4962 702 4968 703
rect 344 607 350 608
rect 354 607 360 608
rect 344 603 346 607
rect 346 603 350 607
rect 354 603 357 607
rect 357 603 360 607
rect 344 602 350 603
rect 354 602 360 603
rect 1368 607 1374 608
rect 1378 607 1384 608
rect 1368 603 1370 607
rect 1370 603 1374 607
rect 1378 603 1381 607
rect 1381 603 1384 607
rect 1368 602 1374 603
rect 1378 602 1384 603
rect 2392 607 2398 608
rect 2402 607 2408 608
rect 2392 603 2394 607
rect 2394 603 2398 607
rect 2402 603 2405 607
rect 2405 603 2408 607
rect 2392 602 2398 603
rect 2402 602 2408 603
rect 3416 607 3422 608
rect 3426 607 3432 608
rect 3416 603 3418 607
rect 3418 603 3422 607
rect 3426 603 3429 607
rect 3429 603 3432 607
rect 3416 602 3422 603
rect 3426 602 3432 603
rect 4440 607 4446 608
rect 4450 607 4456 608
rect 4440 603 4442 607
rect 4442 603 4446 607
rect 4450 603 4453 607
rect 4453 603 4456 607
rect 4440 602 4446 603
rect 4450 602 4456 603
rect 5277 557 5283 563
rect 5261 527 5267 533
rect 856 507 862 508
rect 866 507 872 508
rect 856 503 858 507
rect 858 503 862 507
rect 866 503 869 507
rect 869 503 872 507
rect 856 502 862 503
rect 866 502 872 503
rect 1872 507 1878 508
rect 1882 507 1888 508
rect 1872 503 1874 507
rect 1874 503 1878 507
rect 1882 503 1885 507
rect 1885 503 1888 507
rect 1872 502 1878 503
rect 1882 502 1888 503
rect 2904 507 2910 508
rect 2914 507 2920 508
rect 2904 503 2906 507
rect 2906 503 2910 507
rect 2914 503 2917 507
rect 2917 503 2920 507
rect 2904 502 2910 503
rect 2914 502 2920 503
rect 3928 507 3934 508
rect 3938 507 3944 508
rect 3928 503 3930 507
rect 3930 503 3934 507
rect 3938 503 3941 507
rect 3941 503 3944 507
rect 3928 502 3934 503
rect 3938 502 3944 503
rect 4952 507 4958 508
rect 4962 507 4968 508
rect 4952 503 4954 507
rect 4954 503 4958 507
rect 4962 503 4965 507
rect 4965 503 4968 507
rect 4952 502 4958 503
rect 4962 502 4968 503
rect 344 407 350 408
rect 354 407 360 408
rect 344 403 346 407
rect 346 403 350 407
rect 354 403 357 407
rect 357 403 360 407
rect 344 402 350 403
rect 354 402 360 403
rect 1368 407 1374 408
rect 1378 407 1384 408
rect 1368 403 1370 407
rect 1370 403 1374 407
rect 1378 403 1381 407
rect 1381 403 1384 407
rect 1368 402 1374 403
rect 1378 402 1384 403
rect 2392 407 2398 408
rect 2402 407 2408 408
rect 2392 403 2394 407
rect 2394 403 2398 407
rect 2402 403 2405 407
rect 2405 403 2408 407
rect 2392 402 2398 403
rect 2402 402 2408 403
rect 3416 407 3422 408
rect 3426 407 3432 408
rect 3416 403 3418 407
rect 3418 403 3422 407
rect 3426 403 3429 407
rect 3429 403 3432 407
rect 3416 402 3422 403
rect 3426 402 3432 403
rect 4440 407 4446 408
rect 4450 407 4456 408
rect 4440 403 4442 407
rect 4442 403 4446 407
rect 4450 403 4453 407
rect 4453 403 4456 407
rect 4440 402 4446 403
rect 4450 402 4456 403
rect 856 307 862 308
rect 866 307 872 308
rect 856 303 858 307
rect 858 303 862 307
rect 866 303 869 307
rect 869 303 872 307
rect 856 302 862 303
rect 866 302 872 303
rect 1872 307 1878 308
rect 1882 307 1888 308
rect 1872 303 1874 307
rect 1874 303 1878 307
rect 1882 303 1885 307
rect 1885 303 1888 307
rect 1872 302 1878 303
rect 1882 302 1888 303
rect 2904 307 2910 308
rect 2914 307 2920 308
rect 2904 303 2906 307
rect 2906 303 2910 307
rect 2914 303 2917 307
rect 2917 303 2920 307
rect 2904 302 2910 303
rect 2914 302 2920 303
rect 3928 307 3934 308
rect 3938 307 3944 308
rect 3928 303 3930 307
rect 3930 303 3934 307
rect 3938 303 3941 307
rect 3941 303 3944 307
rect 3928 302 3934 303
rect 3938 302 3944 303
rect 4952 307 4958 308
rect 4962 307 4968 308
rect 4952 303 4954 307
rect 4954 303 4958 307
rect 4962 303 4965 307
rect 4965 303 4968 307
rect 4952 302 4958 303
rect 4962 302 4968 303
rect 344 207 350 208
rect 354 207 360 208
rect 344 203 346 207
rect 346 203 350 207
rect 354 203 357 207
rect 357 203 360 207
rect 344 202 350 203
rect 354 202 360 203
rect 1368 207 1374 208
rect 1378 207 1384 208
rect 1368 203 1370 207
rect 1370 203 1374 207
rect 1378 203 1381 207
rect 1381 203 1384 207
rect 1368 202 1374 203
rect 1378 202 1384 203
rect 2392 207 2398 208
rect 2402 207 2408 208
rect 2392 203 2394 207
rect 2394 203 2398 207
rect 2402 203 2405 207
rect 2405 203 2408 207
rect 2392 202 2398 203
rect 2402 202 2408 203
rect 3416 207 3422 208
rect 3426 207 3432 208
rect 3416 203 3418 207
rect 3418 203 3422 207
rect 3426 203 3429 207
rect 3429 203 3432 207
rect 3416 202 3422 203
rect 3426 202 3432 203
rect 4440 207 4446 208
rect 4450 207 4456 208
rect 4440 203 4442 207
rect 4442 203 4446 207
rect 4450 203 4453 207
rect 4453 203 4456 207
rect 4440 202 4446 203
rect 4450 202 4456 203
rect 856 107 862 108
rect 866 107 872 108
rect 856 103 858 107
rect 858 103 862 107
rect 866 103 869 107
rect 869 103 872 107
rect 856 102 862 103
rect 866 102 872 103
rect 1872 107 1878 108
rect 1882 107 1888 108
rect 1872 103 1874 107
rect 1874 103 1878 107
rect 1882 103 1885 107
rect 1885 103 1888 107
rect 1872 102 1878 103
rect 1882 102 1888 103
rect 2904 107 2910 108
rect 2914 107 2920 108
rect 2904 103 2906 107
rect 2906 103 2910 107
rect 2914 103 2917 107
rect 2917 103 2920 107
rect 2904 102 2910 103
rect 2914 102 2920 103
rect 3928 107 3934 108
rect 3938 107 3944 108
rect 3928 103 3930 107
rect 3930 103 3934 107
rect 3938 103 3941 107
rect 3941 103 3944 107
rect 3928 102 3934 103
rect 3938 102 3944 103
rect 4952 107 4958 108
rect 4962 107 4968 108
rect 4952 103 4954 107
rect 4954 103 4958 107
rect 4962 103 4965 107
rect 4965 103 4968 107
rect 4952 102 4958 103
rect 4962 102 4968 103
rect 5293 77 5299 83
rect 344 7 350 8
rect 354 7 360 8
rect 344 3 346 7
rect 346 3 350 7
rect 354 3 357 7
rect 357 3 360 7
rect 344 2 350 3
rect 354 2 360 3
rect 1368 7 1374 8
rect 1378 7 1384 8
rect 1368 3 1370 7
rect 1370 3 1374 7
rect 1378 3 1381 7
rect 1381 3 1384 7
rect 1368 2 1374 3
rect 1378 2 1384 3
rect 2392 7 2398 8
rect 2402 7 2408 8
rect 2392 3 2394 7
rect 2394 3 2398 7
rect 2402 3 2405 7
rect 2405 3 2408 7
rect 2392 2 2398 3
rect 2402 2 2408 3
rect 3416 7 3422 8
rect 3426 7 3432 8
rect 3416 3 3418 7
rect 3418 3 3422 7
rect 3426 3 3429 7
rect 3429 3 3432 7
rect 3416 2 3422 3
rect 3426 2 3432 3
rect 4440 7 4446 8
rect 4450 7 4456 8
rect 4440 3 4442 7
rect 4442 3 4446 7
rect 4450 3 4453 7
rect 4453 3 4456 7
rect 4440 2 4446 3
rect 4450 2 4456 3
<< metal6 >>
rect 344 3608 360 3730
rect 350 3602 354 3608
rect 344 3408 360 3602
rect 350 3402 354 3408
rect 344 3208 360 3402
rect 350 3202 354 3208
rect 344 3008 360 3202
rect 350 3002 354 3008
rect 344 2808 360 3002
rect 350 2802 354 2808
rect 344 2608 360 2802
rect 350 2602 354 2608
rect 344 2408 360 2602
rect 350 2402 354 2408
rect 344 2208 360 2402
rect 350 2202 354 2208
rect 344 2008 360 2202
rect 350 2002 354 2008
rect 344 1808 360 2002
rect 350 1802 354 1808
rect 344 1608 360 1802
rect 350 1602 354 1608
rect 344 1408 360 1602
rect 350 1402 354 1408
rect 344 1208 360 1402
rect 350 1202 354 1208
rect 344 1008 360 1202
rect 350 1002 354 1008
rect 344 808 360 1002
rect 350 802 354 808
rect 344 608 360 802
rect 350 602 354 608
rect 344 408 360 602
rect 350 402 354 408
rect 344 208 360 402
rect 350 202 354 208
rect 344 8 360 202
rect 350 2 354 8
rect 344 -30 360 2
rect 856 3708 872 3730
rect 862 3702 866 3708
rect 856 3508 872 3702
rect 862 3502 866 3508
rect 856 3308 872 3502
rect 862 3302 866 3308
rect 856 3108 872 3302
rect 862 3102 866 3108
rect 856 2908 872 3102
rect 862 2902 866 2908
rect 856 2708 872 2902
rect 862 2702 866 2708
rect 856 2508 872 2702
rect 862 2502 866 2508
rect 856 2308 872 2502
rect 862 2302 866 2308
rect 856 2108 872 2302
rect 862 2102 866 2108
rect 856 1908 872 2102
rect 862 1902 866 1908
rect 856 1708 872 1902
rect 862 1702 866 1708
rect 856 1508 872 1702
rect 862 1502 866 1508
rect 856 1308 872 1502
rect 862 1302 866 1308
rect 856 1108 872 1302
rect 862 1102 866 1108
rect 856 908 872 1102
rect 862 902 866 908
rect 856 708 872 902
rect 862 702 866 708
rect 856 508 872 702
rect 862 502 866 508
rect 856 308 872 502
rect 862 302 866 308
rect 856 108 872 302
rect 862 102 866 108
rect 856 -30 872 102
rect 1368 3608 1384 3730
rect 1374 3602 1378 3608
rect 1368 3408 1384 3602
rect 1374 3402 1378 3408
rect 1368 3208 1384 3402
rect 1374 3202 1378 3208
rect 1368 3008 1384 3202
rect 1374 3002 1378 3008
rect 1368 2808 1384 3002
rect 1374 2802 1378 2808
rect 1368 2608 1384 2802
rect 1374 2602 1378 2608
rect 1368 2408 1384 2602
rect 1374 2402 1378 2408
rect 1368 2208 1384 2402
rect 1374 2202 1378 2208
rect 1368 2008 1384 2202
rect 1374 2002 1378 2008
rect 1368 1808 1384 2002
rect 1374 1802 1378 1808
rect 1368 1608 1384 1802
rect 1374 1602 1378 1608
rect 1368 1408 1384 1602
rect 1374 1402 1378 1408
rect 1368 1208 1384 1402
rect 1374 1202 1378 1208
rect 1368 1008 1384 1202
rect 1374 1002 1378 1008
rect 1368 808 1384 1002
rect 1374 802 1378 808
rect 1368 608 1384 802
rect 1374 602 1378 608
rect 1368 408 1384 602
rect 1374 402 1378 408
rect 1368 208 1384 402
rect 1374 202 1378 208
rect 1368 8 1384 202
rect 1374 2 1378 8
rect 1368 -30 1384 2
rect 1872 3708 1888 3730
rect 1878 3702 1882 3708
rect 1872 3508 1888 3702
rect 1878 3502 1882 3508
rect 1872 3308 1888 3502
rect 1878 3302 1882 3308
rect 1872 3108 1888 3302
rect 1878 3102 1882 3108
rect 1872 2908 1888 3102
rect 1878 2902 1882 2908
rect 1872 2708 1888 2902
rect 1878 2702 1882 2708
rect 1872 2508 1888 2702
rect 1878 2502 1882 2508
rect 1872 2308 1888 2502
rect 2392 3608 2408 3730
rect 2398 3602 2402 3608
rect 2392 3408 2408 3602
rect 2398 3402 2402 3408
rect 2392 3208 2408 3402
rect 2398 3202 2402 3208
rect 2392 3008 2408 3202
rect 2398 3002 2402 3008
rect 2392 2808 2408 3002
rect 2398 2802 2402 2808
rect 2392 2608 2408 2802
rect 2398 2602 2402 2608
rect 1878 2302 1882 2308
rect 1872 2108 1888 2302
rect 1878 2102 1882 2108
rect 1872 1908 1888 2102
rect 1878 1902 1882 1908
rect 1872 1708 1888 1902
rect 1878 1702 1882 1708
rect 1872 1508 1888 1702
rect 1878 1502 1882 1508
rect 1872 1308 1888 1502
rect 1878 1302 1882 1308
rect 1872 1108 1888 1302
rect 2141 1273 2146 2467
rect 2392 2408 2408 2602
rect 2904 3708 2920 3730
rect 2910 3702 2914 3708
rect 2904 3508 2920 3702
rect 2910 3502 2914 3508
rect 2904 3308 2920 3502
rect 2910 3302 2914 3308
rect 2904 3108 2920 3302
rect 2910 3102 2914 3108
rect 2904 2908 2920 3102
rect 2910 2902 2914 2908
rect 2904 2708 2920 2902
rect 2910 2702 2914 2708
rect 2904 2508 2920 2702
rect 2910 2502 2914 2508
rect 2398 2402 2402 2408
rect 2392 2208 2408 2402
rect 2398 2202 2402 2208
rect 2392 2008 2408 2202
rect 2621 2043 2626 2437
rect 2904 2308 2920 2502
rect 2910 2302 2914 2308
rect 2904 2108 2920 2302
rect 2910 2102 2914 2108
rect 2398 2002 2402 2008
rect 2392 1808 2408 2002
rect 2398 1802 2402 1808
rect 2392 1608 2408 1802
rect 2398 1602 2402 1608
rect 2392 1408 2408 1602
rect 2398 1402 2402 1408
rect 1878 1102 1882 1108
rect 1872 908 1888 1102
rect 1878 902 1882 908
rect 1872 708 1888 902
rect 1878 702 1882 708
rect 1872 508 1888 702
rect 1878 502 1882 508
rect 1872 308 1888 502
rect 1878 302 1882 308
rect 1872 108 1888 302
rect 1878 102 1882 108
rect 1872 -30 1888 102
rect 2392 1208 2408 1402
rect 2398 1202 2402 1208
rect 2392 1008 2408 1202
rect 2398 1002 2402 1008
rect 2392 808 2408 1002
rect 2398 802 2402 808
rect 2392 608 2408 802
rect 2398 602 2402 608
rect 2392 408 2408 602
rect 2398 402 2402 408
rect 2392 208 2408 402
rect 2398 202 2402 208
rect 2392 8 2408 202
rect 2398 2 2402 8
rect 2392 -30 2408 2
rect 2904 1908 2920 2102
rect 2910 1902 2914 1908
rect 2904 1708 2920 1902
rect 2910 1702 2914 1708
rect 2904 1508 2920 1702
rect 2910 1502 2914 1508
rect 2904 1308 2920 1502
rect 2910 1302 2914 1308
rect 2904 1108 2920 1302
rect 2910 1102 2914 1108
rect 2904 908 2920 1102
rect 2910 902 2914 908
rect 2904 708 2920 902
rect 2910 702 2914 708
rect 2904 508 2920 702
rect 2910 502 2914 508
rect 2904 308 2920 502
rect 2910 302 2914 308
rect 2904 108 2920 302
rect 2910 102 2914 108
rect 2904 -30 2920 102
rect 3416 3608 3432 3730
rect 3422 3602 3426 3608
rect 3416 3408 3432 3602
rect 3422 3402 3426 3408
rect 3416 3208 3432 3402
rect 3422 3202 3426 3208
rect 3416 3008 3432 3202
rect 3422 3002 3426 3008
rect 3416 2808 3432 3002
rect 3422 2802 3426 2808
rect 3416 2608 3432 2802
rect 3422 2602 3426 2608
rect 3416 2408 3432 2602
rect 3422 2402 3426 2408
rect 3416 2208 3432 2402
rect 3422 2202 3426 2208
rect 3416 2008 3432 2202
rect 3422 2002 3426 2008
rect 3416 1808 3432 2002
rect 3422 1802 3426 1808
rect 3416 1608 3432 1802
rect 3422 1602 3426 1608
rect 3416 1408 3432 1602
rect 3422 1402 3426 1408
rect 3416 1208 3432 1402
rect 3422 1202 3426 1208
rect 3416 1008 3432 1202
rect 3422 1002 3426 1008
rect 3416 808 3432 1002
rect 3422 802 3426 808
rect 3416 608 3432 802
rect 3422 602 3426 608
rect 3416 408 3432 602
rect 3422 402 3426 408
rect 3416 208 3432 402
rect 3422 202 3426 208
rect 3416 8 3432 202
rect 3422 2 3426 8
rect 3416 -30 3432 2
rect 3928 3708 3944 3730
rect 3934 3702 3938 3708
rect 3928 3508 3944 3702
rect 3934 3502 3938 3508
rect 3928 3308 3944 3502
rect 3934 3302 3938 3308
rect 3928 3108 3944 3302
rect 3934 3102 3938 3108
rect 3928 2908 3944 3102
rect 3934 2902 3938 2908
rect 3928 2708 3944 2902
rect 3934 2702 3938 2708
rect 3928 2508 3944 2702
rect 3934 2502 3938 2508
rect 3928 2308 3944 2502
rect 3934 2302 3938 2308
rect 3928 2108 3944 2302
rect 3934 2102 3938 2108
rect 3928 1908 3944 2102
rect 3934 1902 3938 1908
rect 3928 1708 3944 1902
rect 3934 1702 3938 1708
rect 3928 1508 3944 1702
rect 3934 1502 3938 1508
rect 3928 1308 3944 1502
rect 3934 1302 3938 1308
rect 3928 1108 3944 1302
rect 3934 1102 3938 1108
rect 3928 908 3944 1102
rect 3934 902 3938 908
rect 3928 708 3944 902
rect 3934 702 3938 708
rect 3928 508 3944 702
rect 3934 502 3938 508
rect 3928 308 3944 502
rect 3934 302 3938 308
rect 3928 108 3944 302
rect 3934 102 3938 108
rect 3928 -30 3944 102
rect 4440 3608 4456 3730
rect 4446 3602 4450 3608
rect 4440 3408 4456 3602
rect 4446 3402 4450 3408
rect 4440 3208 4456 3402
rect 4446 3202 4450 3208
rect 4440 3008 4456 3202
rect 4446 3002 4450 3008
rect 4440 2808 4456 3002
rect 4446 2802 4450 2808
rect 4440 2608 4456 2802
rect 4446 2602 4450 2608
rect 4440 2408 4456 2602
rect 4446 2402 4450 2408
rect 4440 2208 4456 2402
rect 4446 2202 4450 2208
rect 4440 2008 4456 2202
rect 4446 2002 4450 2008
rect 4440 1808 4456 2002
rect 4446 1802 4450 1808
rect 4440 1608 4456 1802
rect 4446 1602 4450 1608
rect 4440 1408 4456 1602
rect 4446 1402 4450 1408
rect 4440 1208 4456 1402
rect 4446 1202 4450 1208
rect 4440 1008 4456 1202
rect 4446 1002 4450 1008
rect 4440 808 4456 1002
rect 4446 802 4450 808
rect 4440 608 4456 802
rect 4446 602 4450 608
rect 4440 408 4456 602
rect 4446 402 4450 408
rect 4440 208 4456 402
rect 4446 202 4450 208
rect 4440 8 4456 202
rect 4446 2 4450 8
rect 4440 -30 4456 2
rect 4952 3708 4968 3730
rect 4958 3702 4962 3708
rect 4952 3508 4968 3702
rect 4958 3502 4962 3508
rect 4952 3308 4968 3502
rect 4958 3302 4962 3308
rect 4952 3108 4968 3302
rect 4958 3102 4962 3108
rect 4952 2908 4968 3102
rect 4958 2902 4962 2908
rect 4952 2708 4968 2902
rect 4958 2702 4962 2708
rect 4952 2508 4968 2702
rect 4958 2502 4962 2508
rect 4952 2308 4968 2502
rect 4958 2302 4962 2308
rect 4952 2108 4968 2302
rect 5213 2173 5218 2407
rect 4958 2102 4962 2108
rect 4952 1908 4968 2102
rect 4958 1902 4962 1908
rect 4952 1708 4968 1902
rect 4958 1702 4962 1708
rect 4952 1508 4968 1702
rect 4958 1502 4962 1508
rect 4952 1308 4968 1502
rect 4958 1302 4962 1308
rect 4952 1108 4968 1302
rect 5213 1283 5218 2147
rect 5229 2133 5234 3547
rect 5229 1683 5234 2107
rect 4958 1102 4962 1108
rect 4952 908 4968 1102
rect 4958 902 4962 908
rect 4952 708 4968 902
rect 5245 873 5250 3167
rect 4958 702 4962 708
rect 4952 508 4968 702
rect 5261 533 5266 3457
rect 5277 3063 5282 3437
rect 5277 2643 5282 2987
rect 5293 2683 5298 3067
rect 5277 2143 5282 2627
rect 5277 2103 5282 2127
rect 5277 563 5282 1287
rect 4958 502 4962 508
rect 4952 308 4968 502
rect 4958 302 4962 308
rect 4952 108 4968 302
rect 4958 102 4962 108
rect 4952 -30 4968 102
rect 5293 83 5298 2677
rect 5309 2583 5314 3067
rect 5309 853 5314 2567
rect 5357 863 5362 2517
use BUFX2  BUFX2_106
timestamp 1625156677
transform 1 0 4 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_35
timestamp 1625156677
transform 1 0 28 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_112
timestamp 1625156677
transform 1 0 52 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_98
timestamp 1625156677
transform 1 0 76 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_58
timestamp 1625156677
transform 1 0 100 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_38
timestamp 1625156677
transform -1 0 148 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_56
timestamp 1625156677
transform -1 0 172 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_65
timestamp 1625156677
transform 1 0 172 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_130
timestamp 1625156677
transform 1 0 196 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_137
timestamp 1625156677
transform 1 0 220 0 -1 3705
box -2 -3 26 103
use NAND3X1  NAND3X1_390
timestamp 1625156677
transform -1 0 276 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_259
timestamp 1625156677
transform 1 0 276 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_326
timestamp 1625156677
transform -1 0 324 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_394
timestamp 1625156677
transform -1 0 356 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_0_0
timestamp 1625156677
transform 1 0 356 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_0_1
timestamp 1625156677
transform 1 0 364 0 -1 3705
box -2 -3 10 103
use AOI21X1  AOI21X1_260
timestamp 1625156677
transform 1 0 372 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_268
timestamp 1625156677
transform 1 0 404 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_424
timestamp 1625156677
transform -1 0 460 0 -1 3705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_177
timestamp 1625156677
transform -1 0 516 0 -1 3705
box -2 -3 58 103
use NOR2X1  NOR2X1_269
timestamp 1625156677
transform -1 0 540 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_430
timestamp 1625156677
transform -1 0 572 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_423
timestamp 1625156677
transform -1 0 604 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_261
timestamp 1625156677
transform 1 0 604 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_387
timestamp 1625156677
transform 1 0 636 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_463
timestamp 1625156677
transform -1 0 692 0 -1 3705
box -2 -3 26 103
use NOR3X1  NOR3X1_71
timestamp 1625156677
transform -1 0 756 0 -1 3705
box -2 -3 66 103
use INVX1  INVX1_325
timestamp 1625156677
transform -1 0 772 0 -1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_461
timestamp 1625156677
transform 1 0 772 0 -1 3705
box -2 -3 26 103
use NAND3X1  NAND3X1_385
timestamp 1625156677
transform 1 0 796 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_464
timestamp 1625156677
transform -1 0 852 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_1_0
timestamp 1625156677
transform -1 0 860 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_1_1
timestamp 1625156677
transform -1 0 868 0 -1 3705
box -2 -3 10 103
use NAND3X1  NAND3X1_393
timestamp 1625156677
transform -1 0 900 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_323
timestamp 1625156677
transform -1 0 916 0 -1 3705
box -2 -3 18 103
use NOR2X1  NOR2X1_265
timestamp 1625156677
transform -1 0 940 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_417
timestamp 1625156677
transform -1 0 972 0 -1 3705
box -2 -3 34 103
use NOR2X1  NOR2X1_266
timestamp 1625156677
transform -1 0 996 0 -1 3705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_176
timestamp 1625156677
transform -1 0 1052 0 -1 3705
box -2 -3 58 103
use BUFX2  BUFX2_217
timestamp 1625156677
transform 1 0 1052 0 -1 3705
box -2 -3 26 103
use XOR2X1  XOR2X1_238
timestamp 1625156677
transform 1 0 1076 0 -1 3705
box -2 -3 58 103
use BUFX2  BUFX2_215
timestamp 1625156677
transform -1 0 1156 0 -1 3705
box -2 -3 26 103
use XOR2X1  XOR2X1_237
timestamp 1625156677
transform 1 0 1156 0 -1 3705
box -2 -3 58 103
use INVX1  INVX1_366
timestamp 1625156677
transform 1 0 1212 0 -1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_460
timestamp 1625156677
transform 1 0 1228 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_367
timestamp 1625156677
transform -1 0 1276 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_414
timestamp 1625156677
transform -1 0 1308 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_365
timestamp 1625156677
transform -1 0 1324 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_415
timestamp 1625156677
transform -1 0 1356 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_2_0
timestamp 1625156677
transform -1 0 1364 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_2_1
timestamp 1625156677
transform -1 0 1372 0 -1 3705
box -2 -3 10 103
use XOR2X1  XOR2X1_236
timestamp 1625156677
transform -1 0 1428 0 -1 3705
box -2 -3 58 103
use NOR2X1  NOR2X1_288
timestamp 1625156677
transform -1 0 1452 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_457
timestamp 1625156677
transform 1 0 1452 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_412
timestamp 1625156677
transform -1 0 1516 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_454
timestamp 1625156677
transform 1 0 1516 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_363
timestamp 1625156677
transform 1 0 1548 0 -1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_465
timestamp 1625156677
transform 1 0 1564 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_360
timestamp 1625156677
transform -1 0 1612 0 -1 3705
box -2 -3 18 103
use NAND2X1  NAND2X1_506
timestamp 1625156677
transform 1 0 1612 0 -1 3705
box -2 -3 26 103
use NAND2X1  NAND2X1_498
timestamp 1625156677
transform 1 0 1636 0 -1 3705
box -2 -3 26 103
use AOI21X1  AOI21X1_278
timestamp 1625156677
transform 1 0 1660 0 -1 3705
box -2 -3 34 103
use XOR2X1  XOR2X1_234
timestamp 1625156677
transform 1 0 1692 0 -1 3705
box -2 -3 58 103
use XOR2X1  XOR2X1_256
timestamp 1625156677
transform 1 0 1748 0 -1 3705
box -2 -3 58 103
use NOR2X1  NOR2X1_286
timestamp 1625156677
transform 1 0 1804 0 -1 3705
box -2 -3 26 103
use NAND3X1  NAND3X1_410
timestamp 1625156677
transform 1 0 1828 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_495
timestamp 1625156677
transform -1 0 1884 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_3_0
timestamp 1625156677
transform 1 0 1884 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_3_1
timestamp 1625156677
transform 1 0 1892 0 -1 3705
box -2 -3 10 103
use AND2X2  AND2X2_134
timestamp 1625156677
transform 1 0 1900 0 -1 3705
box -2 -3 34 103
use NAND2X1  NAND2X1_496
timestamp 1625156677
transform -1 0 1956 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_451
timestamp 1625156677
transform 1 0 1956 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_358
timestamp 1625156677
transform -1 0 2004 0 -1 3705
box -2 -3 18 103
use BUFX2  BUFX2_223
timestamp 1625156677
transform 1 0 2004 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_84
timestamp 1625156677
transform -1 0 2052 0 -1 3705
box -2 -3 26 103
use INVX1  INVX1_385
timestamp 1625156677
transform 1 0 2052 0 -1 3705
box -2 -3 18 103
use BUFX2  BUFX2_123
timestamp 1625156677
transform 1 0 2068 0 -1 3705
box -2 -3 26 103
use INVX1  INVX1_384
timestamp 1625156677
transform 1 0 2092 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_428
timestamp 1625156677
transform -1 0 2140 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_427
timestamp 1625156677
transform 1 0 2140 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_478
timestamp 1625156677
transform -1 0 2204 0 -1 3705
box -2 -3 34 103
use BUFX2  BUFX2_67
timestamp 1625156677
transform 1 0 2204 0 -1 3705
box -2 -3 26 103
use INVX1  INVX1_404
timestamp 1625156677
transform 1 0 2228 0 -1 3705
box -2 -3 18 103
use OAI21X1  OAI21X1_498
timestamp 1625156677
transform 1 0 2244 0 -1 3705
box -2 -3 34 103
use OAI21X1  OAI21X1_497
timestamp 1625156677
transform 1 0 2276 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_405
timestamp 1625156677
transform -1 0 2324 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_440
timestamp 1625156677
transform -1 0 2356 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_403
timestamp 1625156677
transform 1 0 2356 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_441
timestamp 1625156677
transform -1 0 2404 0 -1 3705
box -2 -3 34 103
use FILL  FILL_36_4_0
timestamp 1625156677
transform 1 0 2404 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_4_1
timestamp 1625156677
transform 1 0 2412 0 -1 3705
box -2 -3 10 103
use AOI21X1  AOI21X1_291
timestamp 1625156677
transform 1 0 2420 0 -1 3705
box -2 -3 34 103
use NAND3X1  NAND3X1_442
timestamp 1625156677
transform 1 0 2452 0 -1 3705
box -2 -3 34 103
use INVX1  INVX1_402
timestamp 1625156677
transform -1 0 2500 0 -1 3705
box -2 -3 18 103
use NAND3X1  NAND3X1_446
timestamp 1625156677
transform -1 0 2532 0 -1 3705
box -2 -3 34 103
use AOI21X1  AOI21X1_292
timestamp 1625156677
transform 1 0 2532 0 -1 3705
box -2 -3 34 103
use BUFX2  BUFX2_82
timestamp 1625156677
transform -1 0 2588 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_75
timestamp 1625156677
transform 1 0 2588 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_111
timestamp 1625156677
transform 1 0 2612 0 -1 3705
box -2 -3 26 103
use NOR2X1  NOR2X1_316
timestamp 1625156677
transform 1 0 2636 0 -1 3705
box -2 -3 26 103
use OAI21X1  OAI21X1_500
timestamp 1625156677
transform -1 0 2692 0 -1 3705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_193
timestamp 1625156677
transform 1 0 2692 0 -1 3705
box -2 -3 58 103
use BUFX2  BUFX2_8
timestamp 1625156677
transform -1 0 2772 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1625156677
transform -1 0 2868 0 -1 3705
box -2 -3 98 103
use NOR3X1  NOR3X1_8
timestamp 1625156677
transform -1 0 2932 0 -1 3705
box -2 -3 66 103
use FILL  FILL_36_5_0
timestamp 1625156677
transform -1 0 2940 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_5_1
timestamp 1625156677
transform -1 0 2948 0 -1 3705
box -2 -3 10 103
use BUFX2  BUFX2_1
timestamp 1625156677
transform -1 0 2972 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_4
timestamp 1625156677
transform -1 0 2996 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1625156677
transform -1 0 3092 0 -1 3705
box -2 -3 98 103
use NOR3X1  NOR3X1_1
timestamp 1625156677
transform 1 0 3092 0 -1 3705
box -2 -3 66 103
use BUFX2  BUFX2_2
timestamp 1625156677
transform -1 0 3180 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1625156677
transform 1 0 3180 0 -1 3705
box -2 -3 98 103
use BUFX2  BUFX2_6
timestamp 1625156677
transform 1 0 3276 0 -1 3705
box -2 -3 26 103
use NOR3X1  NOR3X1_6
timestamp 1625156677
transform 1 0 3300 0 -1 3705
box -2 -3 66 103
use BUFX2  BUFX2_3
timestamp 1625156677
transform 1 0 3364 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_24
timestamp 1625156677
transform -1 0 3412 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_6_0
timestamp 1625156677
transform -1 0 3420 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_6_1
timestamp 1625156677
transform -1 0 3428 0 -1 3705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1625156677
transform -1 0 3524 0 -1 3705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1625156677
transform 1 0 3524 0 -1 3705
box -2 -3 98 103
use BUFX2  BUFX2_22
timestamp 1625156677
transform -1 0 3644 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_25
timestamp 1625156677
transform 1 0 3644 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_7
timestamp 1625156677
transform 1 0 3668 0 -1 3705
box -2 -3 26 103
use MUX2X1  MUX2X1_7
timestamp 1625156677
transform 1 0 3692 0 -1 3705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1625156677
transform -1 0 3836 0 -1 3705
box -2 -3 98 103
use NOR3X1  NOR3X1_7
timestamp 1625156677
transform 1 0 3836 0 -1 3705
box -2 -3 66 103
use MUX2X1  MUX2X1_21
timestamp 1625156677
transform 1 0 3900 0 -1 3705
box -2 -3 50 103
use FILL  FILL_36_7_0
timestamp 1625156677
transform 1 0 3948 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_7_1
timestamp 1625156677
transform 1 0 3956 0 -1 3705
box -2 -3 10 103
use BUFX2  BUFX2_21
timestamp 1625156677
transform 1 0 3964 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1625156677
transform -1 0 4084 0 -1 3705
box -2 -3 98 103
use NOR3X1  NOR3X1_21
timestamp 1625156677
transform 1 0 4084 0 -1 3705
box -2 -3 66 103
use NOR3X1  NOR3X1_13
timestamp 1625156677
transform -1 0 4212 0 -1 3705
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1625156677
transform 1 0 4212 0 -1 3705
box -2 -3 98 103
use INVX1  INVX1_7
timestamp 1625156677
transform 1 0 4308 0 -1 3705
box -2 -3 18 103
use AOI22X1  AOI22X1_4
timestamp 1625156677
transform 1 0 4324 0 -1 3705
box -2 -3 42 103
use OAI22X1  OAI22X1_9
timestamp 1625156677
transform 1 0 4364 0 -1 3705
box -2 -3 42 103
use INVX1  INVX1_8
timestamp 1625156677
transform -1 0 4420 0 -1 3705
box -2 -3 18 103
use BUFX2  BUFX2_13
timestamp 1625156677
transform 1 0 4420 0 -1 3705
box -2 -3 26 103
use FILL  FILL_36_8_0
timestamp 1625156677
transform -1 0 4452 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_8_1
timestamp 1625156677
transform -1 0 4460 0 -1 3705
box -2 -3 10 103
use MUX2X1  MUX2X1_13
timestamp 1625156677
transform -1 0 4508 0 -1 3705
box -2 -3 50 103
use INVX2  INVX2_1
timestamp 1625156677
transform 1 0 4508 0 -1 3705
box -2 -3 18 103
use MUX2X1  MUX2X1_14
timestamp 1625156677
transform 1 0 4524 0 -1 3705
box -2 -3 50 103
use BUFX2  BUFX2_14
timestamp 1625156677
transform 1 0 4572 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1625156677
transform -1 0 4692 0 -1 3705
box -2 -3 98 103
use NOR3X1  NOR3X1_14
timestamp 1625156677
transform 1 0 4692 0 -1 3705
box -2 -3 66 103
use BUFX2  BUFX2_19
timestamp 1625156677
transform 1 0 4756 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1625156677
transform -1 0 4876 0 -1 3705
box -2 -3 98 103
use NOR3X1  NOR3X1_19
timestamp 1625156677
transform 1 0 4876 0 -1 3705
box -2 -3 66 103
use FILL  FILL_36_9_0
timestamp 1625156677
transform -1 0 4948 0 -1 3705
box -2 -3 10 103
use FILL  FILL_36_9_1
timestamp 1625156677
transform -1 0 4956 0 -1 3705
box -2 -3 10 103
use NOR3X1  NOR3X1_11
timestamp 1625156677
transform -1 0 5020 0 -1 3705
box -2 -3 66 103
use MUX2X1  MUX2X1_11
timestamp 1625156677
transform 1 0 5020 0 -1 3705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1625156677
transform 1 0 5068 0 -1 3705
box -2 -3 98 103
use BUFX2  BUFX2_11
timestamp 1625156677
transform 1 0 5164 0 -1 3705
box -2 -3 26 103
use BUFX2  BUFX2_40
timestamp 1625156677
transform 1 0 5188 0 -1 3705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_205
timestamp 1625156677
transform -1 0 5308 0 -1 3705
box -2 -3 98 103
use FILL  FILL_37_1
timestamp 1625156677
transform -1 0 5316 0 -1 3705
box -2 -3 10 103
use NOR2X1  NOR2X1_252
timestamp 1625156677
transform 1 0 4 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_408
timestamp 1625156677
transform 1 0 28 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_303
timestamp 1625156677
transform -1 0 76 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_441
timestamp 1625156677
transform 1 0 76 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_449
timestamp 1625156677
transform -1 0 124 0 1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_254
timestamp 1625156677
transform 1 0 124 0 1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_388
timestamp 1625156677
transform -1 0 188 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_327
timestamp 1625156677
transform -1 0 204 0 1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_389
timestamp 1625156677
transform -1 0 236 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_328
timestamp 1625156677
transform -1 0 252 0 1 3505
box -2 -3 18 103
use INVX1  INVX1_329
timestamp 1625156677
transform 1 0 252 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_422
timestamp 1625156677
transform -1 0 300 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_474
timestamp 1625156677
transform -1 0 324 0 1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_265
timestamp 1625156677
transform -1 0 356 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_0_0
timestamp 1625156677
transform 1 0 356 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_0_1
timestamp 1625156677
transform 1 0 364 0 1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_467
timestamp 1625156677
transform 1 0 372 0 1 3505
box -2 -3 26 103
use XOR2X1  XOR2X1_233
timestamp 1625156677
transform -1 0 452 0 1 3505
box -2 -3 58 103
use NAND2X1  NAND2X1_469
timestamp 1625156677
transform 1 0 452 0 1 3505
box -2 -3 26 103
use XOR2X1  XOR2X1_239
timestamp 1625156677
transform 1 0 476 0 1 3505
box -2 -3 58 103
use AOI21X1  AOI21X1_264
timestamp 1625156677
transform -1 0 564 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_429
timestamp 1625156677
transform 1 0 564 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_336
timestamp 1625156677
transform -1 0 612 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_420
timestamp 1625156677
transform 1 0 612 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_267
timestamp 1625156677
transform -1 0 668 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_462
timestamp 1625156677
transform -1 0 692 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_324
timestamp 1625156677
transform 1 0 692 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_419
timestamp 1625156677
transform -1 0 740 0 1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_386
timestamp 1625156677
transform -1 0 772 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_332
timestamp 1625156677
transform 1 0 772 0 1 3505
box -2 -3 18 103
use AOI21X1  AOI21X1_263
timestamp 1625156677
transform -1 0 820 0 1 3505
box -2 -3 34 103
use NOR3X1  NOR3X1_72
timestamp 1625156677
transform -1 0 884 0 1 3505
box -2 -3 66 103
use FILL  FILL_35_1_0
timestamp 1625156677
transform -1 0 892 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_1_1
timestamp 1625156677
transform -1 0 900 0 1 3505
box -2 -3 10 103
use INVX2  INVX2_66
timestamp 1625156677
transform -1 0 916 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_418
timestamp 1625156677
transform 1 0 916 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_415
timestamp 1625156677
transform 1 0 948 0 1 3505
box -2 -3 34 103
use AND2X2  AND2X2_128
timestamp 1625156677
transform 1 0 980 0 1 3505
box -2 -3 34 103
use BUFX2  BUFX2_218
timestamp 1625156677
transform -1 0 1036 0 1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_384
timestamp 1625156677
transform -1 0 1068 0 1 3505
box -2 -3 34 103
use AND2X2  AND2X2_126
timestamp 1625156677
transform -1 0 1100 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_457
timestamp 1625156677
transform -1 0 1124 0 1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_262
timestamp 1625156677
transform 1 0 1124 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_458
timestamp 1625156677
transform -1 0 1172 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_320
timestamp 1625156677
transform -1 0 1188 0 1 3505
box -2 -3 18 103
use XOR2X1  XOR2X1_247
timestamp 1625156677
transform 1 0 1188 0 1 3505
box -2 -3 58 103
use OAI21X1  OAI21X1_459
timestamp 1625156677
transform 1 0 1244 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_275
timestamp 1625156677
transform 1 0 1276 0 1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_416
timestamp 1625156677
transform -1 0 1340 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_364
timestamp 1625156677
transform -1 0 1356 0 1 3505
box -2 -3 18 103
use FILL  FILL_35_2_0
timestamp 1625156677
transform -1 0 1364 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_2_1
timestamp 1625156677
transform -1 0 1372 0 1 3505
box -2 -3 10 103
use NAND3X1  NAND3X1_420
timestamp 1625156677
transform -1 0 1404 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_276
timestamp 1625156677
transform 1 0 1404 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_458
timestamp 1625156677
transform 1 0 1436 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_362
timestamp 1625156677
transform 1 0 1468 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_500
timestamp 1625156677
transform 1 0 1484 0 1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_291
timestamp 1625156677
transform -1 0 1532 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_501
timestamp 1625156677
transform 1 0 1532 0 1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_413
timestamp 1625156677
transform -1 0 1588 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_277
timestamp 1625156677
transform 1 0 1588 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_370
timestamp 1625156677
transform 1 0 1620 0 1 3505
box -2 -3 18 103
use AOI21X1  AOI21X1_279
timestamp 1625156677
transform -1 0 1668 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_502
timestamp 1625156677
transform 1 0 1668 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_461
timestamp 1625156677
transform -1 0 1724 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_499
timestamp 1625156677
transform 1 0 1724 0 1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_411
timestamp 1625156677
transform 1 0 1748 0 1 3505
box -2 -3 34 103
use NOR3X1  NOR3X1_75
timestamp 1625156677
transform -1 0 1844 0 1 3505
box -2 -3 66 103
use OAI21X1  OAI21X1_455
timestamp 1625156677
transform -1 0 1876 0 1 3505
box -2 -3 34 103
use FILL  FILL_35_3_0
timestamp 1625156677
transform -1 0 1884 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_3_1
timestamp 1625156677
transform -1 0 1892 0 1 3505
box -2 -3 10 103
use INVX2  INVX2_68
timestamp 1625156677
transform -1 0 1908 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_456
timestamp 1625156677
transform 1 0 1908 0 1 3505
box -2 -3 34 103
use NOR3X1  NOR3X1_76
timestamp 1625156677
transform 1 0 1940 0 1 3505
box -2 -3 66 103
use OAI21X1  OAI21X1_453
timestamp 1625156677
transform 1 0 2004 0 1 3505
box -2 -3 34 103
use AND2X2  AND2X2_136
timestamp 1625156677
transform 1 0 2036 0 1 3505
box -2 -3 34 103
use XOR2X1  XOR2X1_266
timestamp 1625156677
transform -1 0 2124 0 1 3505
box -2 -3 58 103
use NAND2X1  NAND2X1_531
timestamp 1625156677
transform 1 0 2124 0 1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_429
timestamp 1625156677
transform 1 0 2148 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_283
timestamp 1625156677
transform 1 0 2180 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_479
timestamp 1625156677
transform 1 0 2212 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_383
timestamp 1625156677
transform -1 0 2260 0 1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_433
timestamp 1625156677
transform 1 0 2260 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_386
timestamp 1625156677
transform -1 0 2308 0 1 3505
box -2 -3 18 103
use AOI21X1  AOI21X1_284
timestamp 1625156677
transform 1 0 2308 0 1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_477
timestamp 1625156677
transform 1 0 2340 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_382
timestamp 1625156677
transform 1 0 2372 0 1 3505
box -2 -3 18 103
use FILL  FILL_35_4_0
timestamp 1625156677
transform 1 0 2388 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_4_1
timestamp 1625156677
transform 1 0 2396 0 1 3505
box -2 -3 10 103
use AOI21X1  AOI21X1_285
timestamp 1625156677
transform 1 0 2404 0 1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_426
timestamp 1625156677
transform 1 0 2436 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_303
timestamp 1625156677
transform -1 0 2492 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_520
timestamp 1625156677
transform -1 0 2516 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_519
timestamp 1625156677
transform -1 0 2540 0 1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_318
timestamp 1625156677
transform 1 0 2540 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_501
timestamp 1625156677
transform 1 0 2564 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_542
timestamp 1625156677
transform 1 0 2596 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_406
timestamp 1625156677
transform -1 0 2636 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_541
timestamp 1625156677
transform -1 0 2660 0 1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_443
timestamp 1625156677
transform -1 0 2692 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_407
timestamp 1625156677
transform 1 0 2692 0 1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_444
timestamp 1625156677
transform -1 0 2740 0 1 3505
box -2 -3 34 103
use AOI22X1  AOI22X1_19
timestamp 1625156677
transform 1 0 2740 0 1 3505
box -2 -3 42 103
use NAND2X1  NAND2X1_550
timestamp 1625156677
transform 1 0 2780 0 1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_297
timestamp 1625156677
transform -1 0 2836 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_543
timestamp 1625156677
transform 1 0 2836 0 1 3505
box -2 -3 26 103
use XOR2X1  XOR2X1_269
timestamp 1625156677
transform 1 0 2860 0 1 3505
box -2 -3 58 103
use FILL  FILL_35_5_0
timestamp 1625156677
transform 1 0 2916 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_5_1
timestamp 1625156677
transform 1 0 2924 0 1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_545
timestamp 1625156677
transform 1 0 2932 0 1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_315
timestamp 1625156677
transform -1 0 2980 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_495
timestamp 1625156677
transform 1 0 2980 0 1 3505
box -2 -3 34 103
use INVX1  INVX1_400
timestamp 1625156677
transform -1 0 3028 0 1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_538
timestamp 1625156677
transform 1 0 3028 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_539
timestamp 1625156677
transform 1 0 3052 0 1 3505
box -2 -3 26 103
use MUX2X1  MUX2X1_8
timestamp 1625156677
transform -1 0 3124 0 1 3505
box -2 -3 50 103
use AOI21X1  AOI21X1_293
timestamp 1625156677
transform 1 0 3124 0 1 3505
box -2 -3 34 103
use MUX2X1  MUX2X1_1
timestamp 1625156677
transform -1 0 3204 0 1 3505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1625156677
transform -1 0 3300 0 1 3505
box -2 -3 98 103
use MUX2X1  MUX2X1_6
timestamp 1625156677
transform -1 0 3348 0 1 3505
box -2 -3 50 103
use MUX2X1  MUX2X1_4
timestamp 1625156677
transform 1 0 3348 0 1 3505
box -2 -3 50 103
use FILL  FILL_35_6_0
timestamp 1625156677
transform -1 0 3404 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_6_1
timestamp 1625156677
transform -1 0 3412 0 1 3505
box -2 -3 10 103
use NOR3X1  NOR3X1_4
timestamp 1625156677
transform -1 0 3476 0 1 3505
box -2 -3 66 103
use BUFX2  BUFX2_50
timestamp 1625156677
transform -1 0 3500 0 1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1625156677
transform -1 0 3596 0 1 3505
box -2 -3 98 103
use MUX2X1  MUX2X1_24
timestamp 1625156677
transform -1 0 3644 0 1 3505
box -2 -3 50 103
use NOR3X1  NOR3X1_24
timestamp 1625156677
transform 1 0 3644 0 1 3505
box -2 -3 66 103
use NOR3X1  NOR3X1_22
timestamp 1625156677
transform 1 0 3708 0 1 3505
box -2 -3 66 103
use MUX2X1  MUX2X1_22
timestamp 1625156677
transform -1 0 3820 0 1 3505
box -2 -3 50 103
use BUFX4  BUFX4_12
timestamp 1625156677
transform -1 0 3852 0 1 3505
box -2 -3 34 103
use BUFX2  BUFX2_63
timestamp 1625156677
transform 1 0 3852 0 1 3505
box -2 -3 26 103
use NOR3X1  NOR3X1_23
timestamp 1625156677
transform -1 0 3940 0 1 3505
box -2 -3 66 103
use FILL  FILL_35_7_0
timestamp 1625156677
transform 1 0 3940 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_7_1
timestamp 1625156677
transform 1 0 3948 0 1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1625156677
transform 1 0 3956 0 1 3505
box -2 -3 98 103
use MUX2X1  MUX2X1_23
timestamp 1625156677
transform -1 0 4100 0 1 3505
box -2 -3 50 103
use BUFX2  BUFX2_23
timestamp 1625156677
transform 1 0 4100 0 1 3505
box -2 -3 26 103
use INVX1  INVX1_6
timestamp 1625156677
transform 1 0 4124 0 1 3505
box -2 -3 18 103
use AOI22X1  AOI22X1_3
timestamp 1625156677
transform -1 0 4180 0 1 3505
box -2 -3 42 103
use OAI22X1  OAI22X1_7
timestamp 1625156677
transform -1 0 4220 0 1 3505
box -2 -3 42 103
use INVX1  INVX1_5
timestamp 1625156677
transform -1 0 4236 0 1 3505
box -2 -3 18 103
use CLKBUF1  CLKBUF1_43
timestamp 1625156677
transform -1 0 4308 0 1 3505
box -2 -3 74 103
use AOI21X1  AOI21X1_7
timestamp 1625156677
transform 1 0 4308 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_13
timestamp 1625156677
transform 1 0 4340 0 1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_3
timestamp 1625156677
transform 1 0 4364 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_14
timestamp 1625156677
transform -1 0 4420 0 1 3505
box -2 -3 26 103
use INVX4  INVX4_1
timestamp 1625156677
transform -1 0 4444 0 1 3505
box -2 -3 26 103
use FILL  FILL_35_8_0
timestamp 1625156677
transform 1 0 4444 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_8_1
timestamp 1625156677
transform 1 0 4452 0 1 3505
box -2 -3 10 103
use INVX2  INVX2_3
timestamp 1625156677
transform 1 0 4460 0 1 3505
box -2 -3 18 103
use AOI22X1  AOI22X1_2
timestamp 1625156677
transform -1 0 4516 0 1 3505
box -2 -3 42 103
use OAI22X1  OAI22X1_2
timestamp 1625156677
transform -1 0 4556 0 1 3505
box -2 -3 42 103
use AOI22X1  AOI22X1_1
timestamp 1625156677
transform 1 0 4556 0 1 3505
box -2 -3 42 103
use NAND2X1  NAND2X1_9
timestamp 1625156677
transform 1 0 4596 0 1 3505
box -2 -3 26 103
use INVX2  INVX2_2
timestamp 1625156677
transform -1 0 4636 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_3
timestamp 1625156677
transform 1 0 4636 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1625156677
transform 1 0 4668 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_8
timestamp 1625156677
transform -1 0 4716 0 1 3505
box -2 -3 26 103
use BUFX4  BUFX4_25
timestamp 1625156677
transform 1 0 4716 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_9
timestamp 1625156677
transform 1 0 4748 0 1 3505
box -2 -3 34 103
use BUFX2  BUFX2_83
timestamp 1625156677
transform 1 0 4780 0 1 3505
box -2 -3 26 103
use MUX2X1  MUX2X1_19
timestamp 1625156677
transform -1 0 4852 0 1 3505
box -2 -3 50 103
use OAI22X1  OAI22X1_10
timestamp 1625156677
transform 1 0 4852 0 1 3505
box -2 -3 42 103
use INVX1  INVX1_9
timestamp 1625156677
transform 1 0 4892 0 1 3505
box -2 -3 18 103
use AOI22X1  AOI22X1_5
timestamp 1625156677
transform -1 0 4948 0 1 3505
box -2 -3 42 103
use FILL  FILL_35_9_0
timestamp 1625156677
transform 1 0 4948 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_9_1
timestamp 1625156677
transform 1 0 4956 0 1 3505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_3
timestamp 1625156677
transform 1 0 4964 0 1 3505
box -2 -3 58 103
use MUX2X1  MUX2X1_16
timestamp 1625156677
transform 1 0 5020 0 1 3505
box -2 -3 50 103
use NOR3X1  NOR3X1_16
timestamp 1625156677
transform 1 0 5068 0 1 3505
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1625156677
transform 1 0 5132 0 1 3505
box -2 -3 98 103
use BUFX2  BUFX2_16
timestamp 1625156677
transform 1 0 5228 0 1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_122
timestamp 1625156677
transform -1 0 5276 0 1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_195
timestamp 1625156677
transform 1 0 5276 0 1 3505
box -2 -3 34 103
use FILL  FILL_36_1
timestamp 1625156677
transform 1 0 5308 0 1 3505
box -2 -3 10 103
use XOR2X1  XOR2X1_209
timestamp 1625156677
transform -1 0 60 0 -1 3505
box -2 -3 58 103
use OAI21X1  OAI21X1_397
timestamp 1625156677
transform 1 0 60 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_442
timestamp 1625156677
transform 1 0 92 0 -1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_372
timestamp 1625156677
transform 1 0 116 0 -1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_255
timestamp 1625156677
transform 1 0 148 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_304
timestamp 1625156677
transform 1 0 180 0 -1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_380
timestamp 1625156677
transform 1 0 196 0 -1 3505
box -2 -3 34 103
use INVX2  INVX2_65
timestamp 1625156677
transform 1 0 228 0 -1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_421
timestamp 1625156677
transform 1 0 244 0 -1 3505
box -2 -3 34 103
use NOR3X1  NOR3X1_70
timestamp 1625156677
transform -1 0 340 0 -1 3505
box -2 -3 66 103
use FILL  FILL_34_0_0
timestamp 1625156677
transform 1 0 340 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_0_1
timestamp 1625156677
transform 1 0 348 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_396
timestamp 1625156677
transform 1 0 356 0 -1 3505
box -2 -3 34 103
use AND2X2  AND2X2_124
timestamp 1625156677
transform 1 0 388 0 -1 3505
box -2 -3 34 103
use BUFX2  BUFX2_135
timestamp 1625156677
transform -1 0 444 0 -1 3505
box -2 -3 26 103
use AOI22X1  AOI22X1_15
timestamp 1625156677
transform -1 0 484 0 -1 3505
box -2 -3 42 103
use NAND3X1  NAND3X1_392
timestamp 1625156677
transform 1 0 484 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_331
timestamp 1625156677
transform 1 0 516 0 -1 3505
box -2 -3 18 103
use INVX1  INVX1_333
timestamp 1625156677
transform 1 0 532 0 -1 3505
box -2 -3 18 103
use INVX1  INVX1_337
timestamp 1625156677
transform 1 0 548 0 -1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_472
timestamp 1625156677
transform 1 0 564 0 -1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_272
timestamp 1625156677
transform 1 0 588 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_473
timestamp 1625156677
transform 1 0 612 0 -1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_266
timestamp 1625156677
transform 1 0 636 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_395
timestamp 1625156677
transform 1 0 668 0 -1 3505
box -2 -3 34 103
use XOR2X1  XOR2X1_219
timestamp 1625156677
transform -1 0 756 0 -1 3505
box -2 -3 58 103
use OAI21X1  OAI21X1_416
timestamp 1625156677
transform -1 0 788 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_264
timestamp 1625156677
transform -1 0 812 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_460
timestamp 1625156677
transform -1 0 836 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_468
timestamp 1625156677
transform -1 0 860 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_1_0
timestamp 1625156677
transform 1 0 860 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_1_1
timestamp 1625156677
transform 1 0 868 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_427
timestamp 1625156677
transform 1 0 876 0 -1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_262
timestamp 1625156677
transform 1 0 908 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_322
timestamp 1625156677
transform -1 0 956 0 -1 3505
box -2 -3 18 103
use XOR2X1  XOR2X1_217
timestamp 1625156677
transform 1 0 956 0 -1 3505
box -2 -3 58 103
use AND2X2  AND2X2_127
timestamp 1625156677
transform -1 0 1044 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_459
timestamp 1625156677
transform 1 0 1044 0 -1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_263
timestamp 1625156677
transform -1 0 1092 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_414
timestamp 1625156677
transform 1 0 1092 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_321
timestamp 1625156677
transform -1 0 1140 0 -1 3505
box -2 -3 18 103
use BUFX2  BUFX2_216
timestamp 1625156677
transform -1 0 1164 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_413
timestamp 1625156677
transform 1 0 1164 0 -1 3505
box -2 -3 34 103
use XOR2X1  XOR2X1_216
timestamp 1625156677
transform 1 0 1196 0 -1 3505
box -2 -3 58 103
use XOR2X1  XOR2X1_235
timestamp 1625156677
transform -1 0 1308 0 -1 3505
box -2 -3 58 103
use OAI21X1  OAI21X1_463
timestamp 1625156677
transform 1 0 1308 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_417
timestamp 1625156677
transform 1 0 1340 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_2_0
timestamp 1625156677
transform 1 0 1372 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_2_1
timestamp 1625156677
transform 1 0 1380 0 -1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_512
timestamp 1625156677
transform 1 0 1388 0 -1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_292
timestamp 1625156677
transform -1 0 1436 0 -1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_281
timestamp 1625156677
transform -1 0 1468 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_505
timestamp 1625156677
transform 1 0 1468 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_462
timestamp 1625156677
transform -1 0 1524 0 -1 3505
box -2 -3 34 103
use XOR2X1  XOR2X1_251
timestamp 1625156677
transform 1 0 1524 0 -1 3505
box -2 -3 58 103
use NAND2X1  NAND2X1_507
timestamp 1625156677
transform 1 0 1580 0 -1 3505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_185
timestamp 1625156677
transform -1 0 1660 0 -1 3505
box -2 -3 58 103
use AOI21X1  AOI21X1_280
timestamp 1625156677
transform -1 0 1692 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_293
timestamp 1625156677
transform 1 0 1692 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_468
timestamp 1625156677
transform -1 0 1748 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_419
timestamp 1625156677
transform -1 0 1780 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_452
timestamp 1625156677
transform 1 0 1780 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_361
timestamp 1625156677
transform 1 0 1812 0 -1 3505
box -2 -3 18 103
use NOR2X1  NOR2X1_287
timestamp 1625156677
transform -1 0 1852 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_497
timestamp 1625156677
transform -1 0 1876 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_3_0
timestamp 1625156677
transform 1 0 1876 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_3_1
timestamp 1625156677
transform 1 0 1884 0 -1 3505
box -2 -3 10 103
use AND2X2  AND2X2_135
timestamp 1625156677
transform 1 0 1892 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_289
timestamp 1625156677
transform 1 0 1924 0 -1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_290
timestamp 1625156677
transform -1 0 1972 0 -1 3505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_184
timestamp 1625156677
transform -1 0 2028 0 -1 3505
box -2 -3 58 103
use XOR2X1  XOR2X1_246
timestamp 1625156677
transform 1 0 2028 0 -1 3505
box -2 -3 58 103
use NAND2X1  NAND2X1_524
timestamp 1625156677
transform 1 0 2084 0 -1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_289
timestamp 1625156677
transform 1 0 2108 0 -1 3505
box -2 -3 34 103
use XOR2X1  XOR2X1_260
timestamp 1625156677
transform -1 0 2196 0 -1 3505
box -2 -3 58 103
use OAI21X1  OAI21X1_481
timestamp 1625156677
transform -1 0 2228 0 -1 3505
box -2 -3 34 103
use XOR2X1  XOR2X1_257
timestamp 1625156677
transform 1 0 2228 0 -1 3505
box -2 -3 58 103
use NOR2X1  NOR2X1_304
timestamp 1625156677
transform -1 0 2308 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_526
timestamp 1625156677
transform 1 0 2308 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_487
timestamp 1625156677
transform -1 0 2364 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_305
timestamp 1625156677
transform 1 0 2364 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_4_0
timestamp 1625156677
transform -1 0 2396 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_4_1
timestamp 1625156677
transform -1 0 2404 0 -1 3505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_189
timestamp 1625156677
transform -1 0 2460 0 -1 3505
box -2 -3 58 103
use OAI21X1  OAI21X1_480
timestamp 1625156677
transform -1 0 2492 0 -1 3505
box -2 -3 34 103
use NOR3X1  NOR3X1_77
timestamp 1625156677
transform -1 0 2556 0 -1 3505
box -2 -3 66 103
use NAND3X1  NAND3X1_425
timestamp 1625156677
transform -1 0 2588 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_381
timestamp 1625156677
transform 1 0 2588 0 -1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_476
timestamp 1625156677
transform -1 0 2636 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_502
timestamp 1625156677
transform 1 0 2636 0 -1 3505
box -2 -3 34 103
use BUFX2  BUFX2_225
timestamp 1625156677
transform -1 0 2692 0 -1 3505
box -2 -3 26 103
use BUFX2  BUFX2_224
timestamp 1625156677
transform 1 0 2692 0 -1 3505
box -2 -3 26 103
use INVX1  INVX1_409
timestamp 1625156677
transform 1 0 2716 0 -1 3505
box -2 -3 18 103
use XOR2X1  XOR2X1_253
timestamp 1625156677
transform 1 0 2732 0 -1 3505
box -2 -3 58 103
use XOR2X1  XOR2X1_255
timestamp 1625156677
transform 1 0 2788 0 -1 3505
box -2 -3 58 103
use OAI21X1  OAI21X1_505
timestamp 1625156677
transform -1 0 2876 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_413
timestamp 1625156677
transform 1 0 2876 0 -1 3505
box -2 -3 18 103
use NOR2X1  NOR2X1_317
timestamp 1625156677
transform 1 0 2892 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_5_0
timestamp 1625156677
transform -1 0 2924 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_5_1
timestamp 1625156677
transform -1 0 2932 0 -1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_506
timestamp 1625156677
transform -1 0 2964 0 -1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_296
timestamp 1625156677
transform -1 0 2996 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_496
timestamp 1625156677
transform 1 0 2996 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_438
timestamp 1625156677
transform -1 0 3060 0 -1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_295
timestamp 1625156677
transform 1 0 3060 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_408
timestamp 1625156677
transform -1 0 3108 0 -1 3505
box -2 -3 18 103
use NAND3X1  NAND3X1_439
timestamp 1625156677
transform 1 0 3108 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_401
timestamp 1625156677
transform -1 0 3156 0 -1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_499
timestamp 1625156677
transform -1 0 3188 0 -1 3505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1625156677
transform -1 0 3284 0 -1 3505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1625156677
transform 1 0 3284 0 -1 3505
box -2 -3 98 103
use FILL  FILL_34_6_0
timestamp 1625156677
transform -1 0 3388 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_6_1
timestamp 1625156677
transform -1 0 3396 0 -1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1625156677
transform -1 0 3492 0 -1 3505
box -2 -3 98 103
use BUFX2  BUFX2_136
timestamp 1625156677
transform 1 0 3492 0 -1 3505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1625156677
transform 1 0 3516 0 -1 3505
box -2 -3 98 103
use NOR3X1  NOR3X1_2
timestamp 1625156677
transform 1 0 3612 0 -1 3505
box -2 -3 66 103
use BUFX4  BUFX4_24
timestamp 1625156677
transform -1 0 3708 0 -1 3505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_4
timestamp 1625156677
transform -1 0 3780 0 -1 3505
box -2 -3 74 103
use BUFX2  BUFX2_5
timestamp 1625156677
transform -1 0 3804 0 -1 3505
box -2 -3 26 103
use BUFX2  BUFX2_102
timestamp 1625156677
transform -1 0 3828 0 -1 3505
box -2 -3 26 103
use BUFX4  BUFX4_22
timestamp 1625156677
transform -1 0 3860 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1625156677
transform -1 0 3892 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_7_0
timestamp 1625156677
transform -1 0 3900 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_7_1
timestamp 1625156677
transform -1 0 3908 0 -1 3505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1625156677
transform -1 0 4004 0 -1 3505
box -2 -3 98 103
use NOR3X1  NOR3X1_15
timestamp 1625156677
transform -1 0 4068 0 -1 3505
box -2 -3 66 103
use BUFX2  BUFX2_15
timestamp 1625156677
transform -1 0 4092 0 -1 3505
box -2 -3 26 103
use BUFX4  BUFX4_20
timestamp 1625156677
transform 1 0 4092 0 -1 3505
box -2 -3 34 103
use BUFX4  BUFX4_27
timestamp 1625156677
transform 1 0 4124 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_2
timestamp 1625156677
transform -1 0 4188 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_12
timestamp 1625156677
transform 1 0 4188 0 -1 3505
box -2 -3 26 103
use OAI22X1  OAI22X1_6
timestamp 1625156677
transform -1 0 4252 0 -1 3505
box -2 -3 42 103
use NAND2X1  NAND2X1_11
timestamp 1625156677
transform 1 0 4252 0 -1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_13
timestamp 1625156677
transform -1 0 4300 0 -1 3505
box -2 -3 26 103
use AOI22X1  AOI22X1_7
timestamp 1625156677
transform 1 0 4300 0 -1 3505
box -2 -3 42 103
use INVX2  INVX2_8
timestamp 1625156677
transform -1 0 4356 0 -1 3505
box -2 -3 18 103
use NOR2X1  NOR2X1_11
timestamp 1625156677
transform 1 0 4356 0 -1 3505
box -2 -3 26 103
use OAI22X1  OAI22X1_8
timestamp 1625156677
transform 1 0 4380 0 -1 3505
box -2 -3 42 103
use NOR2X1  NOR2X1_14
timestamp 1625156677
transform 1 0 4420 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_8_0
timestamp 1625156677
transform 1 0 4444 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_8_1
timestamp 1625156677
transform 1 0 4452 0 -1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_19
timestamp 1625156677
transform 1 0 4460 0 -1 3505
box -2 -3 26 103
use OAI22X1  OAI22X1_1
timestamp 1625156677
transform -1 0 4524 0 -1 3505
box -2 -3 42 103
use NOR2X1  NOR2X1_8
timestamp 1625156677
transform 1 0 4524 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_2
timestamp 1625156677
transform -1 0 4572 0 -1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_16
timestamp 1625156677
transform 1 0 4572 0 -1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_9
timestamp 1625156677
transform -1 0 4628 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_18
timestamp 1625156677
transform -1 0 4652 0 -1 3505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_48
timestamp 1625156677
transform 1 0 4652 0 -1 3505
box -2 -3 74 103
use BUFX4  BUFX4_21
timestamp 1625156677
transform -1 0 4756 0 -1 3505
box -2 -3 34 103
use INVX2  INVX2_10
timestamp 1625156677
transform 1 0 4756 0 -1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_7
timestamp 1625156677
transform -1 0 4804 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_6
timestamp 1625156677
transform -1 0 4836 0 -1 3505
box -2 -3 34 103
use INVX2  INVX2_6
timestamp 1625156677
transform 1 0 4836 0 -1 3505
box -2 -3 18 103
use AOI22X1  AOI22X1_6
timestamp 1625156677
transform 1 0 4852 0 -1 3505
box -2 -3 42 103
use NAND2X1  NAND2X1_15
timestamp 1625156677
transform -1 0 4916 0 -1 3505
box -2 -3 26 103
use INVX2  INVX2_7
timestamp 1625156677
transform 1 0 4916 0 -1 3505
box -2 -3 18 103
use FILL  FILL_34_9_0
timestamp 1625156677
transform 1 0 4932 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_9_1
timestamp 1625156677
transform 1 0 4940 0 -1 3505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_2
timestamp 1625156677
transform 1 0 4948 0 -1 3505
box -2 -3 58 103
use MUX2X1  MUX2X1_12
timestamp 1625156677
transform 1 0 5004 0 -1 3505
box -2 -3 50 103
use NOR3X1  NOR3X1_12
timestamp 1625156677
transform 1 0 5052 0 -1 3505
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1625156677
transform 1 0 5116 0 -1 3505
box -2 -3 98 103
use BUFX2  BUFX2_12
timestamp 1625156677
transform 1 0 5212 0 -1 3505
box -2 -3 26 103
use BUFX2  BUFX2_120
timestamp 1625156677
transform -1 0 5260 0 -1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_191
timestamp 1625156677
transform 1 0 5260 0 -1 3505
box -2 -3 34 103
use FILL  FILL_35_1
timestamp 1625156677
transform -1 0 5300 0 -1 3505
box -2 -3 10 103
use FILL  FILL_35_2
timestamp 1625156677
transform -1 0 5308 0 -1 3505
box -2 -3 10 103
use FILL  FILL_35_3
timestamp 1625156677
transform -1 0 5316 0 -1 3505
box -2 -3 10 103
use NOR2X1  NOR2X1_255
timestamp 1625156677
transform 1 0 4 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_400
timestamp 1625156677
transform 1 0 28 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_444
timestamp 1625156677
transform -1 0 84 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_305
timestamp 1625156677
transform -1 0 100 0 1 3305
box -2 -3 18 103
use INVX1  INVX1_306
timestamp 1625156677
transform -1 0 116 0 1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_373
timestamp 1625156677
transform 1 0 116 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_443
timestamp 1625156677
transform -1 0 172 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_313
timestamp 1625156677
transform -1 0 188 0 1 3305
box -2 -3 18 103
use AOI21X1  AOI21X1_256
timestamp 1625156677
transform 1 0 188 0 1 3305
box -2 -3 34 103
use NOR3X1  NOR3X1_69
timestamp 1625156677
transform -1 0 284 0 1 3305
box -2 -3 66 103
use OAI21X1  OAI21X1_398
timestamp 1625156677
transform -1 0 316 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_254
timestamp 1625156677
transform 1 0 316 0 1 3305
box -2 -3 26 103
use FILL  FILL_33_0_0
timestamp 1625156677
transform -1 0 348 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_0_1
timestamp 1625156677
transform -1 0 356 0 1 3305
box -2 -3 10 103
use NOR2X1  NOR2X1_253
timestamp 1625156677
transform -1 0 380 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_399
timestamp 1625156677
transform -1 0 412 0 1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_371
timestamp 1625156677
transform 1 0 412 0 1 3305
box -2 -3 34 103
use AND2X2  AND2X2_123
timestamp 1625156677
transform -1 0 476 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_440
timestamp 1625156677
transform -1 0 500 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_302
timestamp 1625156677
transform -1 0 516 0 1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_391
timestamp 1625156677
transform 1 0 516 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_465
timestamp 1625156677
transform -1 0 572 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_466
timestamp 1625156677
transform -1 0 596 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_330
timestamp 1625156677
transform 1 0 596 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_425
timestamp 1625156677
transform -1 0 644 0 1 3305
box -2 -3 34 103
use BUFX2  BUFX2_207
timestamp 1625156677
transform 1 0 644 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_335
timestamp 1625156677
transform -1 0 684 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_431
timestamp 1625156677
transform 1 0 684 0 1 3305
box -2 -3 34 103
use AND2X2  AND2X2_129
timestamp 1625156677
transform 1 0 716 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_338
timestamp 1625156677
transform 1 0 748 0 1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_396
timestamp 1625156677
transform 1 0 764 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_475
timestamp 1625156677
transform 1 0 796 0 1 3305
box -2 -3 26 103
use XOR2X1  XOR2X1_218
timestamp 1625156677
transform -1 0 876 0 1 3305
box -2 -3 58 103
use FILL  FILL_33_1_0
timestamp 1625156677
transform 1 0 876 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_1_1
timestamp 1625156677
transform 1 0 884 0 1 3305
box -2 -3 10 103
use BUFX2  BUFX2_211
timestamp 1625156677
transform 1 0 892 0 1 3305
box -2 -3 26 103
use XOR2X1  XOR2X1_241
timestamp 1625156677
transform 1 0 916 0 1 3305
box -2 -3 58 103
use NAND2X1  NAND2X1_492
timestamp 1625156677
transform 1 0 972 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_354
timestamp 1625156677
transform -1 0 1012 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_450
timestamp 1625156677
transform -1 0 1044 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_357
timestamp 1625156677
transform 1 0 1044 0 1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_409
timestamp 1625156677
transform 1 0 1060 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_494
timestamp 1625156677
transform 1 0 1092 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_274
timestamp 1625156677
transform -1 0 1148 0 1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_408
timestamp 1625156677
transform -1 0 1180 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_356
timestamp 1625156677
transform -1 0 1196 0 1 3305
box -2 -3 18 103
use INVX1  INVX1_355
timestamp 1625156677
transform 1 0 1196 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_448
timestamp 1625156677
transform -1 0 1244 0 1 3305
box -2 -3 34 103
use AND2X2  AND2X2_133
timestamp 1625156677
transform 1 0 1244 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_297
timestamp 1625156677
transform -1 0 1300 0 1 3305
box -2 -3 26 103
use XOR2X1  XOR2X1_250
timestamp 1625156677
transform -1 0 1356 0 1 3305
box -2 -3 58 103
use FILL  FILL_33_2_0
timestamp 1625156677
transform 1 0 1356 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_2_1
timestamp 1625156677
transform 1 0 1364 0 1 3305
box -2 -3 10 103
use XOR2X1  XOR2X1_248
timestamp 1625156677
transform 1 0 1372 0 1 3305
box -2 -3 58 103
use NOR2X1  NOR2X1_294
timestamp 1625156677
transform 1 0 1428 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_503
timestamp 1625156677
transform -1 0 1476 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_464
timestamp 1625156677
transform 1 0 1476 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_368
timestamp 1625156677
transform 1 0 1508 0 1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_504
timestamp 1625156677
transform 1 0 1524 0 1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_418
timestamp 1625156677
transform 1 0 1548 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_369
timestamp 1625156677
transform -1 0 1596 0 1 3305
box -2 -3 18 103
use AOI22X1  AOI22X1_17
timestamp 1625156677
transform -1 0 1636 0 1 3305
box -2 -3 42 103
use INVX1  INVX1_371
timestamp 1625156677
transform 1 0 1636 0 1 3305
box -2 -3 18 103
use XOR2X1  XOR2X1_249
timestamp 1625156677
transform -1 0 1708 0 1 3305
box -2 -3 58 103
use BUFX2  BUFX2_222
timestamp 1625156677
transform 1 0 1708 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_282
timestamp 1625156677
transform -1 0 1764 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_375
timestamp 1625156677
transform -1 0 1780 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_467
timestamp 1625156677
transform 1 0 1780 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_374
timestamp 1625156677
transform -1 0 1828 0 1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_421
timestamp 1625156677
transform 1 0 1828 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_359
timestamp 1625156677
transform 1 0 1860 0 1 3305
box -2 -3 18 103
use FILL  FILL_33_3_0
timestamp 1625156677
transform 1 0 1876 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_3_1
timestamp 1625156677
transform 1 0 1884 0 1 3305
box -2 -3 10 103
use AND2X2  AND2X2_137
timestamp 1625156677
transform 1 0 1892 0 1 3305
box -2 -3 34 103
use BUFX2  BUFX2_221
timestamp 1625156677
transform 1 0 1924 0 1 3305
box -2 -3 26 103
use XOR2X1  XOR2X1_245
timestamp 1625156677
transform -1 0 2004 0 1 3305
box -2 -3 58 103
use NOR2X1  NOR2X1_307
timestamp 1625156677
transform -1 0 2028 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_527
timestamp 1625156677
transform -1 0 2052 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_482
timestamp 1625156677
transform 1 0 2052 0 1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_430
timestamp 1625156677
transform -1 0 2116 0 1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_431
timestamp 1625156677
transform 1 0 2116 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_388
timestamp 1625156677
transform -1 0 2164 0 1 3305
box -2 -3 18 103
use AOI22X1  AOI22X1_18
timestamp 1625156677
transform 1 0 2164 0 1 3305
box -2 -3 42 103
use XOR2X1  XOR2X1_267
timestamp 1625156677
transform -1 0 2260 0 1 3305
box -2 -3 58 103
use AND2X2  AND2X2_141
timestamp 1625156677
transform -1 0 2292 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_394
timestamp 1625156677
transform 1 0 2292 0 1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_434
timestamp 1625156677
transform 1 0 2308 0 1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_290
timestamp 1625156677
transform 1 0 2340 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_393
timestamp 1625156677
transform 1 0 2372 0 1 3305
box -2 -3 18 103
use FILL  FILL_33_4_0
timestamp 1625156677
transform -1 0 2396 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_4_1
timestamp 1625156677
transform -1 0 2404 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_486
timestamp 1625156677
transform -1 0 2436 0 1 3305
box -2 -3 34 103
use XOR2X1  XOR2X1_265
timestamp 1625156677
transform 1 0 2436 0 1 3305
box -2 -3 58 103
use AOI21X1  AOI21X1_288
timestamp 1625156677
transform -1 0 2524 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_389
timestamp 1625156677
transform 1 0 2524 0 1 3305
box -2 -3 18 103
use AOI21X1  AOI21X1_287
timestamp 1625156677
transform -1 0 2572 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_518
timestamp 1625156677
transform 1 0 2572 0 1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_424
timestamp 1625156677
transform 1 0 2596 0 1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_432
timestamp 1625156677
transform -1 0 2660 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_521
timestamp 1625156677
transform 1 0 2660 0 1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_301
timestamp 1625156677
transform 1 0 2684 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_380
timestamp 1625156677
transform -1 0 2724 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_474
timestamp 1625156677
transform -1 0 2756 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_302
timestamp 1625156677
transform -1 0 2780 0 1 3305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_188
timestamp 1625156677
transform -1 0 2836 0 1 3305
box -2 -3 58 103
use BUFX2  BUFX2_226
timestamp 1625156677
transform 1 0 2836 0 1 3305
box -2 -3 26 103
use BUFX2  BUFX2_230
timestamp 1625156677
transform 1 0 2860 0 1 3305
box -2 -3 26 103
use FILL  FILL_33_5_0
timestamp 1625156677
transform 1 0 2884 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_5_1
timestamp 1625156677
transform 1 0 2892 0 1 3305
box -2 -3 10 103
use XOR2X1  XOR2X1_252
timestamp 1625156677
transform 1 0 2900 0 1 3305
box -2 -3 58 103
use NAND3X1  NAND3X1_447
timestamp 1625156677
transform 1 0 2956 0 1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_298
timestamp 1625156677
transform 1 0 2988 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_412
timestamp 1625156677
transform 1 0 3020 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_490
timestamp 1625156677
transform 1 0 3036 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_311
timestamp 1625156677
transform 1 0 3068 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_535
timestamp 1625156677
transform -1 0 3116 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_397
timestamp 1625156677
transform 1 0 3116 0 1 3305
box -2 -3 18 103
use AND2X2  AND2X2_143
timestamp 1625156677
transform 1 0 3132 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_494
timestamp 1625156677
transform 1 0 3164 0 1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_445
timestamp 1625156677
transform -1 0 3228 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_313
timestamp 1625156677
transform 1 0 3228 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_399
timestamp 1625156677
transform -1 0 3268 0 1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_540
timestamp 1625156677
transform 1 0 3268 0 1 3305
box -2 -3 26 103
use NOR3X1  NOR3X1_79
timestamp 1625156677
transform 1 0 3292 0 1 3305
box -2 -3 66 103
use BUFX2  BUFX2_26
timestamp 1625156677
transform 1 0 3356 0 1 3305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_250
timestamp 1625156677
transform -1 0 3436 0 1 3305
box -2 -3 58 103
use FILL  FILL_33_6_0
timestamp 1625156677
transform -1 0 3444 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_6_1
timestamp 1625156677
transform -1 0 3452 0 1 3305
box -2 -3 10 103
use INVX1  INVX1_589
timestamp 1625156677
transform -1 0 3468 0 1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_702
timestamp 1625156677
transform 1 0 3468 0 1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_444
timestamp 1625156677
transform -1 0 3516 0 1 3305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_249
timestamp 1625156677
transform -1 0 3572 0 1 3305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1625156677
transform -1 0 3668 0 1 3305
box -2 -3 98 103
use MUX2X1  MUX2X1_2
timestamp 1625156677
transform -1 0 3716 0 1 3305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1625156677
transform -1 0 3812 0 1 3305
box -2 -3 98 103
use MUX2X1  MUX2X1_5
timestamp 1625156677
transform 1 0 3812 0 1 3305
box -2 -3 50 103
use BUFX4  BUFX4_11
timestamp 1625156677
transform -1 0 3892 0 1 3305
box -2 -3 34 103
use NOR3X1  NOR3X1_5
timestamp 1625156677
transform 1 0 3892 0 1 3305
box -2 -3 66 103
use FILL  FILL_33_7_0
timestamp 1625156677
transform -1 0 3964 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_7_1
timestamp 1625156677
transform -1 0 3972 0 1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1625156677
transform -1 0 4068 0 1 3305
box -2 -3 98 103
use MUX2X1  MUX2X1_15
timestamp 1625156677
transform -1 0 4116 0 1 3305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1625156677
transform -1 0 4212 0 1 3305
box -2 -3 98 103
use INVX2  INVX2_9
timestamp 1625156677
transform 1 0 4212 0 1 3305
box -2 -3 18 103
use NOR2X1  NOR2X1_7
timestamp 1625156677
transform -1 0 4252 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1625156677
transform 1 0 4252 0 1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_1
timestamp 1625156677
transform -1 0 4372 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_1
timestamp 1625156677
transform 1 0 4372 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_5
timestamp 1625156677
transform 1 0 4396 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_8_0
timestamp 1625156677
transform -1 0 4436 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_8_1
timestamp 1625156677
transform -1 0 4444 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_4
timestamp 1625156677
transform -1 0 4476 0 1 3305
box -2 -3 34 103
use BUFX2  BUFX2_81
timestamp 1625156677
transform 1 0 4476 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1625156677
transform -1 0 4596 0 1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_10
timestamp 1625156677
transform 1 0 4596 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_4
timestamp 1625156677
transform -1 0 4652 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_7
timestamp 1625156677
transform 1 0 4652 0 1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_10
timestamp 1625156677
transform 1 0 4676 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1625156677
transform 1 0 4700 0 1 3305
box -2 -3 98 103
use NAND3X1  NAND3X1_4
timestamp 1625156677
transform -1 0 4828 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_15
timestamp 1625156677
transform 1 0 4828 0 1 3305
box -2 -3 26 103
use OAI22X1  OAI22X1_5
timestamp 1625156677
transform 1 0 4852 0 1 3305
box -2 -3 42 103
use NAND2X1  NAND2X1_6
timestamp 1625156677
transform 1 0 4892 0 1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_4
timestamp 1625156677
transform -1 0 4940 0 1 3305
box -2 -3 26 103
use FILL  FILL_33_9_0
timestamp 1625156677
transform -1 0 4948 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_9_1
timestamp 1625156677
transform -1 0 4956 0 1 3305
box -2 -3 10 103
use AOI21X1  AOI21X1_2
timestamp 1625156677
transform -1 0 4988 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_5
timestamp 1625156677
transform -1 0 5012 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_2
timestamp 1625156677
transform -1 0 5044 0 1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_1
timestamp 1625156677
transform -1 0 5076 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1625156677
transform 1 0 5076 0 1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_1
timestamp 1625156677
transform 1 0 5100 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_9
timestamp 1625156677
transform -1 0 5156 0 1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1625156677
transform 1 0 5156 0 1 3305
box -2 -3 98 103
use NAND2X1  NAND2X1_219
timestamp 1625156677
transform 1 0 5252 0 1 3305
box -2 -3 26 103
use AND2X2  AND2X2_64
timestamp 1625156677
transform -1 0 5308 0 1 3305
box -2 -3 34 103
use FILL  FILL_34_1
timestamp 1625156677
transform 1 0 5308 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_401
timestamp 1625156677
transform 1 0 4 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_253
timestamp 1625156677
transform 1 0 36 0 -1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_374
timestamp 1625156677
transform 1 0 68 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_404
timestamp 1625156677
transform -1 0 132 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_257
timestamp 1625156677
transform 1 0 132 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_411
timestamp 1625156677
transform 1 0 156 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_445
timestamp 1625156677
transform -1 0 212 0 -1 3305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_172
timestamp 1625156677
transform -1 0 268 0 -1 3305
box -2 -3 58 103
use BUFX2  BUFX2_214
timestamp 1625156677
transform 1 0 268 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_213
timestamp 1625156677
transform -1 0 316 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_395
timestamp 1625156677
transform 1 0 316 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_0_0
timestamp 1625156677
transform 1 0 348 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_0_1
timestamp 1625156677
transform 1 0 356 0 -1 3305
box -2 -3 10 103
use AND2X2  AND2X2_125
timestamp 1625156677
transform 1 0 364 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_251
timestamp 1625156677
transform -1 0 420 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_212
timestamp 1625156677
transform 1 0 420 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_270
timestamp 1625156677
transform 1 0 444 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_426
timestamp 1625156677
transform 1 0 468 0 -1 3305
box -2 -3 34 103
use XOR2X1  XOR2X1_231
timestamp 1625156677
transform 1 0 500 0 -1 3305
box -2 -3 58 103
use NOR2X1  NOR2X1_283
timestamp 1625156677
transform -1 0 580 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_447
timestamp 1625156677
transform 1 0 580 0 -1 3305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_183
timestamp 1625156677
transform -1 0 668 0 -1 3305
box -2 -3 58 103
use NAND2X1  NAND2X1_490
timestamp 1625156677
transform 1 0 668 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_489
timestamp 1625156677
transform -1 0 716 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_353
timestamp 1625156677
transform -1 0 732 0 -1 3305
box -2 -3 18 103
use XOR2X1  XOR2X1_240
timestamp 1625156677
transform 1 0 732 0 -1 3305
box -2 -3 58 103
use NAND2X1  NAND2X1_491
timestamp 1625156677
transform -1 0 812 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_284
timestamp 1625156677
transform -1 0 836 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_486
timestamp 1625156677
transform 1 0 836 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_1_0
timestamp 1625156677
transform 1 0 860 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_1_1
timestamp 1625156677
transform 1 0 868 0 -1 3305
box -2 -3 10 103
use AOI21X1  AOI21X1_273
timestamp 1625156677
transform 1 0 876 0 -1 3305
box -2 -3 34 103
use XOR2X1  XOR2X1_242
timestamp 1625156677
transform -1 0 964 0 -1 3305
box -2 -3 58 103
use NAND2X1  NAND2X1_493
timestamp 1625156677
transform -1 0 988 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_443
timestamp 1625156677
transform -1 0 1020 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_488
timestamp 1625156677
transform 1 0 1020 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_449
timestamp 1625156677
transform -1 0 1076 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_281
timestamp 1625156677
transform 1 0 1076 0 -1 3305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_181
timestamp 1625156677
transform 1 0 1100 0 -1 3305
box -2 -3 58 103
use NOR3X1  NOR3X1_73
timestamp 1625156677
transform -1 0 1220 0 -1 3305
box -2 -3 66 103
use OAI21X1  OAI21X1_442
timestamp 1625156677
transform 1 0 1220 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_272
timestamp 1625156677
transform -1 0 1284 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_436
timestamp 1625156677
transform 1 0 1284 0 -1 3305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_180
timestamp 1625156677
transform 1 0 1316 0 -1 3305
box -2 -3 58 103
use FILL  FILL_32_2_0
timestamp 1625156677
transform 1 0 1372 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_2_1
timestamp 1625156677
transform 1 0 1380 0 -1 3305
box -2 -3 10 103
use XNOR2X1  XNOR2X1_186
timestamp 1625156677
transform 1 0 1388 0 -1 3305
box -2 -3 58 103
use NOR2X1  NOR2X1_278
timestamp 1625156677
transform 1 0 1444 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_295
timestamp 1625156677
transform 1 0 1468 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_508
timestamp 1625156677
transform -1 0 1516 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_372
timestamp 1625156677
transform -1 0 1532 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_466
timestamp 1625156677
transform 1 0 1532 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_509
timestamp 1625156677
transform -1 0 1588 0 -1 3305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_187
timestamp 1625156677
transform -1 0 1644 0 -1 3305
box -2 -3 58 103
use NAND2X1  NAND2X1_510
timestamp 1625156677
transform 1 0 1644 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_296
timestamp 1625156677
transform -1 0 1692 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_511
timestamp 1625156677
transform 1 0 1692 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_373
timestamp 1625156677
transform 1 0 1716 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_469
timestamp 1625156677
transform 1 0 1732 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_376
timestamp 1625156677
transform 1 0 1764 0 -1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_422
timestamp 1625156677
transform 1 0 1780 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_309
timestamp 1625156677
transform -1 0 1836 0 -1 3305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_190
timestamp 1625156677
transform -1 0 1892 0 -1 3305
box -2 -3 58 103
use FILL  FILL_32_3_0
timestamp 1625156677
transform -1 0 1900 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_3_1
timestamp 1625156677
transform -1 0 1908 0 -1 3305
box -2 -3 10 103
use BUFX2  BUFX2_229
timestamp 1625156677
transform -1 0 1932 0 -1 3305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_191
timestamp 1625156677
transform 1 0 1932 0 -1 3305
box -2 -3 58 103
use OAI21X1  OAI21X1_485
timestamp 1625156677
transform 1 0 1988 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_528
timestamp 1625156677
transform 1 0 2020 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_391
timestamp 1625156677
transform -1 0 2060 0 -1 3305
box -2 -3 18 103
use NOR2X1  NOR2X1_306
timestamp 1625156677
transform -1 0 2084 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_522
timestamp 1625156677
transform -1 0 2108 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_483
timestamp 1625156677
transform 1 0 2108 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_387
timestamp 1625156677
transform 1 0 2140 0 -1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_523
timestamp 1625156677
transform 1 0 2156 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_390
timestamp 1625156677
transform 1 0 2180 0 -1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_529
timestamp 1625156677
transform 1 0 2196 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_308
timestamp 1625156677
transform 1 0 2220 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_530
timestamp 1625156677
transform 1 0 2244 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_392
timestamp 1625156677
transform 1 0 2268 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_488
timestamp 1625156677
transform -1 0 2316 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_395
timestamp 1625156677
transform 1 0 2316 0 -1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_435
timestamp 1625156677
transform 1 0 2332 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_473
timestamp 1625156677
transform 1 0 2364 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_4_0
timestamp 1625156677
transform 1 0 2396 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_4_1
timestamp 1625156677
transform 1 0 2404 0 -1 3305
box -2 -3 10 103
use NOR2X1  NOR2X1_300
timestamp 1625156677
transform 1 0 2412 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_484
timestamp 1625156677
transform 1 0 2436 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_379
timestamp 1625156677
transform -1 0 2484 0 -1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_517
timestamp 1625156677
transform 1 0 2484 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_525
timestamp 1625156677
transform 1 0 2508 0 -1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_286
timestamp 1625156677
transform 1 0 2532 0 -1 3305
box -2 -3 34 103
use INVX2  INVX2_69
timestamp 1625156677
transform 1 0 2564 0 -1 3305
box -2 -3 18 103
use NOR3X1  NOR3X1_78
timestamp 1625156677
transform -1 0 2644 0 -1 3305
box -2 -3 66 103
use OAI21X1  OAI21X1_475
timestamp 1625156677
transform -1 0 2676 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_472
timestamp 1625156677
transform 1 0 2676 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_320
timestamp 1625156677
transform -1 0 2732 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_548
timestamp 1625156677
transform 1 0 2732 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_549
timestamp 1625156677
transform 1 0 2756 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_411
timestamp 1625156677
transform -1 0 2796 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_507
timestamp 1625156677
transform -1 0 2828 0 -1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_448
timestamp 1625156677
transform 1 0 2828 0 -1 3305
box -2 -3 34 103
use AND2X2  AND2X2_145
timestamp 1625156677
transform 1 0 2860 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_310
timestamp 1625156677
transform -1 0 2916 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_5_0
timestamp 1625156677
transform -1 0 2924 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_5_1
timestamp 1625156677
transform -1 0 2932 0 -1 3305
box -2 -3 10 103
use NAND2X1  NAND2X1_533
timestamp 1625156677
transform -1 0 2956 0 -1 3305
box -2 -3 26 103
use AND2X2  AND2X2_142
timestamp 1625156677
transform 1 0 2956 0 -1 3305
box -2 -3 34 103
use NOR3X1  NOR3X1_80
timestamp 1625156677
transform -1 0 3052 0 -1 3305
box -2 -3 66 103
use INVX2  INVX2_70
timestamp 1625156677
transform 1 0 3052 0 -1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_436
timestamp 1625156677
transform 1 0 3068 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_491
timestamp 1625156677
transform 1 0 3100 0 -1 3305
box -2 -3 34 103
use AND2X2  AND2X2_144
timestamp 1625156677
transform 1 0 3132 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_294
timestamp 1625156677
transform -1 0 3196 0 -1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_437
timestamp 1625156677
transform -1 0 3228 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_537
timestamp 1625156677
transform 1 0 3228 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_314
timestamp 1625156677
transform -1 0 3276 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_493
timestamp 1625156677
transform -1 0 3308 0 -1 3305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_192
timestamp 1625156677
transform -1 0 3364 0 -1 3305
box -2 -3 58 103
use BUFX2  BUFX2_232
timestamp 1625156677
transform -1 0 3388 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_703
timestamp 1625156677
transform 1 0 3388 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_6_0
timestamp 1625156677
transform -1 0 3420 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_6_1
timestamp 1625156677
transform -1 0 3428 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_634
timestamp 1625156677
transform -1 0 3460 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_633
timestamp 1625156677
transform -1 0 3492 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_701
timestamp 1625156677
transform -1 0 3516 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1625156677
transform 1 0 3516 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1625156677
transform 1 0 3612 0 -1 3305
box -2 -3 98 103
use MUX2X1  MUX2X1_3
timestamp 1625156677
transform 1 0 3708 0 -1 3305
box -2 -3 50 103
use NOR3X1  NOR3X1_3
timestamp 1625156677
transform 1 0 3756 0 -1 3305
box -2 -3 66 103
use BUFX2  BUFX2_108
timestamp 1625156677
transform -1 0 3844 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1625156677
transform -1 0 3940 0 -1 3305
box -2 -3 98 103
use FILL  FILL_32_7_0
timestamp 1625156677
transform 1 0 3940 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_7_1
timestamp 1625156677
transform 1 0 3948 0 -1 3305
box -2 -3 10 103
use BUFX4  BUFX4_26
timestamp 1625156677
transform 1 0 3956 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_17
timestamp 1625156677
transform 1 0 3988 0 -1 3305
box -2 -3 26 103
use BUFX4  BUFX4_18
timestamp 1625156677
transform -1 0 4044 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1625156677
transform -1 0 4140 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1625156677
transform 1 0 4140 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1625156677
transform 1 0 4236 0 -1 3305
box -2 -3 98 103
use XOR2X1  XOR2X1_1
timestamp 1625156677
transform -1 0 4388 0 -1 3305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_1
timestamp 1625156677
transform -1 0 4444 0 -1 3305
box -2 -3 58 103
use FILL  FILL_32_8_0
timestamp 1625156677
transform -1 0 4452 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_8_1
timestamp 1625156677
transform -1 0 4460 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_1
timestamp 1625156677
transform -1 0 4492 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_1
timestamp 1625156677
transform -1 0 4508 0 -1 3305
box -2 -3 18 103
use INVX1  INVX1_2
timestamp 1625156677
transform 1 0 4508 0 -1 3305
box -2 -3 18 103
use AOI21X1  AOI21X1_3
timestamp 1625156677
transform 1 0 4524 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_2
timestamp 1625156677
transform -1 0 4580 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1625156677
transform 1 0 4580 0 -1 3305
box -2 -3 98 103
use AOI21X1  AOI21X1_5
timestamp 1625156677
transform 1 0 4676 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_10
timestamp 1625156677
transform 1 0 4708 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_10
timestamp 1625156677
transform 1 0 4740 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_19
timestamp 1625156677
transform 1 0 4772 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_10
timestamp 1625156677
transform 1 0 4804 0 -1 3305
box -2 -3 18 103
use AOI21X1  AOI21X1_8
timestamp 1625156677
transform 1 0 4820 0 -1 3305
box -2 -3 34 103
use AND2X2  AND2X2_1
timestamp 1625156677
transform -1 0 4884 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_6
timestamp 1625156677
transform -1 0 4916 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_17
timestamp 1625156677
transform 1 0 4916 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_12
timestamp 1625156677
transform 1 0 4940 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_9_0
timestamp 1625156677
transform 1 0 4964 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_9_1
timestamp 1625156677
transform 1 0 4972 0 -1 3305
box -2 -3 10 103
use NAND2X1  NAND2X1_16
timestamp 1625156677
transform 1 0 4980 0 -1 3305
box -2 -3 26 103
use INVX2  INVX2_5
timestamp 1625156677
transform 1 0 5004 0 -1 3305
box -2 -3 18 103
use NOR2X1  NOR2X1_3
timestamp 1625156677
transform 1 0 5020 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_5
timestamp 1625156677
transform -1 0 5068 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_4
timestamp 1625156677
transform -1 0 5092 0 -1 3305
box -2 -3 26 103
use OAI22X1  OAI22X1_4
timestamp 1625156677
transform -1 0 5132 0 -1 3305
box -2 -3 42 103
use INVX1  INVX1_3
timestamp 1625156677
transform 1 0 5132 0 -1 3305
box -2 -3 18 103
use INVX1  INVX1_4
timestamp 1625156677
transform 1 0 5148 0 -1 3305
box -2 -3 18 103
use OAI22X1  OAI22X1_3
timestamp 1625156677
transform 1 0 5164 0 -1 3305
box -2 -3 42 103
use INVX2  INVX2_4
timestamp 1625156677
transform -1 0 5220 0 -1 3305
box -2 -3 18 103
use BUFX2  BUFX2_114
timestamp 1625156677
transform -1 0 5244 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_62
timestamp 1625156677
transform -1 0 5268 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_120
timestamp 1625156677
transform -1 0 5292 0 -1 3305
box -2 -3 26 103
use FILL  FILL_33_1
timestamp 1625156677
transform -1 0 5300 0 -1 3305
box -2 -3 10 103
use FILL  FILL_33_2
timestamp 1625156677
transform -1 0 5308 0 -1 3305
box -2 -3 10 103
use FILL  FILL_33_3
timestamp 1625156677
transform -1 0 5316 0 -1 3305
box -2 -3 10 103
use INVX1  INVX1_307
timestamp 1625156677
transform -1 0 20 0 1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_377
timestamp 1625156677
transform -1 0 52 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_251
timestamp 1625156677
transform -1 0 84 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_256
timestamp 1625156677
transform 1 0 84 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_405
timestamp 1625156677
transform -1 0 140 0 1 3105
box -2 -3 34 103
use XOR2X1  XOR2X1_224
timestamp 1625156677
transform 1 0 140 0 1 3105
box -2 -3 58 103
use NAND2X1  NAND2X1_450
timestamp 1625156677
transform 1 0 196 0 1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_173
timestamp 1625156677
transform -1 0 276 0 1 3105
box -2 -3 58 103
use OAI21X1  OAI21X1_410
timestamp 1625156677
transform 1 0 276 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_318
timestamp 1625156677
transform 1 0 308 0 1 3105
box -2 -3 18 103
use INVX1  INVX1_317
timestamp 1625156677
transform -1 0 340 0 1 3105
box -2 -3 18 103
use FILL  FILL_31_0_0
timestamp 1625156677
transform -1 0 348 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_0_1
timestamp 1625156677
transform -1 0 356 0 1 3105
box -2 -3 10 103
use NAND3X1  NAND3X1_382
timestamp 1625156677
transform -1 0 388 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_258
timestamp 1625156677
transform 1 0 388 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_454
timestamp 1625156677
transform 1 0 420 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_316
timestamp 1625156677
transform -1 0 460 0 1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_383
timestamp 1625156677
transform -1 0 492 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_319
timestamp 1625156677
transform -1 0 508 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_456
timestamp 1625156677
transform 1 0 508 0 1 3105
box -2 -3 26 103
use BUFX2  BUFX2_208
timestamp 1625156677
transform 1 0 532 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_439
timestamp 1625156677
transform -1 0 580 0 1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_229
timestamp 1625156677
transform 1 0 580 0 1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_232
timestamp 1625156677
transform 1 0 636 0 1 3105
box -2 -3 58 103
use NOR2X1  NOR2X1_285
timestamp 1625156677
transform -1 0 716 0 1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_182
timestamp 1625156677
transform 1 0 716 0 1 3105
box -2 -3 58 103
use BUFX2  BUFX2_210
timestamp 1625156677
transform 1 0 772 0 1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_226
timestamp 1625156677
transform 1 0 796 0 1 3105
box -2 -3 58 103
use FILL  FILL_31_1_0
timestamp 1625156677
transform -1 0 860 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_1_1
timestamp 1625156677
transform -1 0 868 0 1 3105
box -2 -3 10 103
use INVX1  INVX1_352
timestamp 1625156677
transform -1 0 884 0 1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_404
timestamp 1625156677
transform -1 0 916 0 1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_405
timestamp 1625156677
transform 1 0 916 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_350
timestamp 1625156677
transform -1 0 964 0 1 3105
box -2 -3 18 103
use AOI22X1  AOI22X1_16
timestamp 1625156677
transform 1 0 964 0 1 3105
box -2 -3 42 103
use XOR2X1  XOR2X1_227
timestamp 1625156677
transform 1 0 1004 0 1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_228
timestamp 1625156677
transform 1 0 1060 0 1 3105
box -2 -3 58 103
use NOR2X1  NOR2X1_280
timestamp 1625156677
transform 1 0 1116 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_267
timestamp 1625156677
transform -1 0 1172 0 1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_403
timestamp 1625156677
transform 1 0 1172 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_345
timestamp 1625156677
transform -1 0 1220 0 1 3105
box -2 -3 18 103
use AOI21X1  AOI21X1_269
timestamp 1625156677
transform 1 0 1220 0 1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_400
timestamp 1625156677
transform 1 0 1252 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_344
timestamp 1625156677
transform -1 0 1300 0 1 3105
box -2 -3 18 103
use INVX1  INVX1_351
timestamp 1625156677
transform 1 0 1300 0 1 3105
box -2 -3 18 103
use AOI21X1  AOI21X1_271
timestamp 1625156677
transform -1 0 1348 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_483
timestamp 1625156677
transform -1 0 1372 0 1 3105
box -2 -3 26 103
use FILL  FILL_31_2_0
timestamp 1625156677
transform 1 0 1372 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_2_1
timestamp 1625156677
transform 1 0 1380 0 1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_480
timestamp 1625156677
transform 1 0 1388 0 1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_398
timestamp 1625156677
transform 1 0 1412 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_342
timestamp 1625156677
transform 1 0 1444 0 1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_406
timestamp 1625156677
transform 1 0 1460 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_277
timestamp 1625156677
transform -1 0 1516 0 1 3105
box -2 -3 26 103
use INVX2  INVX2_67
timestamp 1625156677
transform -1 0 1532 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_437
timestamp 1625156677
transform -1 0 1564 0 1 3105
box -2 -3 34 103
use NOR3X1  NOR3X1_74
timestamp 1625156677
transform 1 0 1564 0 1 3105
box -2 -3 66 103
use OAI21X1  OAI21X1_434
timestamp 1625156677
transform 1 0 1628 0 1 3105
box -2 -3 34 103
use AND2X2  AND2X2_132
timestamp 1625156677
transform 1 0 1660 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_274
timestamp 1625156677
transform -1 0 1716 0 1 3105
box -2 -3 26 103
use AND2X2  AND2X2_130
timestamp 1625156677
transform -1 0 1748 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_476
timestamp 1625156677
transform -1 0 1772 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_339
timestamp 1625156677
transform -1 0 1788 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_513
timestamp 1625156677
transform 1 0 1788 0 1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_263
timestamp 1625156677
transform -1 0 1868 0 1 3105
box -2 -3 58 103
use BUFX2  BUFX2_219
timestamp 1625156677
transform 1 0 1868 0 1 3105
box -2 -3 26 103
use FILL  FILL_31_3_0
timestamp 1625156677
transform 1 0 1892 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_3_1
timestamp 1625156677
transform 1 0 1900 0 1 3105
box -2 -3 10 103
use XOR2X1  XOR2X1_259
timestamp 1625156677
transform 1 0 1908 0 1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_258
timestamp 1625156677
transform 1 0 1964 0 1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_262
timestamp 1625156677
transform -1 0 2076 0 1 3105
box -2 -3 58 103
use NOR2X1  NOR2X1_330
timestamp 1625156677
transform 1 0 2076 0 1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_264
timestamp 1625156677
transform -1 0 2156 0 1 3105
box -2 -3 58 103
use NOR2X1  NOR2X1_321
timestamp 1625156677
transform -1 0 2180 0 1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_194
timestamp 1625156677
transform 1 0 2180 0 1 3105
box -2 -3 58 103
use BUFX2  BUFX2_220
timestamp 1625156677
transform -1 0 2260 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_429
timestamp 1625156677
transform 1 0 2260 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_565
timestamp 1625156677
transform 1 0 2276 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_566
timestamp 1625156677
transform -1 0 2324 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_523
timestamp 1625156677
transform -1 0 2356 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_331
timestamp 1625156677
transform -1 0 2380 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_532
timestamp 1625156677
transform 1 0 2380 0 1 3105
box -2 -3 26 103
use FILL  FILL_31_4_0
timestamp 1625156677
transform -1 0 2412 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_4_1
timestamp 1625156677
transform -1 0 2420 0 1 3105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_198
timestamp 1625156677
transform -1 0 2476 0 1 3105
box -2 -3 58 103
use NOR2X1  NOR2X1_333
timestamp 1625156677
transform 1 0 2476 0 1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_268
timestamp 1625156677
transform 1 0 2500 0 1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_244
timestamp 1625156677
transform 1 0 2556 0 1 3105
box -2 -3 58 103
use OAI21X1  OAI21X1_471
timestamp 1625156677
transform 1 0 2612 0 1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_423
timestamp 1625156677
transform 1 0 2644 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_299
timestamp 1625156677
transform -1 0 2700 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_516
timestamp 1625156677
transform -1 0 2724 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_378
timestamp 1625156677
transform 1 0 2724 0 1 3105
box -2 -3 18 103
use AND2X2  AND2X2_139
timestamp 1625156677
transform 1 0 2740 0 1 3105
box -2 -3 34 103
use AND2X2  AND2X2_140
timestamp 1625156677
transform 1 0 2772 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_414
timestamp 1625156677
transform 1 0 2804 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_551
timestamp 1625156677
transform 1 0 2820 0 1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_277
timestamp 1625156677
transform 1 0 2844 0 1 3105
box -2 -3 58 103
use FILL  FILL_31_5_0
timestamp 1625156677
transform -1 0 2908 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_5_1
timestamp 1625156677
transform -1 0 2916 0 1 3105
box -2 -3 10 103
use XOR2X1  XOR2X1_276
timestamp 1625156677
transform -1 0 2972 0 1 3105
box -2 -3 58 103
use INVX1  INVX1_396
timestamp 1625156677
transform -1 0 2988 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_489
timestamp 1625156677
transform 1 0 2988 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_534
timestamp 1625156677
transform 1 0 3020 0 1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_275
timestamp 1625156677
transform -1 0 3100 0 1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_254
timestamp 1625156677
transform 1 0 3100 0 1 3105
box -2 -3 58 103
use OAI21X1  OAI21X1_492
timestamp 1625156677
transform -1 0 3188 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_544
timestamp 1625156677
transform 1 0 3188 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_312
timestamp 1625156677
transform 1 0 3212 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_536
timestamp 1625156677
transform -1 0 3260 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_398
timestamp 1625156677
transform 1 0 3260 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_503
timestamp 1625156677
transform -1 0 3308 0 1 3105
box -2 -3 34 103
use AND2X2  AND2X2_154
timestamp 1625156677
transform -1 0 3340 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_590
timestamp 1625156677
transform -1 0 3364 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_453
timestamp 1625156677
transform 1 0 3364 0 1 3105
box -2 -3 18 103
use BUFX2  BUFX2_234
timestamp 1625156677
transform 1 0 3380 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_588
timestamp 1625156677
transform 1 0 3404 0 1 3105
box -2 -3 18 103
use FILL  FILL_31_6_0
timestamp 1625156677
transform 1 0 3420 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_6_1
timestamp 1625156677
transform 1 0 3428 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_632
timestamp 1625156677
transform 1 0 3436 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_587
timestamp 1625156677
transform 1 0 3468 0 1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_531
timestamp 1625156677
transform 1 0 3484 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_699
timestamp 1625156677
transform 1 0 3516 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_700
timestamp 1625156677
transform -1 0 3564 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_586
timestamp 1625156677
transform -1 0 3580 0 1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_443
timestamp 1625156677
transform -1 0 3604 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_698
timestamp 1625156677
transform -1 0 3628 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_697
timestamp 1625156677
transform -1 0 3652 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_585
timestamp 1625156677
transform 1 0 3652 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1625156677
transform 1 0 3668 0 1 3105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_13
timestamp 1625156677
transform -1 0 3836 0 1 3105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1625156677
transform 1 0 3836 0 1 3105
box -2 -3 98 103
use FILL  FILL_31_7_0
timestamp 1625156677
transform -1 0 3940 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_7_1
timestamp 1625156677
transform -1 0 3948 0 1 3105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_35
timestamp 1625156677
transform -1 0 4020 0 1 3105
box -2 -3 74 103
use XNOR2X1  XNOR2X1_247
timestamp 1625156677
transform -1 0 4076 0 1 3105
box -2 -3 58 103
use BUFX2  BUFX2_43
timestamp 1625156677
transform 1 0 4076 0 1 3105
box -2 -3 26 103
use BUFX2  BUFX2_57
timestamp 1625156677
transform 1 0 4100 0 1 3105
box -2 -3 26 103
use AND2X2  AND2X2_191
timestamp 1625156677
transform 1 0 4124 0 1 3105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_28
timestamp 1625156677
transform 1 0 4156 0 1 3105
box -2 -3 74 103
use INVX2  INVX2_91
timestamp 1625156677
transform -1 0 4244 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_696
timestamp 1625156677
transform 1 0 4244 0 1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_246
timestamp 1625156677
transform -1 0 4324 0 1 3105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1625156677
transform 1 0 4324 0 1 3105
box -2 -3 98 103
use FILL  FILL_31_8_0
timestamp 1625156677
transform -1 0 4428 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_8_1
timestamp 1625156677
transform -1 0 4436 0 1 3105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_245
timestamp 1625156677
transform -1 0 4492 0 1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_288
timestamp 1625156677
transform -1 0 4548 0 1 3105
box -2 -3 58 103
use CLKBUF1  CLKBUF1_42
timestamp 1625156677
transform 1 0 4548 0 1 3105
box -2 -3 74 103
use INVX1  INVX1_584
timestamp 1625156677
transform 1 0 4620 0 1 3105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1625156677
transform 1 0 4636 0 1 3105
box -2 -3 98 103
use BUFX4  BUFX4_23
timestamp 1625156677
transform 1 0 4732 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1625156677
transform 1 0 4764 0 1 3105
box -2 -3 98 103
use MUX2X1  MUX2X1_20
timestamp 1625156677
transform 1 0 4860 0 1 3105
box -2 -3 50 103
use NOR3X1  NOR3X1_20
timestamp 1625156677
transform -1 0 4972 0 1 3105
box -2 -3 66 103
use FILL  FILL_31_9_0
timestamp 1625156677
transform 1 0 4972 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_9_1
timestamp 1625156677
transform 1 0 4980 0 1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1625156677
transform 1 0 4988 0 1 3105
box -2 -3 98 103
use MUX2X1  MUX2X1_17
timestamp 1625156677
transform 1 0 5084 0 1 3105
box -2 -3 50 103
use NOR3X1  NOR3X1_17
timestamp 1625156677
transform 1 0 5132 0 1 3105
box -2 -3 66 103
use BUFX2  BUFX2_20
timestamp 1625156677
transform 1 0 5196 0 1 3105
box -2 -3 26 103
use BUFX2  BUFX2_99
timestamp 1625156677
transform -1 0 5244 0 1 3105
box -2 -3 26 103
use BUFX2  BUFX2_17
timestamp 1625156677
transform -1 0 5268 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_185
timestamp 1625156677
transform 1 0 5268 0 1 3105
box -2 -3 34 103
use FILL  FILL_32_1
timestamp 1625156677
transform 1 0 5300 0 1 3105
box -2 -3 10 103
use FILL  FILL_32_2
timestamp 1625156677
transform 1 0 5308 0 1 3105
box -2 -3 10 103
use BUFX2  BUFX2_105
timestamp 1625156677
transform -1 0 28 0 -1 3105
box -2 -3 26 103
use BUFX2  BUFX2_121
timestamp 1625156677
transform 1 0 28 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_252
timestamp 1625156677
transform -1 0 84 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_381
timestamp 1625156677
transform 1 0 84 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_455
timestamp 1625156677
transform 1 0 116 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_257
timestamp 1625156677
transform -1 0 172 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_448
timestamp 1625156677
transform 1 0 172 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_312
timestamp 1625156677
transform 1 0 196 0 -1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_379
timestamp 1625156677
transform -1 0 244 0 -1 3105
box -2 -3 34 103
use AOI22X1  AOI22X1_14
timestamp 1625156677
transform -1 0 284 0 -1 3105
box -2 -3 42 103
use INVX1  INVX1_314
timestamp 1625156677
transform 1 0 284 0 -1 3105
box -2 -3 18 103
use XOR2X1  XOR2X1_208
timestamp 1625156677
transform -1 0 356 0 -1 3105
box -2 -3 58 103
use FILL  FILL_30_0_0
timestamp 1625156677
transform -1 0 364 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_0_1
timestamp 1625156677
transform -1 0 372 0 -1 3105
box -2 -3 10 103
use BUFX2  BUFX2_204
timestamp 1625156677
transform -1 0 396 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_453
timestamp 1625156677
transform 1 0 396 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_260
timestamp 1625156677
transform 1 0 420 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_412
timestamp 1625156677
transform 1 0 444 0 -1 3105
box -2 -3 34 103
use AND2X2  AND2X2_122
timestamp 1625156677
transform -1 0 508 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_250
timestamp 1625156677
transform 1 0 508 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_438
timestamp 1625156677
transform -1 0 556 0 -1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_221
timestamp 1625156677
transform -1 0 612 0 -1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_230
timestamp 1625156677
transform 1 0 612 0 -1 3105
box -2 -3 58 103
use NAND2X1  NAND2X1_471
timestamp 1625156677
transform -1 0 692 0 -1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_179
timestamp 1625156677
transform 1 0 692 0 -1 3105
box -2 -3 58 103
use NOR2X1  NOR2X1_282
timestamp 1625156677
transform -1 0 772 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_444
timestamp 1625156677
transform 1 0 772 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_445
timestamp 1625156677
transform 1 0 804 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_349
timestamp 1625156677
transform -1 0 852 0 -1 3105
box -2 -3 18 103
use FILL  FILL_30_1_0
timestamp 1625156677
transform 1 0 852 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_1_1
timestamp 1625156677
transform 1 0 860 0 -1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_485
timestamp 1625156677
transform 1 0 868 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_484
timestamp 1625156677
transform -1 0 916 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_440
timestamp 1625156677
transform 1 0 916 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_347
timestamp 1625156677
transform 1 0 948 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_441
timestamp 1625156677
transform 1 0 964 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_401
timestamp 1625156677
transform -1 0 1028 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_346
timestamp 1625156677
transform -1 0 1044 0 -1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_402
timestamp 1625156677
transform -1 0 1076 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_407
timestamp 1625156677
transform -1 0 1108 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_268
timestamp 1625156677
transform 1 0 1108 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_438
timestamp 1625156677
transform 1 0 1140 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_276
timestamp 1625156677
transform 1 0 1172 0 -1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_399
timestamp 1625156677
transform -1 0 1228 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_435
timestamp 1625156677
transform 1 0 1228 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_446
timestamp 1625156677
transform 1 0 1260 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_341
timestamp 1625156677
transform -1 0 1308 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_487
timestamp 1625156677
transform 1 0 1308 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_270
timestamp 1625156677
transform 1 0 1332 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_2_0
timestamp 1625156677
transform 1 0 1364 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_2_1
timestamp 1625156677
transform 1 0 1372 0 -1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_479
timestamp 1625156677
transform 1 0 1380 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_433
timestamp 1625156677
transform 1 0 1404 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_275
timestamp 1625156677
transform -1 0 1460 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_478
timestamp 1625156677
transform 1 0 1460 0 -1 3105
box -2 -3 26 103
use AND2X2  AND2X2_131
timestamp 1625156677
transform 1 0 1484 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_397
timestamp 1625156677
transform -1 0 1548 0 -1 3105
box -2 -3 34 103
use XOR2X1  XOR2X1_225
timestamp 1625156677
transform 1 0 1548 0 -1 3105
box -2 -3 58 103
use OAI21X1  OAI21X1_432
timestamp 1625156677
transform 1 0 1604 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_477
timestamp 1625156677
transform 1 0 1636 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_324
timestamp 1625156677
transform -1 0 1756 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_306
timestamp 1625156677
transform -1 0 1852 0 -1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_327
timestamp 1625156677
transform 1 0 1852 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_3_0
timestamp 1625156677
transform 1 0 1876 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_3_1
timestamp 1625156677
transform 1 0 1884 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_353
timestamp 1625156677
transform 1 0 1892 0 -1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_560
timestamp 1625156677
transform 1 0 1988 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_426
timestamp 1625156677
transform -1 0 2028 0 -1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_456
timestamp 1625156677
transform -1 0 2060 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_521
timestamp 1625156677
transform -1 0 2092 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_520
timestamp 1625156677
transform 1 0 2092 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_425
timestamp 1625156677
transform 1 0 2124 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_561
timestamp 1625156677
transform 1 0 2140 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_428
timestamp 1625156677
transform 1 0 2164 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_567
timestamp 1625156677
transform 1 0 2180 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_568
timestamp 1625156677
transform 1 0 2204 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_332
timestamp 1625156677
transform 1 0 2228 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_430
timestamp 1625156677
transform 1 0 2252 0 -1 3105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_199
timestamp 1625156677
transform 1 0 2268 0 -1 3105
box -2 -3 58 103
use OAI21X1  OAI21X1_504
timestamp 1625156677
transform 1 0 2324 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_319
timestamp 1625156677
transform -1 0 2380 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_410
timestamp 1625156677
transform 1 0 2380 0 -1 3105
box -2 -3 18 103
use FILL  FILL_30_4_0
timestamp 1625156677
transform 1 0 2396 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_4_1
timestamp 1625156677
transform 1 0 2404 0 -1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_546
timestamp 1625156677
transform 1 0 2412 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_547
timestamp 1625156677
transform -1 0 2460 0 -1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_195
timestamp 1625156677
transform -1 0 2516 0 -1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_243
timestamp 1625156677
transform 1 0 2516 0 -1 3105
box -2 -3 58 103
use NOR2X1  NOR2X1_298
timestamp 1625156677
transform -1 0 2596 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_470
timestamp 1625156677
transform 1 0 2596 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_515
timestamp 1625156677
transform 1 0 2628 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_514
timestamp 1625156677
transform -1 0 2676 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_377
timestamp 1625156677
transform 1 0 2676 0 -1 3105
box -2 -3 18 103
use AND2X2  AND2X2_138
timestamp 1625156677
transform 1 0 2692 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_608
timestamp 1625156677
transform 1 0 2724 0 -1 3105
box -2 -3 26 103
use BUFX2  BUFX2_228
timestamp 1625156677
transform 1 0 2748 0 -1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_202
timestamp 1625156677
transform -1 0 2828 0 -1 3105
box -2 -3 58 103
use NOR2X1  NOR2X1_345
timestamp 1625156677
transform 1 0 2828 0 -1 3105
box -2 -3 26 103
use AND2X2  AND2X2_157
timestamp 1625156677
transform 1 0 2852 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_5_0
timestamp 1625156677
transform 1 0 2884 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_5_1
timestamp 1625156677
transform 1 0 2892 0 -1 3105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_203
timestamp 1625156677
transform 1 0 2900 0 -1 3105
box -2 -3 58 103
use OAI21X1  OAI21X1_542
timestamp 1625156677
transform 1 0 2956 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_343
timestamp 1625156677
transform -1 0 3012 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_585
timestamp 1625156677
transform 1 0 3012 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_584
timestamp 1625156677
transform -1 0 3060 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_448
timestamp 1625156677
transform 1 0 3060 0 -1 3105
box -2 -3 18 103
use XOR2X1  XOR2X1_274
timestamp 1625156677
transform -1 0 3132 0 -1 3105
box -2 -3 58 103
use BUFX2  BUFX2_235
timestamp 1625156677
transform 1 0 3132 0 -1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_279
timestamp 1625156677
transform -1 0 3212 0 -1 3105
box -2 -3 58 103
use OAI21X1  OAI21X1_546
timestamp 1625156677
transform 1 0 3212 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_591
timestamp 1625156677
transform 1 0 3244 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_346
timestamp 1625156677
transform -1 0 3292 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_342
timestamp 1625156677
transform 1 0 3292 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_535
timestamp 1625156677
transform 1 0 3316 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_442
timestamp 1625156677
transform 1 0 3348 0 -1 3105
box -2 -3 18 103
use INVX1  INVX1_441
timestamp 1625156677
transform 1 0 3364 0 -1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_467
timestamp 1625156677
transform -1 0 3412 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_6_0
timestamp 1625156677
transform 1 0 3412 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_6_1
timestamp 1625156677
transform 1 0 3420 0 -1 3105
box -2 -3 10 103
use NAND3X1  NAND3X1_466
timestamp 1625156677
transform 1 0 3428 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_443
timestamp 1625156677
transform 1 0 3460 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_536
timestamp 1625156677
transform -1 0 3508 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_307
timestamp 1625156677
transform 1 0 3508 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_468
timestamp 1625156677
transform -1 0 3572 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_440
timestamp 1625156677
transform -1 0 3588 0 -1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_472
timestamp 1625156677
transform -1 0 3620 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_308
timestamp 1625156677
transform 1 0 3620 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_340
timestamp 1625156677
transform 1 0 3652 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_538
timestamp 1625156677
transform -1 0 3708 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_583
timestamp 1625156677
transform -1 0 3732 0 -1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_287
timestamp 1625156677
transform -1 0 3788 0 -1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_293
timestamp 1625156677
transform -1 0 3844 0 -1 3105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_201
timestamp 1625156677
transform -1 0 3900 0 -1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_292
timestamp 1625156677
transform -1 0 3956 0 -1 3105
box -2 -3 58 103
use FILL  FILL_30_7_0
timestamp 1625156677
transform 1 0 3956 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_7_1
timestamp 1625156677
transform 1 0 3964 0 -1 3105
box -2 -3 10 103
use BUFX4  BUFX4_2
timestamp 1625156677
transform 1 0 3972 0 -1 3105
box -2 -3 34 103
use AND2X2  AND2X2_192
timestamp 1625156677
transform 1 0 4004 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_582
timestamp 1625156677
transform 1 0 4036 0 -1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_529
timestamp 1625156677
transform 1 0 4052 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_530
timestamp 1625156677
transform 1 0 4084 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_631
timestamp 1625156677
transform -1 0 4148 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_441
timestamp 1625156677
transform -1 0 4172 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_581
timestamp 1625156677
transform -1 0 4188 0 -1 3105
box -2 -3 18 103
use XOR2X1  XOR2X1_290
timestamp 1625156677
transform 1 0 4188 0 -1 3105
box -2 -3 58 103
use XOR2X1  XOR2X1_306
timestamp 1625156677
transform -1 0 4300 0 -1 3105
box -2 -3 58 103
use NAND3X1  NAND3X1_528
timestamp 1625156677
transform -1 0 4332 0 -1 3105
box -2 -3 34 103
use AND2X2  AND2X2_189
timestamp 1625156677
transform 1 0 4332 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_437
timestamp 1625156677
transform 1 0 4364 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_438
timestamp 1625156677
transform 1 0 4388 0 -1 3105
box -2 -3 26 103
use AND2X2  AND2X2_188
timestamp 1625156677
transform -1 0 4444 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_8_0
timestamp 1625156677
transform -1 0 4452 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_8_1
timestamp 1625156677
transform -1 0 4460 0 -1 3105
box -2 -3 10 103
use AND2X2  AND2X2_190
timestamp 1625156677
transform -1 0 4492 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_439
timestamp 1625156677
transform -1 0 4516 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_440
timestamp 1625156677
transform 1 0 4516 0 -1 3105
box -2 -3 26 103
use XOR2X1  XOR2X1_305
timestamp 1625156677
transform -1 0 4596 0 -1 3105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1625156677
transform 1 0 4596 0 -1 3105
box -2 -3 98 103
use INVX1  INVX1_580
timestamp 1625156677
transform 1 0 4692 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_630
timestamp 1625156677
transform 1 0 4708 0 -1 3105
box -2 -3 34 103
use INVX2  INVX2_90
timestamp 1625156677
transform 1 0 4740 0 -1 3105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_244
timestamp 1625156677
transform -1 0 4812 0 -1 3105
box -2 -3 58 103
use NAND2X1  NAND2X1_695
timestamp 1625156677
transform -1 0 4836 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_579
timestamp 1625156677
transform -1 0 4852 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_694
timestamp 1625156677
transform 1 0 4852 0 -1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_243
timestamp 1625156677
transform 1 0 4876 0 -1 3105
box -2 -3 58 103
use FILL  FILL_30_9_0
timestamp 1625156677
transform 1 0 4932 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_9_1
timestamp 1625156677
transform 1 0 4940 0 -1 3105
box -2 -3 10 103
use MUX2X1  MUX2X1_18
timestamp 1625156677
transform 1 0 4948 0 -1 3105
box -2 -3 50 103
use NOR3X1  NOR3X1_18
timestamp 1625156677
transform -1 0 5060 0 -1 3105
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1625156677
transform 1 0 5060 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1625156677
transform 1 0 5156 0 -1 3105
box -2 -3 98 103
use BUFX2  BUFX2_18
timestamp 1625156677
transform 1 0 5252 0 -1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_188
timestamp 1625156677
transform 1 0 5276 0 -1 3105
box -2 -3 34 103
use FILL  FILL_31_1
timestamp 1625156677
transform -1 0 5316 0 -1 3105
box -2 -3 10 103
use BUFX2  BUFX2_30
timestamp 1625156677
transform 1 0 4 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_375
timestamp 1625156677
transform -1 0 60 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_308
timestamp 1625156677
transform -1 0 76 0 1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_376
timestamp 1625156677
transform -1 0 108 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_309
timestamp 1625156677
transform -1 0 124 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_403
timestamp 1625156677
transform -1 0 156 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_310
timestamp 1625156677
transform -1 0 172 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_402
timestamp 1625156677
transform -1 0 204 0 1 2905
box -2 -3 34 103
use BUFX2  BUFX2_205
timestamp 1625156677
transform 1 0 204 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_378
timestamp 1625156677
transform 1 0 228 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_446
timestamp 1625156677
transform -1 0 284 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_447
timestamp 1625156677
transform -1 0 308 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_311
timestamp 1625156677
transform 1 0 308 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_406
timestamp 1625156677
transform -1 0 356 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_0_0
timestamp 1625156677
transform 1 0 356 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_0_1
timestamp 1625156677
transform 1 0 364 0 1 2905
box -2 -3 10 103
use NOR2X1  NOR2X1_258
timestamp 1625156677
transform 1 0 372 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_407
timestamp 1625156677
transform 1 0 396 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_452
timestamp 1625156677
transform 1 0 428 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_451
timestamp 1625156677
transform -1 0 476 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_315
timestamp 1625156677
transform -1 0 492 0 1 2905
box -2 -3 18 103
use XNOR2X1  XNOR2X1_175
timestamp 1625156677
transform -1 0 548 0 1 2905
box -2 -3 58 103
use INVX1  INVX1_301
timestamp 1625156677
transform -1 0 564 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_394
timestamp 1625156677
transform 1 0 564 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_299
timestamp 1625156677
transform -1 0 692 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_470
timestamp 1625156677
transform -1 0 716 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_271
timestamp 1625156677
transform 1 0 716 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_334
timestamp 1625156677
transform -1 0 756 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_428
timestamp 1625156677
transform 1 0 756 0 1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_321
timestamp 1625156677
transform -1 0 884 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_1_0
timestamp 1625156677
transform -1 0 892 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_1_1
timestamp 1625156677
transform -1 0 900 0 1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_301
timestamp 1625156677
transform -1 0 996 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_348
timestamp 1625156677
transform 1 0 996 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_310
timestamp 1625156677
transform -1 0 1108 0 1 2905
box -2 -3 98 103
use OAI21X1  OAI21X1_439
timestamp 1625156677
transform 1 0 1108 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_279
timestamp 1625156677
transform -1 0 1164 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_343
timestamp 1625156677
transform 1 0 1164 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_482
timestamp 1625156677
transform 1 0 1180 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_481
timestamp 1625156677
transform -1 0 1228 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_308
timestamp 1625156677
transform -1 0 1324 0 1 2905
box -2 -3 98 103
use FILL  FILL_29_2_0
timestamp 1625156677
transform -1 0 1332 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_2_1
timestamp 1625156677
transform -1 0 1340 0 1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_317
timestamp 1625156677
transform -1 0 1436 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_550
timestamp 1625156677
transform -1 0 1452 0 1 2905
box -2 -3 18 103
use INVX1  INVX1_340
timestamp 1625156677
transform 1 0 1452 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_325
timestamp 1625156677
transform -1 0 1564 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_563
timestamp 1625156677
transform -1 0 1580 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_327
timestamp 1625156677
transform -1 0 1676 0 1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_349
timestamp 1625156677
transform 1 0 1676 0 1 2905
box -2 -3 98 103
use INVX1  INVX1_419
timestamp 1625156677
transform 1 0 1772 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_558
timestamp 1625156677
transform 1 0 1788 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_514
timestamp 1625156677
transform -1 0 1844 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_557
timestamp 1625156677
transform -1 0 1868 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_3_0
timestamp 1625156677
transform -1 0 1876 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_3_1
timestamp 1625156677
transform -1 0 1884 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_515
timestamp 1625156677
transform -1 0 1916 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_525
timestamp 1625156677
transform 1 0 1916 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_562
timestamp 1625156677
transform -1 0 1972 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_305
timestamp 1625156677
transform 1 0 1972 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_457
timestamp 1625156677
transform -1 0 2036 0 1 2905
box -2 -3 34 103
use AOI22X1  AOI22X1_20
timestamp 1625156677
transform -1 0 2076 0 1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_524
timestamp 1625156677
transform 1 0 2076 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_432
timestamp 1625156677
transform 1 0 2108 0 1 2905
box -2 -3 18 103
use INVX1  INVX1_431
timestamp 1625156677
transform -1 0 2140 0 1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_460
timestamp 1625156677
transform -1 0 2172 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_306
timestamp 1625156677
transform 1 0 2172 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_526
timestamp 1625156677
transform 1 0 2204 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_433
timestamp 1625156677
transform 1 0 2236 0 1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_461
timestamp 1625156677
transform 1 0 2252 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_570
timestamp 1625156677
transform 1 0 2284 0 1 2905
box -2 -3 26 103
use AND2X2  AND2X2_149
timestamp 1625156677
transform 1 0 2308 0 1 2905
box -2 -3 34 103
use XOR2X1  XOR2X1_285
timestamp 1625156677
transform 1 0 2340 0 1 2905
box -2 -3 58 103
use FILL  FILL_29_4_0
timestamp 1625156677
transform -1 0 2404 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_4_1
timestamp 1625156677
transform -1 0 2412 0 1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_322
timestamp 1625156677
transform -1 0 2508 0 1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_604
timestamp 1625156677
transform -1 0 2532 0 1 2905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_207
timestamp 1625156677
transform -1 0 2588 0 1 2905
box -2 -3 58 103
use NAND2X1  NAND2X1_605
timestamp 1625156677
transform -1 0 2612 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_356
timestamp 1625156677
transform -1 0 2636 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_466
timestamp 1625156677
transform -1 0 2652 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_606
timestamp 1625156677
transform 1 0 2652 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_468
timestamp 1625156677
transform -1 0 2692 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_564
timestamp 1625156677
transform -1 0 2724 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_471
timestamp 1625156677
transform 1 0 2724 0 1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_487
timestamp 1625156677
transform 1 0 2740 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_322
timestamp 1625156677
transform -1 0 2804 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_469
timestamp 1625156677
transform 1 0 2804 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_562
timestamp 1625156677
transform -1 0 2852 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_470
timestamp 1625156677
transform 1 0 2852 0 1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_486
timestamp 1625156677
transform 1 0 2868 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_5_0
timestamp 1625156677
transform -1 0 2908 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_5_1
timestamp 1625156677
transform -1 0 2916 0 1 2905
box -2 -3 10 103
use BUFX2  BUFX2_233
timestamp 1625156677
transform -1 0 2940 0 1 2905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_205
timestamp 1625156677
transform 1 0 2940 0 1 2905
box -2 -3 58 103
use NOR3X1  NOR3X1_86
timestamp 1625156677
transform -1 0 3060 0 1 2905
box -2 -3 66 103
use OAI21X1  OAI21X1_548
timestamp 1625156677
transform 1 0 3060 0 1 2905
box -2 -3 34 103
use AND2X2  AND2X2_156
timestamp 1625156677
transform 1 0 3092 0 1 2905
box -2 -3 34 103
use INVX2  INVX2_73
timestamp 1625156677
transform -1 0 3140 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_551
timestamp 1625156677
transform 1 0 3140 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_349
timestamp 1625156677
transform 1 0 3172 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_350
timestamp 1625156677
transform -1 0 3220 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_475
timestamp 1625156677
transform 1 0 3220 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_539
timestamp 1625156677
transform 1 0 3252 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_580
timestamp 1625156677
transform 1 0 3284 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_444
timestamp 1625156677
transform -1 0 3324 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_579
timestamp 1625156677
transform -1 0 3348 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_469
timestamp 1625156677
transform -1 0 3380 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_540
timestamp 1625156677
transform 1 0 3380 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_6_0
timestamp 1625156677
transform -1 0 3420 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_6_1
timestamp 1625156677
transform -1 0 3428 0 1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_586
timestamp 1625156677
transform -1 0 3452 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_344
timestamp 1625156677
transform -1 0 3476 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_447
timestamp 1625156677
transform -1 0 3492 0 1 2905
box -2 -3 18 103
use INVX1  INVX1_445
timestamp 1625156677
transform 1 0 3492 0 1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_470
timestamp 1625156677
transform -1 0 3540 0 1 2905
box -2 -3 34 103
use AOI22X1  AOI22X1_21
timestamp 1625156677
transform 1 0 3540 0 1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_545
timestamp 1625156677
transform -1 0 3612 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_588
timestamp 1625156677
transform 1 0 3612 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_451
timestamp 1625156677
transform 1 0 3636 0 1 2905
box -2 -3 18 103
use AOI21X1  AOI21X1_314
timestamp 1625156677
transform -1 0 3684 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_473
timestamp 1625156677
transform 1 0 3684 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_581
timestamp 1625156677
transform 1 0 3716 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_313
timestamp 1625156677
transform 1 0 3740 0 1 2905
box -2 -3 34 103
use BUFX2  BUFX2_34
timestamp 1625156677
transform 1 0 3772 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_544
timestamp 1625156677
transform -1 0 3828 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_341
timestamp 1625156677
transform -1 0 3852 0 1 2905
box -2 -3 26 103
use XOR2X1  XOR2X1_308
timestamp 1625156677
transform -1 0 3908 0 1 2905
box -2 -3 58 103
use FILL  FILL_29_7_0
timestamp 1625156677
transform -1 0 3916 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_7_1
timestamp 1625156677
transform -1 0 3924 0 1 2905
box -2 -3 10 103
use NOR3X1  NOR3X1_83
timestamp 1625156677
transform -1 0 3988 0 1 2905
box -2 -3 66 103
use XNOR2X1  XNOR2X1_200
timestamp 1625156677
transform -1 0 4044 0 1 2905
box -2 -3 58 103
use INVX1  INVX1_583
timestamp 1625156677
transform 1 0 4044 0 1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_442
timestamp 1625156677
transform 1 0 4060 0 1 2905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_248
timestamp 1625156677
transform -1 0 4140 0 1 2905
box -2 -3 58 103
use NOR2X1  NOR2X1_338
timestamp 1625156677
transform 1 0 4140 0 1 2905
box -2 -3 26 103
use XOR2X1  XOR2X1_291
timestamp 1625156677
transform -1 0 4220 0 1 2905
box -2 -3 58 103
use BUFX2  BUFX2_246
timestamp 1625156677
transform 1 0 4220 0 1 2905
box -2 -3 26 103
use XOR2X1  XOR2X1_307
timestamp 1625156677
transform -1 0 4300 0 1 2905
box -2 -3 58 103
use BUFX2  BUFX2_245
timestamp 1625156677
transform 1 0 4300 0 1 2905
box -2 -3 26 103
use BUFX2  BUFX2_244
timestamp 1625156677
transform 1 0 4324 0 1 2905
box -2 -3 26 103
use XOR2X1  XOR2X1_289
timestamp 1625156677
transform 1 0 4348 0 1 2905
box -2 -3 58 103
use AND2X2  AND2X2_57
timestamp 1625156677
transform 1 0 4404 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_8_0
timestamp 1625156677
transform 1 0 4436 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_8_1
timestamp 1625156677
transform 1 0 4444 0 1 2905
box -2 -3 10 103
use NOR2X1  NOR2X1_109
timestamp 1625156677
transform 1 0 4452 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_194
timestamp 1625156677
transform 1 0 4476 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_111
timestamp 1625156677
transform 1 0 4500 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_163
timestamp 1625156677
transform 1 0 4516 0 1 2905
box -2 -3 34 103
use NOR3X1  NOR3X1_44
timestamp 1625156677
transform 1 0 4548 0 1 2905
box -2 -3 66 103
use BUFX2  BUFX2_64
timestamp 1625156677
transform 1 0 4612 0 1 2905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_41
timestamp 1625156677
transform 1 0 4636 0 1 2905
box -2 -3 74 103
use NOR2X1  NOR2X1_435
timestamp 1625156677
transform -1 0 4732 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_436
timestamp 1625156677
transform 1 0 4732 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1625156677
transform 1 0 4756 0 1 2905
box -2 -3 98 103
use AND2X2  AND2X2_58
timestamp 1625156677
transform -1 0 4884 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_197
timestamp 1625156677
transform 1 0 4884 0 1 2905
box -2 -3 26 103
use NOR3X1  NOR3X1_10
timestamp 1625156677
transform -1 0 4972 0 1 2905
box -2 -3 66 103
use FILL  FILL_29_9_0
timestamp 1625156677
transform 1 0 4972 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_9_1
timestamp 1625156677
transform 1 0 4980 0 1 2905
box -2 -3 10 103
use MUX2X1  MUX2X1_10
timestamp 1625156677
transform 1 0 4988 0 1 2905
box -2 -3 50 103
use BUFX2  BUFX2_10
timestamp 1625156677
transform 1 0 5036 0 1 2905
box -2 -3 26 103
use MUX2X1  MUX2X1_9
timestamp 1625156677
transform 1 0 5060 0 1 2905
box -2 -3 50 103
use NOR3X1  NOR3X1_9
timestamp 1625156677
transform 1 0 5108 0 1 2905
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1625156677
transform 1 0 5172 0 1 2905
box -2 -3 98 103
use AOI21X1  AOI21X1_132
timestamp 1625156677
transform -1 0 5300 0 1 2905
box -2 -3 34 103
use FILL  FILL_30_1
timestamp 1625156677
transform 1 0 5300 0 1 2905
box -2 -3 10 103
use FILL  FILL_30_2
timestamp 1625156677
transform 1 0 5308 0 1 2905
box -2 -3 10 103
use XOR2X1  XOR2X1_210
timestamp 1625156677
transform -1 0 60 0 -1 2905
box -2 -3 58 103
use BUFX2  BUFX2_203
timestamp 1625156677
transform -1 0 84 0 -1 2905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_164
timestamp 1625156677
transform 1 0 84 0 -1 2905
box -2 -3 58 103
use NOR2X1  NOR2X1_230
timestamp 1625156677
transform 1 0 140 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_360
timestamp 1625156677
transform -1 0 196 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_302
timestamp 1625156677
transform -1 0 292 0 -1 2905
box -2 -3 98 103
use XOR2X1  XOR2X1_220
timestamp 1625156677
transform -1 0 348 0 -1 2905
box -2 -3 58 103
use FILL  FILL_28_0_0
timestamp 1625156677
transform 1 0 348 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_0_1
timestamp 1625156677
transform 1 0 356 0 -1 2905
box -2 -3 10 103
use AND2X2  AND2X2_116
timestamp 1625156677
transform 1 0 364 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_259
timestamp 1625156677
transform 1 0 396 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_409
timestamp 1625156677
transform 1 0 420 0 -1 2905
box -2 -3 34 103
use XOR2X1  XOR2X1_207
timestamp 1625156677
transform 1 0 452 0 -1 2905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_311
timestamp 1625156677
transform -1 0 604 0 -1 2905
box -2 -3 98 103
use XOR2X1  XOR2X1_223
timestamp 1625156677
transform -1 0 660 0 -1 2905
box -2 -3 58 103
use NOR2X1  NOR2X1_273
timestamp 1625156677
transform -1 0 684 0 -1 2905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_178
timestamp 1625156677
transform 1 0 684 0 -1 2905
box -2 -3 58 103
use XOR2X1  XOR2X1_222
timestamp 1625156677
transform -1 0 796 0 -1 2905
box -2 -3 58 103
use NAND2X1  NAND2X1_437
timestamp 1625156677
transform -1 0 820 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_1_0
timestamp 1625156677
transform -1 0 828 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_1_1
timestamp 1625156677
transform -1 0 836 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_309
timestamp 1625156677
transform -1 0 932 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_319
timestamp 1625156677
transform -1 0 1028 0 -1 2905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_34
timestamp 1625156677
transform -1 0 1100 0 -1 2905
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_318
timestamp 1625156677
transform -1 0 1196 0 -1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_420
timestamp 1625156677
transform -1 0 1220 0 -1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_316
timestamp 1625156677
transform -1 0 1316 0 -1 2905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_46
timestamp 1625156677
transform 1 0 1316 0 -1 2905
box -2 -3 74 103
use FILL  FILL_28_2_0
timestamp 1625156677
transform -1 0 1396 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_2_1
timestamp 1625156677
transform -1 0 1404 0 -1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_329
timestamp 1625156677
transform -1 0 1500 0 -1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_675
timestamp 1625156677
transform -1 0 1524 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_324
timestamp 1625156677
transform 1 0 1524 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_511
timestamp 1625156677
transform 1 0 1548 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_420
timestamp 1625156677
transform 1 0 1580 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_522
timestamp 1625156677
transform 1 0 1596 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_452
timestamp 1625156677
transform -1 0 1660 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_301
timestamp 1625156677
transform -1 0 1692 0 -1 2905
box -2 -3 34 103
use NOR3X1  NOR3X1_81
timestamp 1625156677
transform -1 0 1756 0 -1 2905
box -2 -3 66 103
use OAI21X1  OAI21X1_518
timestamp 1625156677
transform 1 0 1756 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_329
timestamp 1625156677
transform 1 0 1788 0 -1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_451
timestamp 1625156677
transform 1 0 1812 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_304
timestamp 1625156677
transform 1 0 1844 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_3_0
timestamp 1625156677
transform -1 0 1884 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_3_1
timestamp 1625156677
transform -1 0 1892 0 -1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_564
timestamp 1625156677
transform -1 0 1916 0 -1 2905
box -2 -3 26 103
use XOR2X1  XOR2X1_278
timestamp 1625156677
transform -1 0 1972 0 -1 2905
box -2 -3 58 103
use OAI21X1  OAI21X1_519
timestamp 1625156677
transform 1 0 1972 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_569
timestamp 1625156677
transform -1 0 2028 0 -1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_455
timestamp 1625156677
transform 1 0 2028 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_421
timestamp 1625156677
transform -1 0 2076 0 -1 2905
box -2 -3 18 103
use AOI21X1  AOI21X1_299
timestamp 1625156677
transform -1 0 2108 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_328
timestamp 1625156677
transform -1 0 2132 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_300
timestamp 1625156677
transform -1 0 2164 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_459
timestamp 1625156677
transform 1 0 2164 0 -1 2905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_197
timestamp 1625156677
transform -1 0 2252 0 -1 2905
box -2 -3 58 103
use OAI21X1  OAI21X1_516
timestamp 1625156677
transform -1 0 2284 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_517
timestamp 1625156677
transform 1 0 2284 0 -1 2905
box -2 -3 34 103
use BUFX2  BUFX2_227
timestamp 1625156677
transform -1 0 2340 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_423
timestamp 1625156677
transform 1 0 2340 0 -1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_355
timestamp 1625156677
transform -1 0 2380 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_4_0
timestamp 1625156677
transform 1 0 2380 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_4_1
timestamp 1625156677
transform 1 0 2388 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_561
timestamp 1625156677
transform 1 0 2396 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_467
timestamp 1625156677
transform 1 0 2428 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_603
timestamp 1625156677
transform 1 0 2444 0 -1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_331
timestamp 1625156677
transform 1 0 2468 0 -1 2905
box -2 -3 98 103
use XOR2X1  XOR2X1_284
timestamp 1625156677
transform 1 0 2564 0 -1 2905
box -2 -3 58 103
use OAI21X1  OAI21X1_559
timestamp 1625156677
transform 1 0 2620 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_354
timestamp 1625156677
transform 1 0 2652 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_598
timestamp 1625156677
transform 1 0 2676 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_599
timestamp 1625156677
transform -1 0 2724 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_558
timestamp 1625156677
transform -1 0 2756 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_482
timestamp 1625156677
transform -1 0 2788 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_464
timestamp 1625156677
transform 1 0 2788 0 -1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_483
timestamp 1625156677
transform -1 0 2836 0 -1 2905
box -2 -3 34 103
use AOI22X1  AOI22X1_22
timestamp 1625156677
transform 1 0 2836 0 -1 2905
box -2 -3 42 103
use NAND2X1  NAND2X1_600
timestamp 1625156677
transform 1 0 2876 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_5_0
timestamp 1625156677
transform 1 0 2900 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_5_1
timestamp 1625156677
transform 1 0 2908 0 -1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_321
timestamp 1625156677
transform 1 0 2916 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_607
timestamp 1625156677
transform -1 0 2972 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_557
timestamp 1625156677
transform -1 0 3004 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_602
timestamp 1625156677
transform 1 0 3004 0 -1 2905
box -2 -3 26 103
use XOR2X1  XOR2X1_296
timestamp 1625156677
transform -1 0 3084 0 -1 2905
box -2 -3 58 103
use OAI21X1  OAI21X1_563
timestamp 1625156677
transform -1 0 3116 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_353
timestamp 1625156677
transform 1 0 3116 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_320
timestamp 1625156677
transform -1 0 3172 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_484
timestamp 1625156677
transform -1 0 3204 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_556
timestamp 1625156677
transform -1 0 3236 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_597
timestamp 1625156677
transform 1 0 3236 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_456
timestamp 1625156677
transform -1 0 3276 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_550
timestamp 1625156677
transform -1 0 3308 0 -1 2905
box -2 -3 34 103
use NOR3X1  NOR3X1_85
timestamp 1625156677
transform 1 0 3308 0 -1 2905
box -2 -3 66 103
use XNOR2X1  XNOR2X1_204
timestamp 1625156677
transform -1 0 3428 0 -1 2905
box -2 -3 58 103
use FILL  FILL_28_6_0
timestamp 1625156677
transform 1 0 3428 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_6_1
timestamp 1625156677
transform 1 0 3436 0 -1 2905
box -2 -3 10 103
use INVX1  INVX1_454
timestamp 1625156677
transform 1 0 3444 0 -1 2905
box -2 -3 18 103
use AND2X2  AND2X2_155
timestamp 1625156677
transform -1 0 3492 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_592
timestamp 1625156677
transform -1 0 3516 0 -1 2905
box -2 -3 26 103
use BUFX2  BUFX2_236
timestamp 1625156677
transform -1 0 3540 0 -1 2905
box -2 -3 26 103
use XOR2X1  XOR2X1_295
timestamp 1625156677
transform -1 0 3596 0 -1 2905
box -2 -3 58 103
use NAND2X1  NAND2X1_589
timestamp 1625156677
transform 1 0 3596 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_449
timestamp 1625156677
transform 1 0 3620 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_587
timestamp 1625156677
transform 1 0 3636 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_452
timestamp 1625156677
transform 1 0 3660 0 -1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_474
timestamp 1625156677
transform 1 0 3676 0 -1 2905
box -2 -3 34 103
use XOR2X1  XOR2X1_294
timestamp 1625156677
transform -1 0 3764 0 -1 2905
box -2 -3 58 103
use AND2X2  AND2X2_153
timestamp 1625156677
transform -1 0 3796 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_450
timestamp 1625156677
transform 1 0 3796 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_543
timestamp 1625156677
transform -1 0 3844 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_312
timestamp 1625156677
transform -1 0 3876 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_311
timestamp 1625156677
transform 1 0 3876 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_446
timestamp 1625156677
transform -1 0 3924 0 -1 2905
box -2 -3 18 103
use FILL  FILL_28_7_0
timestamp 1625156677
transform -1 0 3932 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_7_1
timestamp 1625156677
transform -1 0 3940 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_537
timestamp 1625156677
transform -1 0 3972 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_578
timestamp 1625156677
transform -1 0 3996 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_575
timestamp 1625156677
transform 1 0 3996 0 -1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_463
timestamp 1625156677
transform 1 0 4020 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_531
timestamp 1625156677
transform -1 0 4084 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_437
timestamp 1625156677
transform 1 0 4084 0 -1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_471
timestamp 1625156677
transform 1 0 4100 0 -1 2905
box -2 -3 34 103
use INVX2  INVX2_72
timestamp 1625156677
transform 1 0 4132 0 -1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_337
timestamp 1625156677
transform -1 0 4172 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_532
timestamp 1625156677
transform -1 0 4204 0 -1 2905
box -2 -3 34 103
use NOR3X1  NOR3X1_84
timestamp 1625156677
transform 1 0 4204 0 -1 2905
box -2 -3 66 103
use OAI21X1  OAI21X1_529
timestamp 1625156677
transform 1 0 4268 0 -1 2905
box -2 -3 34 103
use AND2X2  AND2X2_152
timestamp 1625156677
transform 1 0 4300 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_196
timestamp 1625156677
transform 1 0 4332 0 -1 2905
box -2 -3 98 103
use FILL  FILL_28_8_0
timestamp 1625156677
transform -1 0 4436 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_8_1
timestamp 1625156677
transform -1 0 4444 0 -1 2905
box -2 -3 10 103
use XOR2X1  XOR2X1_84
timestamp 1625156677
transform -1 0 4500 0 -1 2905
box -2 -3 58 103
use BUFX2  BUFX2_243
timestamp 1625156677
transform -1 0 4524 0 -1 2905
box -2 -3 26 103
use BUFX2  BUFX2_115
timestamp 1625156677
transform -1 0 4548 0 -1 2905
box -2 -3 26 103
use OR2X2  OR2X2_74
timestamp 1625156677
transform 1 0 4548 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_169
timestamp 1625156677
transform -1 0 4612 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_119
timestamp 1625156677
transform 1 0 4612 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_170
timestamp 1625156677
transform -1 0 4676 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_164
timestamp 1625156677
transform -1 0 4708 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_162
timestamp 1625156677
transform -1 0 4740 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_171
timestamp 1625156677
transform 1 0 4740 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_113
timestamp 1625156677
transform 1 0 4772 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_121
timestamp 1625156677
transform -1 0 4828 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_167
timestamp 1625156677
transform -1 0 4860 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_110
timestamp 1625156677
transform -1 0 4884 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_166
timestamp 1625156677
transform 1 0 4884 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_112
timestamp 1625156677
transform 1 0 4916 0 -1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_173
timestamp 1625156677
transform 1 0 4932 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_9_0
timestamp 1625156677
transform 1 0 4964 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_9_1
timestamp 1625156677
transform 1 0 4972 0 -1 2905
box -2 -3 10 103
use NAND3X1  NAND3X1_172
timestamp 1625156677
transform 1 0 4980 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_122
timestamp 1625156677
transform 1 0 5012 0 -1 2905
box -2 -3 34 103
use OR2X2  OR2X2_75
timestamp 1625156677
transform -1 0 5076 0 -1 2905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1625156677
transform -1 0 5172 0 -1 2905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_197
timestamp 1625156677
transform -1 0 5268 0 -1 2905
box -2 -3 98 103
use BUFX2  BUFX2_9
timestamp 1625156677
transform 1 0 5268 0 -1 2905
box -2 -3 26 103
use BUFX2  BUFX2_132
timestamp 1625156677
transform -1 0 5316 0 -1 2905
box -2 -3 26 103
use BUFX2  BUFX2_61
timestamp 1625156677
transform -1 0 28 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_237
timestamp 1625156677
transform 1 0 28 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_348
timestamp 1625156677
transform 1 0 60 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_268
timestamp 1625156677
transform -1 0 108 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_366
timestamp 1625156677
transform -1 0 140 0 1 2705
box -2 -3 34 103
use NOR3X1  NOR3X1_65
timestamp 1625156677
transform -1 0 204 0 1 2705
box -2 -3 66 103
use NAND2X1  NAND2X1_404
timestamp 1625156677
transform 1 0 204 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_266
timestamp 1625156677
transform 1 0 228 0 1 2705
box -2 -3 18 103
use NAND3X1  NAND3X1_346
timestamp 1625156677
transform 1 0 244 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_229
timestamp 1625156677
transform -1 0 300 0 1 2705
box -2 -3 26 103
use INVX2  INVX2_63
timestamp 1625156677
transform -1 0 316 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_361
timestamp 1625156677
transform -1 0 348 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_0_0
timestamp 1625156677
transform 1 0 348 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_0_1
timestamp 1625156677
transform 1 0 356 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_358
timestamp 1625156677
transform 1 0 364 0 1 2705
box -2 -3 34 103
use NOR3X1  NOR3X1_66
timestamp 1625156677
transform 1 0 396 0 1 2705
box -2 -3 66 103
use NAND3X1  NAND3X1_345
timestamp 1625156677
transform 1 0 460 0 1 2705
box -2 -3 34 103
use AND2X2  AND2X2_115
timestamp 1625156677
transform -1 0 524 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_402
timestamp 1625156677
transform -1 0 548 0 1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_303
timestamp 1625156677
transform -1 0 644 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_300
timestamp 1625156677
transform -1 0 740 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_300
timestamp 1625156677
transform 1 0 740 0 1 2705
box -2 -3 18 103
use NAND3X1  NAND3X1_370
timestamp 1625156677
transform -1 0 788 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_297
timestamp 1625156677
transform -1 0 804 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_393
timestamp 1625156677
transform -1 0 836 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_435
timestamp 1625156677
transform 1 0 836 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_1_0
timestamp 1625156677
transform -1 0 868 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_1_1
timestamp 1625156677
transform -1 0 876 0 1 2705
box -2 -3 10 103
use BUFX2  BUFX2_209
timestamp 1625156677
transform -1 0 900 0 1 2705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_168
timestamp 1625156677
transform 1 0 900 0 1 2705
box -2 -3 58 103
use NOR2X1  NOR2X1_242
timestamp 1625156677
transform 1 0 956 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_298
timestamp 1625156677
transform 1 0 980 0 1 2705
box -2 -3 18 103
use BUFX2  BUFX2_143
timestamp 1625156677
transform 1 0 996 0 1 2705
box -2 -3 26 103
use XOR2X1  XOR2X1_198
timestamp 1625156677
transform 1 0 1020 0 1 2705
box -2 -3 58 103
use NOR3X1  NOR3X1_68
timestamp 1625156677
transform -1 0 1140 0 1 2705
box -2 -3 66 103
use NOR2X1  NOR2X1_238
timestamp 1625156677
transform -1 0 1164 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_118
timestamp 1625156677
transform -1 0 1196 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_419
timestamp 1625156677
transform -1 0 1220 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_375
timestamp 1625156677
transform 1 0 1220 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_282
timestamp 1625156677
transform -1 0 1268 0 1 2705
box -2 -3 18 103
use CLKBUF1  CLKBUF1_39
timestamp 1625156677
transform 1 0 1268 0 1 2705
box -2 -3 74 103
use FILL  FILL_27_2_0
timestamp 1625156677
transform -1 0 1348 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_2_1
timestamp 1625156677
transform -1 0 1356 0 1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_326
timestamp 1625156677
transform -1 0 1452 0 1 2705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_8
timestamp 1625156677
transform -1 0 1524 0 1 2705
box -2 -3 74 103
use BUFX4  BUFX4_5
timestamp 1625156677
transform -1 0 1556 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_363
timestamp 1625156677
transform 1 0 1556 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_554
timestamp 1625156677
transform -1 0 1668 0 1 2705
box -2 -3 18 103
use INVX1  INVX1_417
timestamp 1625156677
transform 1 0 1668 0 1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_555
timestamp 1625156677
transform 1 0 1684 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_563
timestamp 1625156677
transform -1 0 1732 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_302
timestamp 1625156677
transform 1 0 1732 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_556
timestamp 1625156677
transform 1 0 1764 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_573
timestamp 1625156677
transform -1 0 1804 0 1 2705
box -2 -3 18 103
use NAND3X1  NAND3X1_450
timestamp 1625156677
transform 1 0 1804 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_303
timestamp 1625156677
transform 1 0 1836 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_427
timestamp 1625156677
transform -1 0 1884 0 1 2705
box -2 -3 18 103
use FILL  FILL_27_3_0
timestamp 1625156677
transform -1 0 1892 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_3_1
timestamp 1625156677
transform -1 0 1900 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_512
timestamp 1625156677
transform -1 0 1932 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_559
timestamp 1625156677
transform -1 0 1956 0 1 2705
box -2 -3 26 103
use INVX2  INVX2_71
timestamp 1625156677
transform -1 0 1972 0 1 2705
box -2 -3 18 103
use INVX1  INVX1_418
timestamp 1625156677
transform 1 0 1972 0 1 2705
box -2 -3 18 103
use NAND3X1  NAND3X1_458
timestamp 1625156677
transform 1 0 1988 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_325
timestamp 1625156677
transform -1 0 2044 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_326
timestamp 1625156677
transform -1 0 2068 0 1 2705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_196
timestamp 1625156677
transform -1 0 2124 0 1 2705
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_336
timestamp 1625156677
transform -1 0 2220 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_350
timestamp 1625156677
transform 1 0 2220 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_424
timestamp 1625156677
transform 1 0 2316 0 1 2705
box -2 -3 18 103
use NAND3X1  NAND3X1_454
timestamp 1625156677
transform 1 0 2332 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_453
timestamp 1625156677
transform 1 0 2364 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_4_0
timestamp 1625156677
transform -1 0 2404 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_4_1
timestamp 1625156677
transform -1 0 2412 0 1 2705
box -2 -3 10 103
use INVX1  INVX1_422
timestamp 1625156677
transform -1 0 2428 0 1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_332
timestamp 1625156677
transform 1 0 2428 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_333
timestamp 1625156677
transform 1 0 2524 0 1 2705
box -2 -3 98 103
use INVX1  INVX1_568
timestamp 1625156677
transform -1 0 2636 0 1 2705
box -2 -3 18 103
use XOR2X1  XOR2X1_286
timestamp 1625156677
transform 1 0 2636 0 1 2705
box -2 -3 58 103
use INVX1  INVX1_463
timestamp 1625156677
transform 1 0 2692 0 1 2705
box -2 -3 18 103
use BUFX2  BUFX2_95
timestamp 1625156677
transform -1 0 2732 0 1 2705
box -2 -3 26 103
use XOR2X1  XOR2X1_283
timestamp 1625156677
transform 1 0 2732 0 1 2705
box -2 -3 58 103
use INVX1  INVX1_462
timestamp 1625156677
transform 1 0 2788 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_555
timestamp 1625156677
transform 1 0 2804 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_461
timestamp 1625156677
transform 1 0 2836 0 1 2705
box -2 -3 18 103
use NAND3X1  NAND3X1_479
timestamp 1625156677
transform -1 0 2884 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_481
timestamp 1625156677
transform 1 0 2884 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_5_0
timestamp 1625156677
transform 1 0 2916 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_5_1
timestamp 1625156677
transform 1 0 2924 0 1 2705
box -2 -3 10 103
use NAND3X1  NAND3X1_480
timestamp 1625156677
transform 1 0 2932 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_460
timestamp 1625156677
transform -1 0 2980 0 1 2705
box -2 -3 18 103
use NAND3X1  NAND3X1_485
timestamp 1625156677
transform 1 0 2980 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_352
timestamp 1625156677
transform -1 0 3036 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_316
timestamp 1625156677
transform 1 0 3036 0 1 2705
box -2 -3 34 103
use XOR2X1  XOR2X1_281
timestamp 1625156677
transform -1 0 3124 0 1 2705
box -2 -3 58 103
use AOI21X1  AOI21X1_317
timestamp 1625156677
transform 1 0 3124 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_478
timestamp 1625156677
transform 1 0 3156 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_458
timestamp 1625156677
transform -1 0 3204 0 1 2705
box -2 -3 18 103
use INVX1  INVX1_465
timestamp 1625156677
transform 1 0 3204 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_319
timestamp 1625156677
transform -1 0 3252 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_476
timestamp 1625156677
transform -1 0 3284 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_594
timestamp 1625156677
transform 1 0 3284 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_547
timestamp 1625156677
transform -1 0 3340 0 1 2705
box -2 -3 34 103
use XOR2X1  XOR2X1_272
timestamp 1625156677
transform 1 0 3340 0 1 2705
box -2 -3 58 103
use BUFX2  BUFX2_231
timestamp 1625156677
transform -1 0 3420 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_6_0
timestamp 1625156677
transform -1 0 3428 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_6_1
timestamp 1625156677
transform -1 0 3436 0 1 2705
box -2 -3 10 103
use BUFX2  BUFX2_237
timestamp 1625156677
transform -1 0 3460 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_347
timestamp 1625156677
transform -1 0 3484 0 1 2705
box -2 -3 26 103
use XOR2X1  XOR2X1_271
timestamp 1625156677
transform 1 0 3484 0 1 2705
box -2 -3 58 103
use XOR2X1  XOR2X1_273
timestamp 1625156677
transform 1 0 3540 0 1 2705
box -2 -3 58 103
use OAI21X1  OAI21X1_534
timestamp 1625156677
transform -1 0 3628 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_438
timestamp 1625156677
transform 1 0 3628 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_533
timestamp 1625156677
transform 1 0 3644 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_464
timestamp 1625156677
transform -1 0 3708 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_309
timestamp 1625156677
transform 1 0 3708 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_465
timestamp 1625156677
transform 1 0 3740 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_439
timestamp 1625156677
transform -1 0 3788 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_528
timestamp 1625156677
transform 1 0 3788 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_335
timestamp 1625156677
transform -1 0 3844 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_435
timestamp 1625156677
transform 1 0 3844 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_310
timestamp 1625156677
transform 1 0 3860 0 1 2705
box -2 -3 34 103
use XOR2X1  XOR2X1_270
timestamp 1625156677
transform 1 0 3892 0 1 2705
box -2 -3 58 103
use FILL  FILL_27_7_0
timestamp 1625156677
transform 1 0 3948 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_7_1
timestamp 1625156677
transform 1 0 3956 0 1 2705
box -2 -3 10 103
use NAND2X1  NAND2X1_573
timestamp 1625156677
transform 1 0 3964 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_151
timestamp 1625156677
transform 1 0 3988 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_462
timestamp 1625156677
transform -1 0 4052 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_334
timestamp 1625156677
transform -1 0 4076 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_572
timestamp 1625156677
transform 1 0 4076 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_571
timestamp 1625156677
transform -1 0 4124 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_434
timestamp 1625156677
transform 1 0 4124 0 1 2705
box -2 -3 18 103
use AND2X2  AND2X2_150
timestamp 1625156677
transform 1 0 4140 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_194
timestamp 1625156677
transform 1 0 4172 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_195
timestamp 1625156677
transform 1 0 4268 0 1 2705
box -2 -3 98 103
use OR2X2  OR2X2_73
timestamp 1625156677
transform 1 0 4364 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_167
timestamp 1625156677
transform -1 0 4428 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_110
timestamp 1625156677
transform 1 0 4428 0 1 2705
box -2 -3 18 103
use FILL  FILL_27_8_0
timestamp 1625156677
transform -1 0 4452 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_8_1
timestamp 1625156677
transform -1 0 4460 0 1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_108
timestamp 1625156677
transform -1 0 4484 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_161
timestamp 1625156677
transform 1 0 4484 0 1 2705
box -2 -3 34 103
use NOR3X1  NOR3X1_43
timestamp 1625156677
transform 1 0 4516 0 1 2705
box -2 -3 66 103
use NAND2X1  NAND2X1_193
timestamp 1625156677
transform 1 0 4580 0 1 2705
box -2 -3 26 103
use NAND3X1  NAND3X1_168
timestamp 1625156677
transform -1 0 4636 0 1 2705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_87
timestamp 1625156677
transform -1 0 4692 0 1 2705
box -2 -3 58 103
use NAND2X1  NAND2X1_195
timestamp 1625156677
transform 1 0 4692 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_196
timestamp 1625156677
transform -1 0 4740 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_111
timestamp 1625156677
transform -1 0 4764 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_123
timestamp 1625156677
transform 1 0 4764 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_118
timestamp 1625156677
transform 1 0 4796 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_128
timestamp 1625156677
transform -1 0 4844 0 1 2705
box -2 -3 34 103
use INVX2  INVX2_39
timestamp 1625156677
transform 1 0 4844 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_120
timestamp 1625156677
transform -1 0 4892 0 1 2705
box -2 -3 34 103
use OR2X2  OR2X2_76
timestamp 1625156677
transform 1 0 4892 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_198
timestamp 1625156677
transform -1 0 4948 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_9_0
timestamp 1625156677
transform 1 0 4948 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_9_1
timestamp 1625156677
transform 1 0 4956 0 1 2705
box -2 -3 10 103
use AOI21X1  AOI21X1_124
timestamp 1625156677
transform 1 0 4964 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_112
timestamp 1625156677
transform 1 0 4996 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_59
timestamp 1625156677
transform 1 0 5020 0 1 2705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_198
timestamp 1625156677
transform -1 0 5148 0 1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1625156677
transform -1 0 5244 0 1 2705
box -2 -3 98 103
use BUFX2  BUFX2_142
timestamp 1625156677
transform -1 0 5268 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_578
timestamp 1625156677
transform -1 0 5284 0 1 2705
box -2 -3 18 103
use BUFX2  BUFX2_49
timestamp 1625156677
transform -1 0 5308 0 1 2705
box -2 -3 26 103
use FILL  FILL_28_1
timestamp 1625156677
transform 1 0 5308 0 1 2705
box -2 -3 10 103
use BUFX2  BUFX2_77
timestamp 1625156677
transform 1 0 4 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_231
timestamp 1625156677
transform 1 0 28 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_406
timestamp 1625156677
transform -1 0 76 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_362
timestamp 1625156677
transform 1 0 76 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_267
timestamp 1625156677
transform -1 0 124 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_405
timestamp 1625156677
transform -1 0 148 0 -1 2705
box -2 -3 26 103
use NAND3X1  NAND3X1_347
timestamp 1625156677
transform -1 0 180 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_407
timestamp 1625156677
transform -1 0 204 0 -1 2705
box -2 -3 26 103
use XOR2X1  XOR2X1_211
timestamp 1625156677
transform 1 0 204 0 -1 2705
box -2 -3 58 103
use INVX1  INVX1_275
timestamp 1625156677
transform 1 0 260 0 -1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_239
timestamp 1625156677
transform -1 0 308 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_354
timestamp 1625156677
transform 1 0 308 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_0_0
timestamp 1625156677
transform -1 0 348 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_0_1
timestamp 1625156677
transform -1 0 356 0 -1 2705
box -2 -3 10 103
use AOI21X1  AOI21X1_238
timestamp 1625156677
transform -1 0 388 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_403
timestamp 1625156677
transform -1 0 412 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_411
timestamp 1625156677
transform -1 0 436 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_370
timestamp 1625156677
transform -1 0 468 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_265
timestamp 1625156677
transform -1 0 484 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_359
timestamp 1625156677
transform -1 0 516 0 -1 2705
box -2 -3 34 103
use AND2X2  AND2X2_114
timestamp 1625156677
transform -1 0 548 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_400
timestamp 1625156677
transform 1 0 548 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_401
timestamp 1625156677
transform -1 0 596 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_227
timestamp 1625156677
transform -1 0 620 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_357
timestamp 1625156677
transform 1 0 620 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_264
timestamp 1625156677
transform -1 0 668 0 -1 2705
box -2 -3 18 103
use XOR2X1  XOR2X1_215
timestamp 1625156677
transform 1 0 668 0 -1 2705
box -2 -3 58 103
use NAND2X1  NAND2X1_431
timestamp 1625156677
transform 1 0 724 0 -1 2705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_169
timestamp 1625156677
transform -1 0 804 0 -1 2705
box -2 -3 58 103
use NOR2X1  NOR2X1_248
timestamp 1625156677
transform -1 0 828 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_434
timestamp 1625156677
transform -1 0 852 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_1_0
timestamp 1625156677
transform -1 0 860 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_1_1
timestamp 1625156677
transform -1 0 868 0 -1 2705
box -2 -3 10 103
use AND2X2  AND2X2_121
timestamp 1625156677
transform -1 0 900 0 -1 2705
box -2 -3 34 103
use BUFX2  BUFX2_199
timestamp 1625156677
transform -1 0 924 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_250
timestamp 1625156677
transform -1 0 956 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_369
timestamp 1625156677
transform -1 0 988 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_299
timestamp 1625156677
transform -1 0 1004 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_391
timestamp 1625156677
transform -1 0 1036 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_426
timestamp 1625156677
transform -1 0 1060 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_248
timestamp 1625156677
transform -1 0 1092 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_379
timestamp 1625156677
transform -1 0 1124 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_367
timestamp 1625156677
transform -1 0 1156 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_285
timestamp 1625156677
transform 1 0 1156 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_241
timestamp 1625156677
transform -1 0 1196 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_380
timestamp 1625156677
transform -1 0 1228 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_377
timestamp 1625156677
transform -1 0 1260 0 -1 2705
box -2 -3 34 103
use AND2X2  AND2X2_120
timestamp 1625156677
transform 1 0 1260 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_358
timestamp 1625156677
transform 1 0 1292 0 -1 2705
box -2 -3 34 103
use AND2X2  AND2X2_119
timestamp 1625156677
transform -1 0 1356 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_421
timestamp 1625156677
transform -1 0 1380 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_2_0
timestamp 1625156677
transform -1 0 1388 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_2_1
timestamp 1625156677
transform -1 0 1396 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_312
timestamp 1625156677
transform -1 0 1492 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_315
timestamp 1625156677
transform -1 0 1588 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_307
timestamp 1625156677
transform -1 0 1684 0 -1 2705
box -2 -3 98 103
use BUFX2  BUFX2_80
timestamp 1625156677
transform -1 0 1708 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_323
timestamp 1625156677
transform 1 0 1708 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_339
timestamp 1625156677
transform 1 0 1804 0 -1 2705
box -2 -3 98 103
use FILL  FILL_26_3_0
timestamp 1625156677
transform 1 0 1900 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_3_1
timestamp 1625156677
transform 1 0 1908 0 -1 2705
box -2 -3 10 103
use INVX1  INVX1_416
timestamp 1625156677
transform 1 0 1916 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_509
timestamp 1625156677
transform -1 0 1964 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_323
timestamp 1625156677
transform 1 0 1964 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_554
timestamp 1625156677
transform 1 0 1988 0 -1 2705
box -2 -3 26 103
use AND2X2  AND2X2_147
timestamp 1625156677
transform 1 0 2012 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_449
timestamp 1625156677
transform -1 0 2076 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_513
timestamp 1625156677
transform -1 0 2108 0 -1 2705
box -2 -3 34 103
use NOR3X1  NOR3X1_82
timestamp 1625156677
transform 1 0 2108 0 -1 2705
box -2 -3 66 103
use OAI21X1  OAI21X1_510
timestamp 1625156677
transform 1 0 2172 0 -1 2705
box -2 -3 34 103
use AND2X2  AND2X2_148
timestamp 1625156677
transform 1 0 2204 0 -1 2705
box -2 -3 34 103
use AND2X2  AND2X2_146
timestamp 1625156677
transform -1 0 2268 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_552
timestamp 1625156677
transform 1 0 2268 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_415
timestamp 1625156677
transform -1 0 2308 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_322
timestamp 1625156677
transform 1 0 2308 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_553
timestamp 1625156677
transform -1 0 2356 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_508
timestamp 1625156677
transform -1 0 2388 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_4_0
timestamp 1625156677
transform 1 0 2388 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_4_1
timestamp 1625156677
transform 1 0 2396 0 -1 2705
box -2 -3 10 103
use NAND2X1  NAND2X1_680
timestamp 1625156677
transform 1 0 2404 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_368
timestamp 1625156677
transform 1 0 2428 0 -1 2705
box -2 -3 98 103
use XOR2X1  XOR2X1_261
timestamp 1625156677
transform 1 0 2524 0 -1 2705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_206
timestamp 1625156677
transform -1 0 2636 0 -1 2705
box -2 -3 58 103
use NOR2X1  NOR2X1_357
timestamp 1625156677
transform 1 0 2636 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_343
timestamp 1625156677
transform -1 0 2756 0 -1 2705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_334
timestamp 1625156677
transform -1 0 2852 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_554
timestamp 1625156677
transform 1 0 2852 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_315
timestamp 1625156677
transform 1 0 2884 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_5_0
timestamp 1625156677
transform -1 0 2924 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_5_1
timestamp 1625156677
transform -1 0 2932 0 -1 2705
box -2 -3 10 103
use INVX1  INVX1_459
timestamp 1625156677
transform -1 0 2948 0 -1 2705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_340
timestamp 1625156677
transform 1 0 2948 0 -1 2705
box -2 -3 98 103
use XOR2X1  XOR2X1_282
timestamp 1625156677
transform -1 0 3100 0 -1 2705
box -2 -3 58 103
use BUFX2  BUFX2_238
timestamp 1625156677
transform -1 0 3124 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_596
timestamp 1625156677
transform 1 0 3124 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_351
timestamp 1625156677
transform -1 0 3172 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_549
timestamp 1625156677
transform -1 0 3204 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_601
timestamp 1625156677
transform 1 0 3204 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_318
timestamp 1625156677
transform -1 0 3260 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_455
timestamp 1625156677
transform 1 0 3260 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_593
timestamp 1625156677
transform 1 0 3276 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_560
timestamp 1625156677
transform -1 0 3332 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_348
timestamp 1625156677
transform -1 0 3356 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_358
timestamp 1625156677
transform 1 0 3356 0 -1 2705
box -2 -3 98 103
use FILL  FILL_26_6_0
timestamp 1625156677
transform -1 0 3460 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_6_1
timestamp 1625156677
transform -1 0 3468 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_359
timestamp 1625156677
transform -1 0 3564 0 -1 2705
box -2 -3 98 103
use XOR2X1  XOR2X1_280
timestamp 1625156677
transform -1 0 3620 0 -1 2705
box -2 -3 58 103
use NOR2X1  NOR2X1_339
timestamp 1625156677
transform 1 0 3620 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_576
timestamp 1625156677
transform 1 0 3644 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_577
timestamp 1625156677
transform 1 0 3668 0 -1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_228
timestamp 1625156677
transform 1 0 3692 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_530
timestamp 1625156677
transform 1 0 3788 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_436
timestamp 1625156677
transform 1 0 3820 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_582
timestamp 1625156677
transform 1 0 3836 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_541
timestamp 1625156677
transform -1 0 3892 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_336
timestamp 1625156677
transform -1 0 3916 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_574
timestamp 1625156677
transform 1 0 3916 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_7_0
timestamp 1625156677
transform 1 0 3940 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_7_1
timestamp 1625156677
transform 1 0 3948 0 -1 2705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_199
timestamp 1625156677
transform 1 0 3956 0 -1 2705
box -2 -3 98 103
use OAI21X1  OAI21X1_527
timestamp 1625156677
transform 1 0 4052 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_155
timestamp 1625156677
transform 1 0 4084 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_231
timestamp 1625156677
transform -1 0 4132 0 -1 2705
box -2 -3 34 103
use NOR3X1  NOR3X1_52
timestamp 1625156677
transform 1 0 4132 0 -1 2705
box -2 -3 66 103
use AOI21X1  AOI21X1_167
timestamp 1625156677
transform -1 0 4228 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_241
timestamp 1625156677
transform 1 0 4228 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_149
timestamp 1625156677
transform -1 0 4284 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_270
timestamp 1625156677
transform -1 0 4308 0 -1 2705
box -2 -3 26 103
use AND2X2  AND2X2_81
timestamp 1625156677
transform -1 0 4340 0 -1 2705
box -2 -3 34 103
use OR2X2  OR2X2_106
timestamp 1625156677
transform -1 0 4372 0 -1 2705
box -2 -3 34 103
use INVX2  INVX2_38
timestamp 1625156677
transform 1 0 4372 0 -1 2705
box -2 -3 18 103
use BUFX2  BUFX2_88
timestamp 1625156677
transform 1 0 4388 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_192
timestamp 1625156677
transform -1 0 4436 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_8_0
timestamp 1625156677
transform 1 0 4436 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_8_1
timestamp 1625156677
transform 1 0 4444 0 -1 2705
box -2 -3 10 103
use AND2X2  AND2X2_56
timestamp 1625156677
transform 1 0 4452 0 -1 2705
box -2 -3 34 103
use XOR2X1  XOR2X1_82
timestamp 1625156677
transform -1 0 4540 0 -1 2705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_85
timestamp 1625156677
transform -1 0 4596 0 -1 2705
box -2 -3 58 103
use NAND2X1  NAND2X1_191
timestamp 1625156677
transform 1 0 4596 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_129
timestamp 1625156677
transform 1 0 4620 0 -1 2705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_86
timestamp 1625156677
transform -1 0 4708 0 -1 2705
box -2 -3 58 103
use NAND3X1  NAND3X1_183
timestamp 1625156677
transform 1 0 4708 0 -1 2705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_88
timestamp 1625156677
transform 1 0 4740 0 -1 2705
box -2 -3 58 103
use OAI21X1  OAI21X1_165
timestamp 1625156677
transform -1 0 4828 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_170
timestamp 1625156677
transform 1 0 4828 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_199
timestamp 1625156677
transform -1 0 4884 0 -1 2705
box -2 -3 26 103
use NAND3X1  NAND3X1_182
timestamp 1625156677
transform 1 0 4884 0 -1 2705
box -2 -3 34 103
use XOR2X1  XOR2X1_85
timestamp 1625156677
transform 1 0 4916 0 -1 2705
box -2 -3 58 103
use FILL  FILL_26_9_0
timestamp 1625156677
transform 1 0 4972 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_9_1
timestamp 1625156677
transform 1 0 4980 0 -1 2705
box -2 -3 10 103
use NAND3X1  NAND3X1_177
timestamp 1625156677
transform 1 0 4988 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_176
timestamp 1625156677
transform -1 0 5052 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_174
timestamp 1625156677
transform -1 0 5084 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_175
timestamp 1625156677
transform 1 0 5084 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_169
timestamp 1625156677
transform -1 0 5148 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_168
timestamp 1625156677
transform 1 0 5148 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_113
timestamp 1625156677
transform 1 0 5180 0 -1 2705
box -2 -3 18 103
use BUFX2  BUFX2_155
timestamp 1625156677
transform 1 0 5196 0 -1 2705
box -2 -3 26 103
use BUFX2  BUFX2_156
timestamp 1625156677
transform -1 0 5244 0 -1 2705
box -2 -3 26 103
use BUFX2  BUFX2_53
timestamp 1625156677
transform -1 0 5268 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_184
timestamp 1625156677
transform -1 0 5300 0 -1 2705
box -2 -3 34 103
use FILL  FILL_27_1
timestamp 1625156677
transform -1 0 5308 0 -1 2705
box -2 -3 10 103
use FILL  FILL_27_2
timestamp 1625156677
transform -1 0 5316 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_363
timestamp 1625156677
transform 1 0 4 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_232
timestamp 1625156677
transform 1 0 36 0 1 2505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_165
timestamp 1625156677
transform -1 0 116 0 1 2505
box -2 -3 58 103
use OAI21X1  OAI21X1_367
timestamp 1625156677
transform 1 0 116 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_233
timestamp 1625156677
transform 1 0 148 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_373
timestamp 1625156677
transform 1 0 172 0 1 2505
box -2 -3 34 103
use XOR2X1  XOR2X1_206
timestamp 1625156677
transform 1 0 204 0 1 2505
box -2 -3 58 103
use NAND2X1  NAND2X1_412
timestamp 1625156677
transform 1 0 260 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_240
timestamp 1625156677
transform -1 0 316 0 1 2505
box -2 -3 34 103
use XOR2X1  XOR2X1_212
timestamp 1625156677
transform 1 0 316 0 1 2505
box -2 -3 58 103
use FILL  FILL_25_0_0
timestamp 1625156677
transform 1 0 372 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_0_1
timestamp 1625156677
transform 1 0 380 0 1 2505
box -2 -3 10 103
use BUFX2  BUFX2_200
timestamp 1625156677
transform 1 0 388 0 1 2505
box -2 -3 26 103
use BUFX2  BUFX2_206
timestamp 1625156677
transform 1 0 412 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_228
timestamp 1625156677
transform 1 0 436 0 1 2505
box -2 -3 26 103
use BUFX2  BUFX2_139
timestamp 1625156677
transform -1 0 484 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_551
timestamp 1625156677
transform -1 0 500 0 1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_261
timestamp 1625156677
transform -1 0 524 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_226
timestamp 1625156677
transform 1 0 524 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_263
timestamp 1625156677
transform -1 0 564 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_356
timestamp 1625156677
transform 1 0 564 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_436
timestamp 1625156677
transform 1 0 596 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_249
timestamp 1625156677
transform -1 0 652 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_429
timestamp 1625156677
transform 1 0 652 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_386
timestamp 1625156677
transform -1 0 708 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_244
timestamp 1625156677
transform -1 0 732 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_293
timestamp 1625156677
transform -1 0 748 0 1 2505
box -2 -3 18 103
use NAND3X1  NAND3X1_366
timestamp 1625156677
transform -1 0 780 0 1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_13
timestamp 1625156677
transform -1 0 820 0 1 2505
box -2 -3 42 103
use INVX1  INVX1_295
timestamp 1625156677
transform -1 0 836 0 1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_245
timestamp 1625156677
transform 1 0 836 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_1_0
timestamp 1625156677
transform -1 0 868 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_1_1
timestamp 1625156677
transform -1 0 876 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_392
timestamp 1625156677
transform -1 0 908 0 1 2505
box -2 -3 34 103
use NOR3X1  NOR3X1_67
timestamp 1625156677
transform -1 0 972 0 1 2505
box -2 -3 66 103
use OAI21X1  OAI21X1_385
timestamp 1625156677
transform 1 0 972 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_552
timestamp 1625156677
transform -1 0 1020 0 1 2505
box -2 -3 18 103
use INVX1  INVX1_294
timestamp 1625156677
transform 1 0 1020 0 1 2505
box -2 -3 18 103
use AOI21X1  AOI21X1_247
timestamp 1625156677
transform -1 0 1068 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_423
timestamp 1625156677
transform 1 0 1068 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_359
timestamp 1625156677
transform 1 0 1092 0 1 2505
box -2 -3 34 103
use XOR2X1  XOR2X1_199
timestamp 1625156677
transform 1 0 1124 0 1 2505
box -2 -3 58 103
use INVX1  INVX1_555
timestamp 1625156677
transform -1 0 1196 0 1 2505
box -2 -3 18 103
use INVX2  INVX2_64
timestamp 1625156677
transform -1 0 1212 0 1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_285
timestamp 1625156677
transform -1 0 1308 0 1 2505
box -2 -3 98 103
use INVX1  INVX1_561
timestamp 1625156677
transform -1 0 1324 0 1 2505
box -2 -3 18 103
use INVX1  INVX1_283
timestamp 1625156677
transform 1 0 1324 0 1 2505
box -2 -3 18 103
use FILL  FILL_25_2_0
timestamp 1625156677
transform -1 0 1348 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_2_1
timestamp 1625156677
transform -1 0 1356 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_284
timestamp 1625156677
transform -1 0 1452 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_290
timestamp 1625156677
transform -1 0 1548 0 1 2505
box -2 -3 98 103
use INVX1  INVX1_560
timestamp 1625156677
transform 1 0 1548 0 1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_347
timestamp 1625156677
transform 1 0 1564 0 1 2505
box -2 -3 98 103
use OR2X2  OR2X2_137
timestamp 1625156677
transform -1 0 1692 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_427
timestamp 1625156677
transform 1 0 1692 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_569
timestamp 1625156677
transform 1 0 1716 0 1 2505
box -2 -3 18 103
use INVX1  INVX1_556
timestamp 1625156677
transform -1 0 1748 0 1 2505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_314
timestamp 1625156677
transform -1 0 1844 0 1 2505
box -2 -3 98 103
use FILL  FILL_25_3_0
timestamp 1625156677
transform 1 0 1844 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_3_1
timestamp 1625156677
transform 1 0 1852 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_351
timestamp 1625156677
transform 1 0 1860 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_282
timestamp 1625156677
transform -1 0 2052 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_335
timestamp 1625156677
transform 1 0 2052 0 1 2505
box -2 -3 98 103
use BUFX2  BUFX2_78
timestamp 1625156677
transform -1 0 2172 0 1 2505
box -2 -3 26 103
use BUFX2  BUFX2_116
timestamp 1625156677
transform 1 0 2172 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_565
timestamp 1625156677
transform 1 0 2196 0 1 2505
box -2 -3 18 103
use OR2X2  OR2X2_152
timestamp 1625156677
transform 1 0 2212 0 1 2505
box -2 -3 34 103
use OR2X2  OR2X2_146
timestamp 1625156677
transform 1 0 2244 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_344
timestamp 1625156677
transform 1 0 2276 0 1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_691
timestamp 1625156677
transform 1 0 2372 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_4_0
timestamp 1625156677
transform -1 0 2404 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_4_1
timestamp 1625156677
transform -1 0 2412 0 1 2505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_19
timestamp 1625156677
transform -1 0 2484 0 1 2505
box -2 -3 74 103
use OR2X2  OR2X2_147
timestamp 1625156677
transform 1 0 2484 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_342
timestamp 1625156677
transform -1 0 2612 0 1 2505
box -2 -3 98 103
use INVX1  INVX1_558
timestamp 1625156677
transform -1 0 2628 0 1 2505
box -2 -3 18 103
use OR2X2  OR2X2_153
timestamp 1625156677
transform 1 0 2628 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_330
timestamp 1625156677
transform -1 0 2756 0 1 2505
box -2 -3 98 103
use OR2X2  OR2X2_145
timestamp 1625156677
transform -1 0 2788 0 1 2505
box -2 -3 34 103
use OR2X2  OR2X2_135
timestamp 1625156677
transform 1 0 2788 0 1 2505
box -2 -3 34 103
use OR2X2  OR2X2_150
timestamp 1625156677
transform 1 0 2820 0 1 2505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_45
timestamp 1625156677
transform 1 0 2852 0 1 2505
box -2 -3 74 103
use FILL  FILL_25_5_0
timestamp 1625156677
transform 1 0 2924 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_5_1
timestamp 1625156677
transform 1 0 2932 0 1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_338
timestamp 1625156677
transform 1 0 2940 0 1 2505
box -2 -3 98 103
use OAI21X1  OAI21X1_553
timestamp 1625156677
transform -1 0 3068 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_457
timestamp 1625156677
transform 1 0 3068 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_552
timestamp 1625156677
transform 1 0 3084 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_595
timestamp 1625156677
transform 1 0 3116 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_477
timestamp 1625156677
transform -1 0 3172 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_357
timestamp 1625156677
transform 1 0 3172 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_179
timestamp 1625156677
transform 1 0 3268 0 1 2505
box -2 -3 98 103
use INVX1  INVX1_88
timestamp 1625156677
transform 1 0 3364 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_127
timestamp 1625156677
transform -1 0 3412 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_6_0
timestamp 1625156677
transform 1 0 3412 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_6_1
timestamp 1625156677
transform 1 0 3420 0 1 2505
box -2 -3 10 103
use NOR2X1  NOR2X1_88
timestamp 1625156677
transform 1 0 3428 0 1 2505
box -2 -3 26 103
use NOR3X1  NOR3X1_39
timestamp 1625156677
transform 1 0 3452 0 1 2505
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_354
timestamp 1625156677
transform 1 0 3516 0 1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_356
timestamp 1625156677
transform 1 0 3612 0 1 2505
box -2 -3 98 103
use INVX8  INVX8_1
timestamp 1625156677
transform -1 0 3748 0 1 2505
box -2 -3 42 103
use BUFX2  BUFX2_44
timestamp 1625156677
transform -1 0 3772 0 1 2505
box -2 -3 26 103
use BUFX2  BUFX2_33
timestamp 1625156677
transform 1 0 3772 0 1 2505
box -2 -3 26 103
use BUFX2  BUFX2_68
timestamp 1625156677
transform -1 0 3820 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_169
timestamp 1625156677
transform -1 0 3852 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_235
timestamp 1625156677
transform -1 0 3884 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_150
timestamp 1625156677
transform 1 0 3884 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_234
timestamp 1625156677
transform 1 0 3908 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_7_0
timestamp 1625156677
transform 1 0 3940 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_7_1
timestamp 1625156677
transform 1 0 3948 0 1 2505
box -2 -3 10 103
use INVX1  INVX1_156
timestamp 1625156677
transform 1 0 3956 0 1 2505
box -2 -3 18 103
use NAND3X1  NAND3X1_245
timestamp 1625156677
transform 1 0 3972 0 1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_244
timestamp 1625156677
transform -1 0 4036 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_170
timestamp 1625156677
transform -1 0 4068 0 1 2505
box -2 -3 34 103
use OR2X2  OR2X2_107
timestamp 1625156677
transform -1 0 4100 0 1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_230
timestamp 1625156677
transform 1 0 4100 0 1 2505
box -2 -3 98 103
use BUFX2  BUFX2_267
timestamp 1625156677
transform 1 0 4196 0 1 2505
box -2 -3 26 103
use BUFX2  BUFX2_165
timestamp 1625156677
transform -1 0 4244 0 1 2505
box -2 -3 26 103
use XOR2X1  XOR2X1_124
timestamp 1625156677
transform 1 0 4244 0 1 2505
box -2 -3 58 103
use XOR2X1  XOR2X1_83
timestamp 1625156677
transform -1 0 4356 0 1 2505
box -2 -3 58 103
use OR2X2  OR2X2_77
timestamp 1625156677
transform 1 0 4356 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_201
timestamp 1625156677
transform 1 0 4388 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_180
timestamp 1625156677
transform 1 0 4412 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_8_0
timestamp 1625156677
transform -1 0 4452 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_8_1
timestamp 1625156677
transform -1 0 4460 0 1 2505
box -2 -3 10 103
use NAND3X1  NAND3X1_178
timestamp 1625156677
transform -1 0 4492 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_114
timestamp 1625156677
transform 1 0 4492 0 1 2505
box -2 -3 18 103
use AND2X2  AND2X2_61
timestamp 1625156677
transform -1 0 4540 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_114
timestamp 1625156677
transform -1 0 4564 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_172
timestamp 1625156677
transform -1 0 4596 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_173
timestamp 1625156677
transform 1 0 4596 0 1 2505
box -2 -3 34 103
use BUFX2  BUFX2_268
timestamp 1625156677
transform 1 0 4628 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_179
timestamp 1625156677
transform -1 0 4684 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_203
timestamp 1625156677
transform 1 0 4684 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_130
timestamp 1625156677
transform 1 0 4708 0 1 2505
box -2 -3 34 103
use XOR2X1  XOR2X1_100
timestamp 1625156677
transform -1 0 4796 0 1 2505
box -2 -3 58 103
use AOI21X1  AOI21X1_126
timestamp 1625156677
transform 1 0 4796 0 1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_181
timestamp 1625156677
transform 1 0 4828 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_202
timestamp 1625156677
transform -1 0 4884 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_125
timestamp 1625156677
transform 1 0 4884 0 1 2505
box -2 -3 34 103
use AND2X2  AND2X2_60
timestamp 1625156677
transform -1 0 4948 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_9_0
timestamp 1625156677
transform 1 0 4948 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_9_1
timestamp 1625156677
transform 1 0 4956 0 1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_200
timestamp 1625156677
transform 1 0 4964 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_171
timestamp 1625156677
transform 1 0 4988 0 1 2505
box -2 -3 34 103
use XOR2X1  XOR2X1_105
timestamp 1625156677
transform 1 0 5020 0 1 2505
box -2 -3 58 103
use OR2X2  OR2X2_93
timestamp 1625156677
transform -1 0 5108 0 1 2505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_90
timestamp 1625156677
transform -1 0 5164 0 1 2505
box -2 -3 58 103
use OR2X2  OR2X2_65
timestamp 1625156677
transform -1 0 5196 0 1 2505
box -2 -3 34 103
use XOR2X1  XOR2X1_107
timestamp 1625156677
transform 1 0 5196 0 1 2505
box -2 -3 58 103
use NOR2X1  NOR2X1_134
timestamp 1625156677
transform -1 0 5276 0 1 2505
box -2 -3 26 103
use AND2X2  AND2X2_73
timestamp 1625156677
transform 1 0 5276 0 1 2505
box -2 -3 34 103
use FILL  FILL_26_1
timestamp 1625156677
transform 1 0 5308 0 1 2505
box -2 -3 10 103
use BUFX2  BUFX2_29
timestamp 1625156677
transform 1 0 4 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_236
timestamp 1625156677
transform -1 0 60 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_355
timestamp 1625156677
transform -1 0 92 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_269
timestamp 1625156677
transform 1 0 92 0 -1 2505
box -2 -3 18 103
use AOI21X1  AOI21X1_235
timestamp 1625156677
transform -1 0 140 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_351
timestamp 1625156677
transform -1 0 172 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_417
timestamp 1625156677
transform 1 0 172 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_241
timestamp 1625156677
transform -1 0 228 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_410
timestamp 1625156677
transform 1 0 228 0 -1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_353
timestamp 1625156677
transform -1 0 284 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_274
timestamp 1625156677
transform -1 0 300 0 -1 2505
box -2 -3 18 103
use AOI22X1  AOI22X1_12
timestamp 1625156677
transform -1 0 340 0 -1 2505
box -2 -3 42 103
use FILL  FILL_24_0_0
timestamp 1625156677
transform -1 0 348 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_0_1
timestamp 1625156677
transform -1 0 356 0 -1 2505
box -2 -3 10 103
use INVX1  INVX1_280
timestamp 1625156677
transform -1 0 372 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_372
timestamp 1625156677
transform 1 0 372 0 -1 2505
box -2 -3 34 103
use AND2X2  AND2X2_117
timestamp 1625156677
transform 1 0 404 0 -1 2505
box -2 -3 34 103
use XOR2X1  XOR2X1_213
timestamp 1625156677
transform 1 0 436 0 -1 2505
box -2 -3 58 103
use XOR2X1  XOR2X1_191
timestamp 1625156677
transform 1 0 492 0 -1 2505
box -2 -3 58 103
use BUFX2  BUFX2_192
timestamp 1625156677
transform 1 0 548 0 -1 2505
box -2 -3 26 103
use XOR2X1  XOR2X1_190
timestamp 1625156677
transform 1 0 572 0 -1 2505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_174
timestamp 1625156677
transform 1 0 628 0 -1 2505
box -2 -3 58 103
use NAND3X1  NAND3X1_368
timestamp 1625156677
transform -1 0 716 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_244
timestamp 1625156677
transform 1 0 716 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_243
timestamp 1625156677
transform 1 0 748 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_364
timestamp 1625156677
transform 1 0 780 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_288
timestamp 1625156677
transform 1 0 812 0 -1 2505
box -2 -3 18 103
use INVX1  INVX1_292
timestamp 1625156677
transform -1 0 844 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_428
timestamp 1625156677
transform 1 0 844 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_1_0
timestamp 1625156677
transform -1 0 876 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_1_1
timestamp 1625156677
transform -1 0 884 0 -1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_427
timestamp 1625156677
transform -1 0 908 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_388
timestamp 1625156677
transform -1 0 940 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_246
timestamp 1625156677
transform -1 0 964 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_283
timestamp 1625156677
transform -1 0 1060 0 -1 2505
box -2 -3 98 103
use XOR2X1  XOR2X1_200
timestamp 1625156677
transform 1 0 1060 0 -1 2505
box -2 -3 58 103
use OAI21X1  OAI21X1_378
timestamp 1625156677
transform 1 0 1116 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_240
timestamp 1625156677
transform 1 0 1148 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_422
timestamp 1625156677
transform -1 0 1196 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_284
timestamp 1625156677
transform -1 0 1212 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_389
timestamp 1625156677
transform 1 0 1212 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_246
timestamp 1625156677
transform -1 0 1276 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_430
timestamp 1625156677
transform -1 0 1300 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_376
timestamp 1625156677
transform -1 0 1332 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_239
timestamp 1625156677
transform -1 0 1356 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_2_0
timestamp 1625156677
transform -1 0 1364 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_2_1
timestamp 1625156677
transform -1 0 1372 0 -1 2505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_23
timestamp 1625156677
transform -1 0 1444 0 -1 2505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_32
timestamp 1625156677
transform 1 0 1444 0 -1 2505
box -2 -3 74 103
use OR2X2  OR2X2_136
timestamp 1625156677
transform 1 0 1516 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_521
timestamp 1625156677
transform -1 0 1580 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_684
timestamp 1625156677
transform 1 0 1580 0 -1 2505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_2
timestamp 1625156677
transform 1 0 1604 0 -1 2505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_292
timestamp 1625156677
transform -1 0 1772 0 -1 2505
box -2 -3 98 103
use NOR2X1  NOR2X1_428
timestamp 1625156677
transform 1 0 1772 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_677
timestamp 1625156677
transform -1 0 1820 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_348
timestamp 1625156677
transform -1 0 1916 0 -1 2505
box -2 -3 98 103
use FILL  FILL_24_3_0
timestamp 1625156677
transform 1 0 1916 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_3_1
timestamp 1625156677
transform 1 0 1924 0 -1 2505
box -2 -3 10 103
use INVX1  INVX1_537
timestamp 1625156677
transform 1 0 1932 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_685
timestamp 1625156677
transform 1 0 1948 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_676
timestamp 1625156677
transform -1 0 1996 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_692
timestamp 1625156677
transform 1 0 1996 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_681
timestamp 1625156677
transform 1 0 2020 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_367
timestamp 1625156677
transform 1 0 2044 0 -1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_682
timestamp 1625156677
transform 1 0 2140 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_345
timestamp 1625156677
transform 1 0 2164 0 -1 2505
box -2 -3 98 103
use OR2X2  OR2X2_151
timestamp 1625156677
transform 1 0 2260 0 -1 2505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_364
timestamp 1625156677
transform 1 0 2292 0 -1 2505
box -2 -3 98 103
use FILL  FILL_24_4_0
timestamp 1625156677
transform 1 0 2388 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_4_1
timestamp 1625156677
transform 1 0 2396 0 -1 2505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_369
timestamp 1625156677
transform 1 0 2404 0 -1 2505
box -2 -3 98 103
use NAND3X1  NAND3X1_524
timestamp 1625156677
transform -1 0 2532 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_687
timestamp 1625156677
transform 1 0 2532 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_346
timestamp 1625156677
transform -1 0 2652 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_366
timestamp 1625156677
transform 1 0 2652 0 -1 2505
box -2 -3 98 103
use OR2X2  OR2X2_148
timestamp 1625156677
transform 1 0 2748 0 -1 2505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_40
timestamp 1625156677
transform 1 0 2780 0 -1 2505
box -2 -3 74 103
use NAND2X1  NAND2X1_683
timestamp 1625156677
transform 1 0 2852 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_5_0
timestamp 1625156677
transform 1 0 2876 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_5_1
timestamp 1625156677
transform 1 0 2884 0 -1 2505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_51
timestamp 1625156677
transform 1 0 2892 0 -1 2505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_341
timestamp 1625156677
transform 1 0 2964 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_355
timestamp 1625156677
transform 1 0 3060 0 -1 2505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_362
timestamp 1625156677
transform 1 0 3156 0 -1 2505
box -2 -3 98 103
use BUFX2  BUFX2_96
timestamp 1625156677
transform -1 0 3276 0 -1 2505
box -2 -3 26 103
use XOR2X1  XOR2X1_63
timestamp 1625156677
transform 1 0 3276 0 -1 2505
box -2 -3 58 103
use NAND2X1  NAND2X1_154
timestamp 1625156677
transform 1 0 3332 0 -1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_131
timestamp 1625156677
transform 1 0 3356 0 -1 2505
box -2 -3 34 103
use OR2X2  OR2X2_57
timestamp 1625156677
transform -1 0 3420 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_6_0
timestamp 1625156677
transform 1 0 3420 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_6_1
timestamp 1625156677
transform 1 0 3428 0 -1 2505
box -2 -3 10 103
use AND2X2  AND2X2_44
timestamp 1625156677
transform 1 0 3436 0 -1 2505
box -2 -3 34 103
use OR2X2  OR2X2_105
timestamp 1625156677
transform 1 0 3468 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_239
timestamp 1625156677
transform -1 0 3532 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_268
timestamp 1625156677
transform -1 0 3556 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_154
timestamp 1625156677
transform 1 0 3556 0 -1 2505
box -2 -3 18 103
use AND2X2  AND2X2_80
timestamp 1625156677
transform 1 0 3572 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_229
timestamp 1625156677
transform -1 0 3636 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_148
timestamp 1625156677
transform -1 0 3660 0 -1 2505
box -2 -3 26 103
use NOR3X1  NOR3X1_51
timestamp 1625156677
transform 1 0 3660 0 -1 2505
box -2 -3 66 103
use NAND3X1  NAND3X1_255
timestamp 1625156677
transform 1 0 3724 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_232
timestamp 1625156677
transform -1 0 3788 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_230
timestamp 1625156677
transform 1 0 3788 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_271
timestamp 1625156677
transform -1 0 3844 0 -1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_242
timestamp 1625156677
transform -1 0 3876 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_243
timestamp 1625156677
transform 1 0 3876 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_171
timestamp 1625156677
transform 1 0 3908 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_7_0
timestamp 1625156677
transform -1 0 3948 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_7_1
timestamp 1625156677
transform -1 0 3956 0 -1 2505
box -2 -3 10 103
use NOR2X1  NOR2X1_153
timestamp 1625156677
transform -1 0 3980 0 -1 2505
box -2 -3 26 103
use AND2X2  AND2X2_82
timestamp 1625156677
transform -1 0 4012 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_168
timestamp 1625156677
transform -1 0 4044 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_247
timestamp 1625156677
transform 1 0 4044 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_273
timestamp 1625156677
transform -1 0 4100 0 -1 2505
box -2 -3 26 103
use XOR2X1  XOR2X1_125
timestamp 1625156677
transform -1 0 4156 0 -1 2505
box -2 -3 58 103
use OAI21X1  OAI21X1_237
timestamp 1625156677
transform -1 0 4188 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_236
timestamp 1625156677
transform -1 0 4220 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_152
timestamp 1625156677
transform -1 0 4244 0 -1 2505
box -2 -3 26 103
use AND2X2  AND2X2_83
timestamp 1625156677
transform -1 0 4276 0 -1 2505
box -2 -3 34 103
use BUFX2  BUFX2_163
timestamp 1625156677
transform 1 0 4276 0 -1 2505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_214
timestamp 1625156677
transform 1 0 4300 0 -1 2505
box -2 -3 98 103
use NAND2X1  NAND2X1_206
timestamp 1625156677
transform -1 0 4420 0 -1 2505
box -2 -3 26 103
use OR2X2  OR2X2_80
timestamp 1625156677
transform 1 0 4420 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_8_0
timestamp 1625156677
transform 1 0 4452 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_8_1
timestamp 1625156677
transform 1 0 4460 0 -1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_207
timestamp 1625156677
transform 1 0 4468 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_119
timestamp 1625156677
transform 1 0 4492 0 -1 2505
box -2 -3 18 103
use INVX1  INVX1_120
timestamp 1625156677
transform 1 0 4508 0 -1 2505
box -2 -3 18 103
use NAND3X1  NAND3X1_184
timestamp 1625156677
transform 1 0 4524 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_177
timestamp 1625156677
transform -1 0 4588 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_117
timestamp 1625156677
transform 1 0 4588 0 -1 2505
box -2 -3 18 103
use AOI21X1  AOI21X1_127
timestamp 1625156677
transform -1 0 4636 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_176
timestamp 1625156677
transform -1 0 4668 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_117
timestamp 1625156677
transform 1 0 4668 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_116
timestamp 1625156677
transform 1 0 4692 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_174
timestamp 1625156677
transform -1 0 4748 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_115
timestamp 1625156677
transform -1 0 4772 0 -1 2505
box -2 -3 26 103
use INVX1  INVX1_115
timestamp 1625156677
transform -1 0 4788 0 -1 2505
box -2 -3 18 103
use OR2X2  OR2X2_78
timestamp 1625156677
transform 1 0 4788 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_175
timestamp 1625156677
transform -1 0 4852 0 -1 2505
box -2 -3 34 103
use INVX2  INVX2_40
timestamp 1625156677
transform -1 0 4868 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_208
timestamp 1625156677
transform 1 0 4868 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_235
timestamp 1625156677
transform -1 0 4916 0 -1 2505
box -2 -3 26 103
use OR2X2  OR2X2_91
timestamp 1625156677
transform -1 0 4948 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_9_0
timestamp 1625156677
transform -1 0 4956 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_9_1
timestamp 1625156677
transform -1 0 4964 0 -1 2505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_89
timestamp 1625156677
transform -1 0 5020 0 -1 2505
box -2 -3 58 103
use NAND2X1  NAND2X1_239
timestamp 1625156677
transform 1 0 5020 0 -1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_216
timestamp 1625156677
transform -1 0 5076 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_214
timestamp 1625156677
transform -1 0 5108 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_215
timestamp 1625156677
transform -1 0 5140 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_136
timestamp 1625156677
transform 1 0 5140 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_206
timestamp 1625156677
transform -1 0 5188 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_207
timestamp 1625156677
transform -1 0 5220 0 -1 2505
box -2 -3 34 103
use BUFX2  BUFX2_150
timestamp 1625156677
transform -1 0 5244 0 -1 2505
box -2 -3 26 103
use BUFX2  BUFX2_100
timestamp 1625156677
transform 1 0 5244 0 -1 2505
box -2 -3 26 103
use OR2X2  OR2X2_83
timestamp 1625156677
transform -1 0 5300 0 -1 2505
box -2 -3 34 103
use FILL  FILL_25_1
timestamp 1625156677
transform -1 0 5308 0 -1 2505
box -2 -3 10 103
use FILL  FILL_25_2
timestamp 1625156677
transform -1 0 5316 0 -1 2505
box -2 -3 10 103
use INVX1  INVX1_271
timestamp 1625156677
transform -1 0 20 0 1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_350
timestamp 1625156677
transform -1 0 52 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_272
timestamp 1625156677
transform 1 0 52 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_365
timestamp 1625156677
transform -1 0 100 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_349
timestamp 1625156677
transform -1 0 132 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_270
timestamp 1625156677
transform -1 0 148 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_364
timestamp 1625156677
transform 1 0 148 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_352
timestamp 1625156677
transform -1 0 212 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_368
timestamp 1625156677
transform 1 0 212 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_273
timestamp 1625156677
transform -1 0 260 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_369
timestamp 1625156677
transform 1 0 260 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_356
timestamp 1625156677
transform -1 0 324 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_242
timestamp 1625156677
transform 1 0 324 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_0_0
timestamp 1625156677
transform 1 0 356 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_0_1
timestamp 1625156677
transform 1 0 364 0 1 2305
box -2 -3 10 103
use INVX1  INVX1_279
timestamp 1625156677
transform 1 0 372 0 1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_416
timestamp 1625156677
transform 1 0 388 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_278
timestamp 1625156677
transform 1 0 412 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_374
timestamp 1625156677
transform 1 0 428 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_418
timestamp 1625156677
transform 1 0 460 0 1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_357
timestamp 1625156677
transform 1 0 484 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_281
timestamp 1625156677
transform 1 0 516 0 1 2305
box -2 -3 18 103
use XOR2X1  XOR2X1_189
timestamp 1625156677
transform 1 0 532 0 1 2305
box -2 -3 58 103
use INVX1  INVX1_290
timestamp 1625156677
transform 1 0 588 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_289
timestamp 1625156677
transform -1 0 620 0 1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_363
timestamp 1625156677
transform -1 0 652 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_362
timestamp 1625156677
transform 1 0 652 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_384
timestamp 1625156677
transform 1 0 684 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_291
timestamp 1625156677
transform -1 0 732 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_383
timestamp 1625156677
transform 1 0 732 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_365
timestamp 1625156677
transform 1 0 764 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_387
timestamp 1625156677
transform 1 0 796 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_1_0
timestamp 1625156677
transform -1 0 836 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_1_1
timestamp 1625156677
transform -1 0 844 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_295
timestamp 1625156677
transform -1 0 940 0 1 2305
box -2 -3 98 103
use INVX1  INVX1_546
timestamp 1625156677
transform -1 0 956 0 1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_245
timestamp 1625156677
transform 1 0 956 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_361
timestamp 1625156677
transform 1 0 988 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_287
timestamp 1625156677
transform -1 0 1036 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_243
timestamp 1625156677
transform -1 0 1060 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_425
timestamp 1625156677
transform -1 0 1084 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_424
timestamp 1625156677
transform -1 0 1108 0 1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_360
timestamp 1625156677
transform -1 0 1140 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_381
timestamp 1625156677
transform 1 0 1140 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_286
timestamp 1625156677
transform -1 0 1188 0 1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_294
timestamp 1625156677
transform -1 0 1284 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_291
timestamp 1625156677
transform -1 0 1380 0 1 2305
box -2 -3 98 103
use FILL  FILL_23_2_0
timestamp 1625156677
transform -1 0 1388 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_2_1
timestamp 1625156677
transform -1 0 1396 0 1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_287
timestamp 1625156677
transform -1 0 1492 0 1 2305
box -2 -3 98 103
use AOI21X1  AOI21X1_380
timestamp 1625156677
transform 1 0 1492 0 1 2305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_240
timestamp 1625156677
transform 1 0 1524 0 1 2305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_242
timestamp 1625156677
transform -1 0 1636 0 1 2305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_210
timestamp 1625156677
transform 1 0 1636 0 1 2305
box -2 -3 58 103
use NAND3X1  NAND3X1_516
timestamp 1625156677
transform -1 0 1724 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_652
timestamp 1625156677
transform 1 0 1724 0 1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_505
timestamp 1625156677
transform 1 0 1748 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_570
timestamp 1625156677
transform -1 0 1796 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_536
timestamp 1625156677
transform 1 0 1796 0 1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_518
timestamp 1625156677
transform -1 0 1844 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_376
timestamp 1625156677
transform 1 0 1844 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_3_0
timestamp 1625156677
transform 1 0 1876 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_3_1
timestamp 1625156677
transform 1 0 1884 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_612
timestamp 1625156677
transform 1 0 1892 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_381
timestamp 1625156677
transform -1 0 1956 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_522
timestamp 1625156677
transform 1 0 1956 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_517
timestamp 1625156677
transform -1 0 2020 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_572
timestamp 1625156677
transform -1 0 2036 0 1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_352
timestamp 1625156677
transform 1 0 2036 0 1 2305
box -2 -3 98 103
use XNOR2X1  XNOR2X1_238
timestamp 1625156677
transform 1 0 2132 0 1 2305
box -2 -3 58 103
use AOI21X1  AOI21X1_383
timestamp 1625156677
transform -1 0 2220 0 1 2305
box -2 -3 34 103
use OR2X2  OR2X2_138
timestamp 1625156677
transform 1 0 2220 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_361
timestamp 1625156677
transform 1 0 2252 0 1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_668
timestamp 1625156677
transform 1 0 2348 0 1 2305
box -2 -3 26 103
use BUFX2  BUFX2_73
timestamp 1625156677
transform 1 0 2372 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_4_0
timestamp 1625156677
transform -1 0 2404 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_4_1
timestamp 1625156677
transform -1 0 2412 0 1 2305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_22
timestamp 1625156677
transform -1 0 2484 0 1 2305
box -2 -3 74 103
use BUFX4  BUFX4_4
timestamp 1625156677
transform -1 0 2516 0 1 2305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_360
timestamp 1625156677
transform 1 0 2516 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_246
timestamp 1625156677
transform 1 0 2612 0 1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_180
timestamp 1625156677
transform 1 0 2708 0 1 2305
box -2 -3 98 103
use NAND3X1  NAND3X1_520
timestamp 1625156677
transform -1 0 2836 0 1 2305
box -2 -3 34 103
use OR2X2  OR2X2_58
timestamp 1625156677
transform 1 0 2836 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_133
timestamp 1625156677
transform 1 0 2868 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_5_0
timestamp 1625156677
transform 1 0 2900 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_5_1
timestamp 1625156677
transform 1 0 2908 0 1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_95
timestamp 1625156677
transform 1 0 2916 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_89
timestamp 1625156677
transform 1 0 2948 0 1 2305
box -2 -3 18 103
use AND2X2  AND2X2_45
timestamp 1625156677
transform 1 0 2964 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_89
timestamp 1625156677
transform -1 0 3020 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_129
timestamp 1625156677
transform 1 0 3020 0 1 2305
box -2 -3 34 103
use NOR3X1  NOR3X1_40
timestamp 1625156677
transform 1 0 3052 0 1 2305
box -2 -3 66 103
use NAND2X1  NAND2X1_158
timestamp 1625156677
transform 1 0 3116 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_99
timestamp 1625156677
transform -1 0 3172 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_93
timestamp 1625156677
transform 1 0 3172 0 1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_135
timestamp 1625156677
transform 1 0 3196 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_134
timestamp 1625156677
transform -1 0 3260 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_130
timestamp 1625156677
transform -1 0 3292 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_157
timestamp 1625156677
transform 1 0 3292 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_128
timestamp 1625156677
transform 1 0 3316 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_132
timestamp 1625156677
transform 1 0 3348 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_155
timestamp 1625156677
transform -1 0 3404 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_6_0
timestamp 1625156677
transform -1 0 3412 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_6_1
timestamp 1625156677
transform -1 0 3420 0 1 2305
box -2 -3 10 103
use XNOR2X1  XNOR2X1_69
timestamp 1625156677
transform -1 0 3476 0 1 2305
box -2 -3 58 103
use NAND2X1  NAND2X1_269
timestamp 1625156677
transform -1 0 3500 0 1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_240
timestamp 1625156677
transform -1 0 3532 0 1 2305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_124
timestamp 1625156677
transform -1 0 3588 0 1 2305
box -2 -3 58 103
use XOR2X1  XOR2X1_140
timestamp 1625156677
transform 1 0 3588 0 1 2305
box -2 -3 58 103
use OAI21X1  OAI21X1_233
timestamp 1625156677
transform -1 0 3676 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_272
timestamp 1625156677
transform 1 0 3676 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_238
timestamp 1625156677
transform 1 0 3700 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_275
timestamp 1625156677
transform -1 0 3756 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_178
timestamp 1625156677
transform -1 0 3788 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_51
timestamp 1625156677
transform -1 0 3804 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_151
timestamp 1625156677
transform -1 0 3828 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_176
timestamp 1625156677
transform -1 0 3860 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_162
timestamp 1625156677
transform -1 0 3876 0 1 2305
box -2 -3 18 103
use AND2X2  AND2X2_84
timestamp 1625156677
transform -1 0 3908 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_276
timestamp 1625156677
transform -1 0 3932 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_7_0
timestamp 1625156677
transform -1 0 3940 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_7_1
timestamp 1625156677
transform -1 0 3948 0 1 2305
box -2 -3 10 103
use NAND3X1  NAND3X1_249
timestamp 1625156677
transform -1 0 3980 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_248
timestamp 1625156677
transform -1 0 4012 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_172
timestamp 1625156677
transform -1 0 4044 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_246
timestamp 1625156677
transform -1 0 4076 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_274
timestamp 1625156677
transform 1 0 4076 0 1 2305
box -2 -3 26 103
use OR2X2  OR2X2_108
timestamp 1625156677
transform -1 0 4132 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_157
timestamp 1625156677
transform -1 0 4148 0 1 2305
box -2 -3 18 103
use BUFX2  BUFX2_166
timestamp 1625156677
transform -1 0 4172 0 1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_212
timestamp 1625156677
transform 1 0 4172 0 1 2305
box -2 -3 98 103
use INVX1  INVX1_133
timestamp 1625156677
transform 1 0 4268 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_129
timestamp 1625156677
transform 1 0 4284 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_197
timestamp 1625156677
transform -1 0 4340 0 1 2305
box -2 -3 34 103
use NOR3X1  NOR3X1_48
timestamp 1625156677
transform 1 0 4340 0 1 2305
box -2 -3 66 103
use AND2X2  AND2X2_69
timestamp 1625156677
transform -1 0 4436 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_8_0
timestamp 1625156677
transform 1 0 4436 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_8_1
timestamp 1625156677
transform 1 0 4444 0 1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_232
timestamp 1625156677
transform 1 0 4452 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_143
timestamp 1625156677
transform -1 0 4508 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_205
timestamp 1625156677
transform 1 0 4508 0 1 2305
box -2 -3 34 103
use OR2X2  OR2X2_90
timestamp 1625156677
transform -1 0 4572 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_209
timestamp 1625156677
transform 1 0 4572 0 1 2305
box -2 -3 26 103
use XOR2X1  XOR2X1_104
timestamp 1625156677
transform -1 0 4652 0 1 2305
box -2 -3 58 103
use AOI21X1  AOI21X1_145
timestamp 1625156677
transform -1 0 4684 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_144
timestamp 1625156677
transform -1 0 4716 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_208
timestamp 1625156677
transform -1 0 4748 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_209
timestamp 1625156677
transform -1 0 4780 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_134
timestamp 1625156677
transform -1 0 4796 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_200
timestamp 1625156677
transform -1 0 4828 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_201
timestamp 1625156677
transform -1 0 4860 0 1 2305
box -2 -3 34 103
use AND2X2  AND2X2_70
timestamp 1625156677
transform -1 0 4892 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_130
timestamp 1625156677
transform -1 0 4916 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_146
timestamp 1625156677
transform 1 0 4916 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_9_0
timestamp 1625156677
transform -1 0 4956 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_9_1
timestamp 1625156677
transform -1 0 4964 0 1 2305
box -2 -3 10 103
use AND2X2  AND2X2_72
timestamp 1625156677
transform -1 0 4996 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_238
timestamp 1625156677
transform -1 0 5020 0 1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_213
timestamp 1625156677
transform -1 0 5052 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_212
timestamp 1625156677
transform 1 0 5052 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_211
timestamp 1625156677
transform 1 0 5084 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_210
timestamp 1625156677
transform -1 0 5148 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_135
timestamp 1625156677
transform 1 0 5148 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_203
timestamp 1625156677
transform -1 0 5196 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_202
timestamp 1625156677
transform -1 0 5228 0 1 2305
box -2 -3 34 103
use BUFX2  BUFX2_27
timestamp 1625156677
transform 1 0 5228 0 1 2305
box -2 -3 26 103
use BUFX2  BUFX2_37
timestamp 1625156677
transform 1 0 5252 0 1 2305
box -2 -3 26 103
use AND2X2  AND2X2_66
timestamp 1625156677
transform -1 0 5308 0 1 2305
box -2 -3 34 103
use FILL  FILL_24_1
timestamp 1625156677
transform 1 0 5308 0 1 2305
box -2 -3 10 103
use XOR2X1  XOR2X1_192
timestamp 1625156677
transform -1 0 60 0 -1 2305
box -2 -3 58 103
use BUFX2  BUFX2_110
timestamp 1625156677
transform 1 0 60 0 -1 2305
box -2 -3 26 103
use BUFX2  BUFX2_191
timestamp 1625156677
transform -1 0 108 0 -1 2305
box -2 -3 26 103
use XOR2X1  XOR2X1_202
timestamp 1625156677
transform 1 0 108 0 -1 2305
box -2 -3 58 103
use NOR2X1  NOR2X1_234
timestamp 1625156677
transform -1 0 188 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_408
timestamp 1625156677
transform -1 0 212 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_409
timestamp 1625156677
transform -1 0 236 0 -1 2305
box -2 -3 26 103
use XOR2X1  XOR2X1_203
timestamp 1625156677
transform 1 0 236 0 -1 2305
box -2 -3 58 103
use BUFX2  BUFX2_193
timestamp 1625156677
transform -1 0 316 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_276
timestamp 1625156677
transform 1 0 316 0 -1 2305
box -2 -3 18 103
use FILL  FILL_22_0_0
timestamp 1625156677
transform -1 0 340 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_0_1
timestamp 1625156677
transform -1 0 348 0 -1 2305
box -2 -3 10 103
use AND2X2  AND2X2_112
timestamp 1625156677
transform -1 0 380 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_415
timestamp 1625156677
transform 1 0 380 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_236
timestamp 1625156677
transform 1 0 404 0 -1 2305
box -2 -3 26 103
use XOR2X1  XOR2X1_204
timestamp 1625156677
transform -1 0 484 0 -1 2305
box -2 -3 58 103
use XOR2X1  XOR2X1_214
timestamp 1625156677
transform 1 0 484 0 -1 2305
box -2 -3 58 103
use NOR2X1  NOR2X1_247
timestamp 1625156677
transform 1 0 540 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_390
timestamp 1625156677
transform 1 0 564 0 -1 2305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_171
timestamp 1625156677
transform -1 0 652 0 -1 2305
box -2 -3 58 103
use NAND2X1  NAND2X1_433
timestamp 1625156677
transform 1 0 652 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_432
timestamp 1625156677
transform -1 0 700 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_296
timestamp 1625156677
transform -1 0 716 0 -1 2305
box -2 -3 18 103
use BUFX2  BUFX2_41
timestamp 1625156677
transform -1 0 740 0 -1 2305
box -2 -3 26 103
use BUFX2  BUFX2_36
timestamp 1625156677
transform -1 0 764 0 -1 2305
box -2 -3 26 103
use BUFX2  BUFX2_103
timestamp 1625156677
transform 1 0 764 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_320
timestamp 1625156677
transform -1 0 884 0 -1 2305
box -2 -3 98 103
use FILL  FILL_22_1_0
timestamp 1625156677
transform -1 0 892 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_1_1
timestamp 1625156677
transform -1 0 900 0 -1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_382
timestamp 1625156677
transform -1 0 924 0 -1 2305
box -2 -3 26 103
use XOR2X1  XOR2X1_201
timestamp 1625156677
transform 1 0 924 0 -1 2305
box -2 -3 58 103
use OAI21X1  OAI21X1_382
timestamp 1625156677
transform 1 0 980 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_670
timestamp 1625156677
transform -1 0 1036 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_286
timestamp 1625156677
transform -1 0 1132 0 -1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_313
timestamp 1625156677
transform -1 0 1228 0 -1 2305
box -2 -3 98 103
use XNOR2X1  XNOR2X1_209
timestamp 1625156677
transform 1 0 1228 0 -1 2305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_236
timestamp 1625156677
transform 1 0 1284 0 -1 2305
box -2 -3 58 103
use NAND2X1  NAND2X1_651
timestamp 1625156677
transform 1 0 1340 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_2_0
timestamp 1625156677
transform 1 0 1364 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_2_1
timestamp 1625156677
transform 1 0 1372 0 -1 2305
box -2 -3 10 103
use NAND3X1  NAND3X1_504
timestamp 1625156677
transform 1 0 1380 0 -1 2305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_220
timestamp 1625156677
transform 1 0 1412 0 -1 2305
box -2 -3 58 103
use NAND2X1  NAND2X1_664
timestamp 1625156677
transform -1 0 1492 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_559
timestamp 1625156677
transform -1 0 1508 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_663
timestamp 1625156677
transform 1 0 1508 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_591
timestamp 1625156677
transform 1 0 1532 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_352
timestamp 1625156677
transform 1 0 1564 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_495
timestamp 1625156677
transform -1 0 1612 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_686
timestamp 1625156677
transform -1 0 1636 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_296
timestamp 1625156677
transform -1 0 1732 0 -1 2305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_337
timestamp 1625156677
transform -1 0 1828 0 -1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_673
timestamp 1625156677
transform -1 0 1852 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_388
timestamp 1625156677
transform 1 0 1852 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_3_0
timestamp 1625156677
transform -1 0 1892 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_3_1
timestamp 1625156677
transform -1 0 1900 0 -1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_674
timestamp 1625156677
transform -1 0 1924 0 -1 2305
box -2 -3 26 103
use OR2X2  OR2X2_139
timestamp 1625156677
transform -1 0 1956 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_665
timestamp 1625156677
transform 1 0 1956 0 -1 2305
box -2 -3 26 103
use BUFX2  BUFX2_260
timestamp 1625156677
transform -1 0 2004 0 -1 2305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_221
timestamp 1625156677
transform 1 0 2004 0 -1 2305
box -2 -3 58 103
use AOI21X1  AOI21X1_372
timestamp 1625156677
transform 1 0 2060 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_609
timestamp 1625156677
transform 1 0 2092 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_531
timestamp 1625156677
transform -1 0 2140 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_654
timestamp 1625156677
transform -1 0 2164 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_507
timestamp 1625156677
transform -1 0 2196 0 -1 2305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_223
timestamp 1625156677
transform 1 0 2196 0 -1 2305
box -2 -3 58 103
use NAND2X1  NAND2X1_669
timestamp 1625156677
transform -1 0 2276 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_564
timestamp 1625156677
transform -1 0 2292 0 -1 2305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_21
timestamp 1625156677
transform -1 0 2364 0 -1 2305
box -2 -3 74 103
use INVX1  INVX1_504
timestamp 1625156677
transform 1 0 2364 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_649
timestamp 1625156677
transform 1 0 2380 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_4_0
timestamp 1625156677
transform 1 0 2404 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_4_1
timestamp 1625156677
transform 1 0 2412 0 -1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_182
timestamp 1625156677
transform 1 0 2420 0 -1 2305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_18
timestamp 1625156677
transform 1 0 2516 0 -1 2305
box -2 -3 74 103
use XNOR2X1  XNOR2X1_239
timestamp 1625156677
transform 1 0 2588 0 -1 2305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_178
timestamp 1625156677
transform 1 0 2644 0 -1 2305
box -2 -3 98 103
use INVX2  INVX2_32
timestamp 1625156677
transform 1 0 2740 0 -1 2305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_227
timestamp 1625156677
transform 1 0 2756 0 -1 2305
box -2 -3 98 103
use NAND2X1  NAND2X1_156
timestamp 1625156677
transform 1 0 2852 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_96
timestamp 1625156677
transform -1 0 2908 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_5_0
timestamp 1625156677
transform -1 0 2916 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_5_1
timestamp 1625156677
transform -1 0 2924 0 -1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_104
timestamp 1625156677
transform -1 0 2956 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_96
timestamp 1625156677
transform -1 0 2972 0 -1 2305
box -2 -3 18 103
use INVX2  INVX2_33
timestamp 1625156677
transform -1 0 2988 0 -1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_91
timestamp 1625156677
transform -1 0 3012 0 -1 2305
box -2 -3 26 103
use XOR2X1  XOR2X1_80
timestamp 1625156677
transform -1 0 3068 0 -1 2305
box -2 -3 58 103
use OAI21X1  OAI21X1_131
timestamp 1625156677
transform -1 0 3100 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_97
timestamp 1625156677
transform -1 0 3132 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_136
timestamp 1625156677
transform 1 0 3132 0 -1 2305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_123
timestamp 1625156677
transform 1 0 3164 0 -1 2305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_70
timestamp 1625156677
transform -1 0 3276 0 -1 2305
box -2 -3 58 103
use NAND3X1  NAND3X1_147
timestamp 1625156677
transform -1 0 3308 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_105
timestamp 1625156677
transform -1 0 3340 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_153
timestamp 1625156677
transform 1 0 3340 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_267
timestamp 1625156677
transform 1 0 3364 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_177
timestamp 1625156677
transform 1 0 3388 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_6_0
timestamp 1625156677
transform 1 0 3420 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_6_1
timestamp 1625156677
transform 1 0 3428 0 -1 2305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_229
timestamp 1625156677
transform 1 0 3436 0 -1 2305
box -2 -3 98 103
use XOR2X1  XOR2X1_123
timestamp 1625156677
transform -1 0 3588 0 -1 2305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_125
timestamp 1625156677
transform 1 0 3588 0 -1 2305
box -2 -3 58 103
use NAND2X1  NAND2X1_284
timestamp 1625156677
transform -1 0 3668 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_242
timestamp 1625156677
transform 1 0 3668 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_254
timestamp 1625156677
transform -1 0 3732 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_239
timestamp 1625156677
transform 1 0 3732 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_173
timestamp 1625156677
transform -1 0 3796 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_278
timestamp 1625156677
transform -1 0 3820 0 -1 2305
box -2 -3 26 103
use INVX2  INVX2_52
timestamp 1625156677
transform 1 0 3820 0 -1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_155
timestamp 1625156677
transform -1 0 3860 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_159
timestamp 1625156677
transform -1 0 3876 0 -1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_174
timestamp 1625156677
transform -1 0 3908 0 -1 2305
box -2 -3 34 103
use OR2X2  OR2X2_110
timestamp 1625156677
transform -1 0 3940 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_7_0
timestamp 1625156677
transform -1 0 3948 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_7_1
timestamp 1625156677
transform -1 0 3956 0 -1 2305
box -2 -3 10 103
use NAND3X1  NAND3X1_253
timestamp 1625156677
transform -1 0 3988 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_279
timestamp 1625156677
transform -1 0 4012 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_251
timestamp 1625156677
transform 1 0 4012 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_241
timestamp 1625156677
transform -1 0 4076 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_240
timestamp 1625156677
transform 1 0 4076 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_154
timestamp 1625156677
transform 1 0 4108 0 -1 2305
box -2 -3 26 103
use AND2X2  AND2X2_85
timestamp 1625156677
transform -1 0 4164 0 -1 2305
box -2 -3 34 103
use XOR2X1  XOR2X1_120
timestamp 1625156677
transform 1 0 4164 0 -1 2305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_106
timestamp 1625156677
transform 1 0 4220 0 -1 2305
box -2 -3 58 103
use NAND3X1  NAND3X1_219
timestamp 1625156677
transform -1 0 4308 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_233
timestamp 1625156677
transform -1 0 4332 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_206
timestamp 1625156677
transform 1 0 4332 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_207
timestamp 1625156677
transform 1 0 4364 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_199
timestamp 1625156677
transform -1 0 4428 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_8_0
timestamp 1625156677
transform -1 0 4436 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_8_1
timestamp 1625156677
transform -1 0 4444 0 -1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_196
timestamp 1625156677
transform -1 0 4476 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_198
timestamp 1625156677
transform 1 0 4476 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_234
timestamp 1625156677
transform -1 0 4532 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_133
timestamp 1625156677
transform 1 0 4532 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_140
timestamp 1625156677
transform 1 0 4556 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_204
timestamp 1625156677
transform 1 0 4572 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_147
timestamp 1625156677
transform 1 0 4604 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_131
timestamp 1625156677
transform 1 0 4636 0 -1 2305
box -2 -3 26 103
use INVX2  INVX2_45
timestamp 1625156677
transform 1 0 4660 0 -1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_152
timestamp 1625156677
transform 1 0 4676 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_154
timestamp 1625156677
transform 1 0 4708 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_237
timestamp 1625156677
transform 1 0 4740 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_218
timestamp 1625156677
transform 1 0 4764 0 -1 2305
box -2 -3 34 103
use XOR2X1  XOR2X1_126
timestamp 1625156677
transform -1 0 4852 0 -1 2305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_107
timestamp 1625156677
transform 1 0 4852 0 -1 2305
box -2 -3 58 103
use OAI21X1  OAI21X1_208
timestamp 1625156677
transform 1 0 4908 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_246
timestamp 1625156677
transform -1 0 4964 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_9_0
timestamp 1625156677
transform 1 0 4964 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_9_1
timestamp 1625156677
transform 1 0 4972 0 -1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_205
timestamp 1625156677
transform 1 0 4980 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_149
timestamp 1625156677
transform -1 0 5044 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_240
timestamp 1625156677
transform 1 0 5044 0 -1 2305
box -2 -3 26 103
use INVX2  INVX2_46
timestamp 1625156677
transform 1 0 5068 0 -1 2305
box -2 -3 18 103
use XOR2X1  XOR2X1_106
timestamp 1625156677
transform 1 0 5084 0 -1 2305
box -2 -3 58 103
use OR2X2  OR2X2_92
timestamp 1625156677
transform 1 0 5140 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_148
timestamp 1625156677
transform 1 0 5172 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_132
timestamp 1625156677
transform 1 0 5204 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_236
timestamp 1625156677
transform -1 0 5252 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_221
timestamp 1625156677
transform -1 0 5276 0 -1 2305
box -2 -3 26 103
use AND2X2  AND2X2_71
timestamp 1625156677
transform 1 0 5276 0 -1 2305
box -2 -3 34 103
use FILL  FILL_23_1
timestamp 1625156677
transform -1 0 5316 0 -1 2305
box -2 -3 10 103
use BUFX2  BUFX2_109
timestamp 1625156677
transform 1 0 4 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_219
timestamp 1625156677
transform 1 0 28 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_387
timestamp 1625156677
transform 1 0 52 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_386
timestamp 1625156677
transform -1 0 100 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_229
timestamp 1625156677
transform 1 0 100 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_335
timestamp 1625156677
transform 1 0 132 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_249
timestamp 1625156677
transform -1 0 180 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_347
timestamp 1625156677
transform -1 0 212 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_256
timestamp 1625156677
transform 1 0 212 0 1 2105
box -2 -3 18 103
use NOR3X1  NOR3X1_63
timestamp 1625156677
transform -1 0 292 0 1 2105
box -2 -3 66 103
use XNOR2X1  XNOR2X1_160
timestamp 1625156677
transform -1 0 348 0 1 2105
box -2 -3 58 103
use FILL  FILL_21_0_0
timestamp 1625156677
transform -1 0 356 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_0_1
timestamp 1625156677
transform -1 0 364 0 1 2105
box -2 -3 10 103
use NOR2X1  NOR2X1_218
timestamp 1625156677
transform -1 0 388 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_341
timestamp 1625156677
transform -1 0 420 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_385
timestamp 1625156677
transform -1 0 444 0 1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_333
timestamp 1625156677
transform 1 0 444 0 1 2105
box -2 -3 34 103
use INVX2  INVX2_62
timestamp 1625156677
transform 1 0 476 0 1 2105
box -2 -3 18 103
use NOR3X1  NOR3X1_64
timestamp 1625156677
transform -1 0 556 0 1 2105
box -2 -3 66 103
use OAI21X1  OAI21X1_339
timestamp 1625156677
transform 1 0 556 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_342
timestamp 1625156677
transform 1 0 588 0 1 2105
box -2 -3 34 103
use AND2X2  AND2X2_111
timestamp 1625156677
transform -1 0 652 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_332
timestamp 1625156677
transform 1 0 652 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_383
timestamp 1625156677
transform 1 0 684 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_215
timestamp 1625156677
transform 1 0 708 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_338
timestamp 1625156677
transform 1 0 732 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_245
timestamp 1625156677
transform -1 0 780 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_249
timestamp 1625156677
transform -1 0 804 0 1 2105
box -2 -3 26 103
use AND2X2  AND2X2_110
timestamp 1625156677
transform -1 0 836 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_214
timestamp 1625156677
transform 1 0 836 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_1_0
timestamp 1625156677
transform -1 0 868 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_1_1
timestamp 1625156677
transform -1 0 876 0 1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_381
timestamp 1625156677
transform -1 0 900 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_337
timestamp 1625156677
transform 1 0 900 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_244
timestamp 1625156677
transform -1 0 948 0 1 2105
box -2 -3 18 103
use BUFX2  BUFX2_202
timestamp 1625156677
transform 1 0 948 0 1 2105
box -2 -3 26 103
use BUFX2  BUFX2_201
timestamp 1625156677
transform -1 0 996 0 1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_268
timestamp 1625156677
transform -1 0 1092 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_277
timestamp 1625156677
transform -1 0 1188 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_275
timestamp 1625156677
transform -1 0 1284 0 1 2105
box -2 -3 98 103
use INVX1  INVX1_538
timestamp 1625156677
transform -1 0 1300 0 1 2105
box -2 -3 18 103
use BUFX2  BUFX2_55
timestamp 1625156677
transform -1 0 1324 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_2_0
timestamp 1625156677
transform -1 0 1332 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_2_1
timestamp 1625156677
transform -1 0 1340 0 1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_267
timestamp 1625156677
transform -1 0 1436 0 1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_293
timestamp 1625156677
transform -1 0 1532 0 1 2105
box -2 -3 98 103
use OAI21X1  OAI21X1_624
timestamp 1625156677
transform 1 0 1532 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_567
timestamp 1625156677
transform -1 0 1580 0 1 2105
box -2 -3 18 103
use OR2X2  OR2X2_143
timestamp 1625156677
transform 1 0 1580 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_387
timestamp 1625156677
transform 1 0 1612 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_511
timestamp 1625156677
transform 1 0 1644 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_658
timestamp 1625156677
transform 1 0 1676 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_627
timestamp 1625156677
transform -1 0 1732 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_432
timestamp 1625156677
transform -1 0 1756 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_571
timestamp 1625156677
transform 1 0 1756 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_243
timestamp 1625156677
transform -1 0 1868 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_3_0
timestamp 1625156677
transform -1 0 1876 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_3_1
timestamp 1625156677
transform -1 0 1884 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_628
timestamp 1625156677
transform -1 0 1916 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_392
timestamp 1625156677
transform -1 0 1948 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_512
timestamp 1625156677
transform 1 0 1948 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_365
timestamp 1625156677
transform 1 0 1980 0 1 2105
box -2 -3 98 103
use INVX1  INVX1_566
timestamp 1625156677
transform -1 0 2092 0 1 2105
box -2 -3 18 103
use INVX1  INVX1_574
timestamp 1625156677
transform 1 0 2092 0 1 2105
box -2 -3 18 103
use NAND3X1  NAND3X1_514
timestamp 1625156677
transform 1 0 2108 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_544
timestamp 1625156677
transform 1 0 2140 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_616
timestamp 1625156677
transform -1 0 2188 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_418
timestamp 1625156677
transform -1 0 2212 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_643
timestamp 1625156677
transform -1 0 2236 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_502
timestamp 1625156677
transform -1 0 2252 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_419
timestamp 1625156677
transform 1 0 2252 0 1 2105
box -2 -3 26 103
use INVX2  INVX2_85
timestamp 1625156677
transform 1 0 2276 0 1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_244
timestamp 1625156677
transform -1 0 2388 0 1 2105
box -2 -3 98 103
use FILL  FILL_21_4_0
timestamp 1625156677
transform -1 0 2396 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_4_1
timestamp 1625156677
transform -1 0 2404 0 1 2105
box -2 -3 10 103
use INVX1  INVX1_530
timestamp 1625156677
transform -1 0 2420 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_597
timestamp 1625156677
transform 1 0 2420 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_358
timestamp 1625156677
transform 1 0 2452 0 1 2105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_212
timestamp 1625156677
transform 1 0 2484 0 1 2105
box -2 -3 58 103
use AND2X2  AND2X2_94
timestamp 1625156677
transform -1 0 2572 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_311
timestamp 1625156677
transform -1 0 2596 0 1 2105
box -2 -3 26 103
use XOR2X1  XOR2X1_145
timestamp 1625156677
transform -1 0 2652 0 1 2105
box -2 -3 58 103
use BUFX2  BUFX2_97
timestamp 1625156677
transform -1 0 2676 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_312
timestamp 1625156677
transform 1 0 2676 0 1 2105
box -2 -3 26 103
use OR2X2  OR2X2_124
timestamp 1625156677
transform -1 0 2732 0 1 2105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_208
timestamp 1625156677
transform 1 0 2732 0 1 2105
box -2 -3 58 103
use AND2X2  AND2X2_95
timestamp 1625156677
transform -1 0 2820 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_379
timestamp 1625156677
transform -1 0 2852 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_503
timestamp 1625156677
transform 1 0 2852 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_650
timestamp 1625156677
transform 1 0 2884 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_5_0
timestamp 1625156677
transform 1 0 2908 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_5_1
timestamp 1625156677
transform 1 0 2916 0 1 2105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_219
timestamp 1625156677
transform 1 0 2924 0 1 2105
box -2 -3 58 103
use XOR2X1  XOR2X1_64
timestamp 1625156677
transform 1 0 2980 0 1 2105
box -2 -3 58 103
use NAND2X1  NAND2X1_159
timestamp 1625156677
transform 1 0 3036 0 1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_136
timestamp 1625156677
transform 1 0 3060 0 1 2105
box -2 -3 34 103
use OR2X2  OR2X2_59
timestamp 1625156677
transform 1 0 3092 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_137
timestamp 1625156677
transform -1 0 3156 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_98
timestamp 1625156677
transform 1 0 3156 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_90
timestamp 1625156677
transform 1 0 3188 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_133
timestamp 1625156677
transform -1 0 3236 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_132
timestamp 1625156677
transform -1 0 3268 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_90
timestamp 1625156677
transform -1 0 3292 0 1 2105
box -2 -3 26 103
use AND2X2  AND2X2_46
timestamp 1625156677
transform -1 0 3324 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_106
timestamp 1625156677
transform 1 0 3324 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_146
timestamp 1625156677
transform -1 0 3388 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_161
timestamp 1625156677
transform 1 0 3388 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_6_0
timestamp 1625156677
transform -1 0 3420 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_6_1
timestamp 1625156677
transform -1 0 3428 0 1 2105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_122
timestamp 1625156677
transform -1 0 3484 0 1 2105
box -2 -3 58 103
use XOR2X1  XOR2X1_62
timestamp 1625156677
transform 1 0 3484 0 1 2105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_67
timestamp 1625156677
transform -1 0 3596 0 1 2105
box -2 -3 58 103
use BUFX2  BUFX2_174
timestamp 1625156677
transform 1 0 3596 0 1 2105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_68
timestamp 1625156677
transform -1 0 3676 0 1 2105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_121
timestamp 1625156677
transform 1 0 3676 0 1 2105
box -2 -3 58 103
use CLKBUF1  CLKBUF1_10
timestamp 1625156677
transform -1 0 3804 0 1 2105
box -2 -3 74 103
use NOR2X1  NOR2X1_156
timestamp 1625156677
transform -1 0 3828 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_157
timestamp 1625156677
transform -1 0 3852 0 1 2105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_126
timestamp 1625156677
transform 1 0 3852 0 1 2105
box -2 -3 58 103
use OAI21X1  OAI21X1_243
timestamp 1625156677
transform 1 0 3908 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_7_0
timestamp 1625156677
transform 1 0 3940 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_7_1
timestamp 1625156677
transform 1 0 3948 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_244
timestamp 1625156677
transform 1 0 3956 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_175
timestamp 1625156677
transform 1 0 3988 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_161
timestamp 1625156677
transform -1 0 4036 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_283
timestamp 1625156677
transform -1 0 4060 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_282
timestamp 1625156677
transform 1 0 4060 0 1 2105
box -2 -3 26 103
use OR2X2  OR2X2_112
timestamp 1625156677
transform 1 0 4084 0 1 2105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_231
timestamp 1625156677
transform 1 0 4116 0 1 2105
box -2 -3 98 103
use INVX1  INVX1_158
timestamp 1625156677
transform 1 0 4212 0 1 2105
box -2 -3 18 103
use NAND3X1  NAND3X1_252
timestamp 1625156677
transform 1 0 4228 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_250
timestamp 1625156677
transform 1 0 4260 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_277
timestamp 1625156677
transform -1 0 4316 0 1 2105
box -2 -3 26 103
use OR2X2  OR2X2_109
timestamp 1625156677
transform -1 0 4348 0 1 2105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_104
timestamp 1625156677
transform 1 0 4348 0 1 2105
box -2 -3 58 103
use AOI21X1  AOI21X1_153
timestamp 1625156677
transform 1 0 4404 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_8_0
timestamp 1625156677
transform -1 0 4444 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_8_1
timestamp 1625156677
transform -1 0 4452 0 1 2105
box -2 -3 10 103
use INVX2  INVX2_44
timestamp 1625156677
transform -1 0 4468 0 1 2105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_105
timestamp 1625156677
transform 1 0 4468 0 1 2105
box -2 -3 58 103
use NAND2X1  NAND2X1_229
timestamp 1625156677
transform 1 0 4524 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_231
timestamp 1625156677
transform -1 0 4572 0 1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_204
timestamp 1625156677
transform -1 0 4604 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_203
timestamp 1625156677
transform 1 0 4604 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_230
timestamp 1625156677
transform 1 0 4636 0 1 2105
box -2 -3 26 103
use OR2X2  OR2X2_89
timestamp 1625156677
transform -1 0 4692 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_132
timestamp 1625156677
transform 1 0 4692 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_195
timestamp 1625156677
transform -1 0 4740 0 1 2105
box -2 -3 34 103
use NOR3X1  NOR3X1_47
timestamp 1625156677
transform 1 0 4740 0 1 2105
box -2 -3 66 103
use NOR2X1  NOR2X1_128
timestamp 1625156677
transform 1 0 4804 0 1 2105
box -2 -3 26 103
use AND2X2  AND2X2_68
timestamp 1625156677
transform -1 0 4860 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_151
timestamp 1625156677
transform 1 0 4860 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_139
timestamp 1625156677
transform 1 0 4892 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_136
timestamp 1625156677
transform 1 0 4908 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_210
timestamp 1625156677
transform -1 0 4964 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_9_0
timestamp 1625156677
transform -1 0 4972 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_9_1
timestamp 1625156677
transform -1 0 4980 0 1 2105
box -2 -3 10 103
use NAND3X1  NAND3X1_220
timestamp 1625156677
transform -1 0 5012 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_245
timestamp 1625156677
transform -1 0 5036 0 1 2105
box -2 -3 26 103
use OR2X2  OR2X2_96
timestamp 1625156677
transform -1 0 5068 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_244
timestamp 1625156677
transform -1 0 5092 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_209
timestamp 1625156677
transform 1 0 5092 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_137
timestamp 1625156677
transform 1 0 5124 0 1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_135
timestamp 1625156677
transform -1 0 5164 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_150
timestamp 1625156677
transform -1 0 5196 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_217
timestamp 1625156677
transform 1 0 5196 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_241
timestamp 1625156677
transform -1 0 5252 0 1 2105
box -2 -3 26 103
use OR2X2  OR2X2_94
timestamp 1625156677
transform 1 0 5252 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_186
timestamp 1625156677
transform -1 0 5316 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_344
timestamp 1625156677
transform 1 0 4 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_343
timestamp 1625156677
transform 1 0 36 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_248
timestamp 1625156677
transform -1 0 84 0 -1 2105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_161
timestamp 1625156677
transform -1 0 140 0 -1 2105
box -2 -3 58 103
use NAND3X1  NAND3X1_334
timestamp 1625156677
transform -1 0 172 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_221
timestamp 1625156677
transform -1 0 196 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_354
timestamp 1625156677
transform 1 0 196 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_388
timestamp 1625156677
transform -1 0 252 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_231
timestamp 1625156677
transform -1 0 284 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_341
timestamp 1625156677
transform 1 0 284 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_247
timestamp 1625156677
transform 1 0 316 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_217
timestamp 1625156677
transform -1 0 356 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_0_0
timestamp 1625156677
transform 1 0 356 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1625156677
transform 1 0 364 0 -1 2105
box -2 -3 10 103
use NOR2X1  NOR2X1_216
timestamp 1625156677
transform 1 0 372 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_384
timestamp 1625156677
transform -1 0 420 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_392
timestamp 1625156677
transform -1 0 444 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_230
timestamp 1625156677
transform 1 0 444 0 -1 2105
box -2 -3 34 103
use AND2X2  AND2X2_113
timestamp 1625156677
transform -1 0 508 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_351
timestamp 1625156677
transform -1 0 540 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_340
timestamp 1625156677
transform 1 0 540 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_246
timestamp 1625156677
transform -1 0 588 0 -1 2105
box -2 -3 18 103
use XOR2X1  XOR2X1_205
timestamp 1625156677
transform -1 0 644 0 -1 2105
box -2 -3 58 103
use BUFX2  BUFX2_187
timestamp 1625156677
transform 1 0 644 0 -1 2105
box -2 -3 26 103
use BUFX2  BUFX2_188
timestamp 1625156677
transform -1 0 692 0 -1 2105
box -2 -3 26 103
use XOR2X1  XOR2X1_181
timestamp 1625156677
transform 1 0 692 0 -1 2105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_170
timestamp 1625156677
transform 1 0 748 0 -1 2105
box -2 -3 58 103
use XOR2X1  XOR2X1_180
timestamp 1625156677
transform 1 0 804 0 -1 2105
box -2 -3 58 103
use FILL  FILL_20_1_0
timestamp 1625156677
transform -1 0 868 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1625156677
transform -1 0 876 0 -1 2105
box -2 -3 10 103
use XOR2X1  XOR2X1_162
timestamp 1625156677
transform -1 0 932 0 -1 2105
box -2 -3 58 103
use AND2X2  AND2X2_102
timestamp 1625156677
transform -1 0 964 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_190
timestamp 1625156677
transform -1 0 988 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_343
timestamp 1625156677
transform -1 0 1012 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_344
timestamp 1625156677
transform -1 0 1036 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_299
timestamp 1625156677
transform 1 0 1036 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_206
timestamp 1625156677
transform -1 0 1084 0 -1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_305
timestamp 1625156677
transform -1 0 1180 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_258
timestamp 1625156677
transform -1 0 1276 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_276
timestamp 1625156677
transform -1 0 1372 0 -1 2105
box -2 -3 98 103
use FILL  FILL_20_2_0
timestamp 1625156677
transform 1 0 1372 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1625156677
transform 1 0 1380 0 -1 2105
box -2 -3 10 103
use XOR2X1  XOR2X1_299
timestamp 1625156677
transform 1 0 1388 0 -1 2105
box -2 -3 58 103
use AND2X2  AND2X2_183
timestamp 1625156677
transform 1 0 1444 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_411
timestamp 1625156677
transform -1 0 1500 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_615
timestamp 1625156677
transform -1 0 1532 0 -1 2105
box -2 -3 34 103
use AND2X2  AND2X2_179
timestamp 1625156677
transform -1 0 1564 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_417
timestamp 1625156677
transform -1 0 1588 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_328
timestamp 1625156677
transform -1 0 1684 0 -1 2105
box -2 -3 98 103
use AOI21X1  AOI21X1_391
timestamp 1625156677
transform 1 0 1684 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_510
timestamp 1625156677
transform -1 0 1732 0 -1 2105
box -2 -3 18 103
use INVX1  INVX1_497
timestamp 1625156677
transform -1 0 1748 0 -1 2105
box -2 -3 18 103
use INVX1  INVX1_176
timestamp 1625156677
transform -1 0 1764 0 -1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_306
timestamp 1625156677
transform 1 0 1764 0 -1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_275
timestamp 1625156677
transform 1 0 1788 0 -1 2105
box -2 -3 34 103
use OR2X2  OR2X2_121
timestamp 1625156677
transform -1 0 1852 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_659
timestamp 1625156677
transform -1 0 1876 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_3_0
timestamp 1625156677
transform -1 0 1884 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1625156677
transform -1 0 1892 0 -1 2105
box -2 -3 10 103
use NOR2X1  NOR2X1_433
timestamp 1625156677
transform -1 0 1916 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_513
timestamp 1625156677
transform -1 0 1932 0 -1 2105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_228
timestamp 1625156677
transform 1 0 1932 0 -1 2105
box -2 -3 58 103
use AOI21X1  AOI21X1_371
timestamp 1625156677
transform -1 0 2020 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_641
timestamp 1625156677
transform -1 0 2044 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_642
timestamp 1625156677
transform 1 0 2044 0 -1 2105
box -2 -3 26 103
use OR2X2  OR2X2_132
timestamp 1625156677
transform -1 0 2100 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_690
timestamp 1625156677
transform -1 0 2124 0 -1 2105
box -2 -3 26 103
use XOR2X1  XOR2X1_143
timestamp 1625156677
transform -1 0 2180 0 -1 2105
box -2 -3 58 103
use NAND2X1  NAND2X1_693
timestamp 1625156677
transform -1 0 2204 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_245
timestamp 1625156677
transform 1 0 2204 0 -1 2105
box -2 -3 98 103
use INVX1  INVX1_177
timestamp 1625156677
transform 1 0 2300 0 -1 2105
box -2 -3 18 103
use INVX1  INVX1_178
timestamp 1625156677
transform 1 0 2316 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_269
timestamp 1625156677
transform -1 0 2364 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_268
timestamp 1625156677
transform 1 0 2364 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_4_0
timestamp 1625156677
transform 1 0 2396 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_4_1
timestamp 1625156677
transform 1 0 2404 0 -1 2105
box -2 -3 10 103
use NAND3X1  NAND3X1_281
timestamp 1625156677
transform 1 0 2412 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_280
timestamp 1625156677
transform 1 0 2444 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_194
timestamp 1625156677
transform -1 0 2508 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_285
timestamp 1625156677
transform -1 0 2540 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_170
timestamp 1625156677
transform 1 0 2540 0 -1 2105
box -2 -3 26 103
use OR2X2  OR2X2_123
timestamp 1625156677
transform -1 0 2596 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_283
timestamp 1625156677
transform 1 0 2596 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_196
timestamp 1625156677
transform -1 0 2660 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_284
timestamp 1625156677
transform 1 0 2660 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_282
timestamp 1625156677
transform -1 0 2724 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_179
timestamp 1625156677
transform 1 0 2724 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_271
timestamp 1625156677
transform -1 0 2772 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_270
timestamp 1625156677
transform -1 0 2804 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_172
timestamp 1625156677
transform 1 0 2804 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_661
timestamp 1625156677
transform 1 0 2828 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_662
timestamp 1625156677
transform -1 0 2876 0 -1 2105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_235
timestamp 1625156677
transform -1 0 2932 0 -1 2105
box -2 -3 58 103
use FILL  FILL_20_5_0
timestamp 1625156677
transform -1 0 2940 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_5_1
timestamp 1625156677
transform -1 0 2948 0 -1 2105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_266
timestamp 1625156677
transform -1 0 3044 0 -1 2105
box -2 -3 98 103
use AND2X2  AND2X2_47
timestamp 1625156677
transform -1 0 3076 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_92
timestamp 1625156677
transform -1 0 3100 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_134
timestamp 1625156677
transform 1 0 3100 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_135
timestamp 1625156677
transform 1 0 3132 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_91
timestamp 1625156677
transform -1 0 3180 0 -1 2105
box -2 -3 18 103
use NAND3X1  NAND3X1_138
timestamp 1625156677
transform 1 0 3180 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_140
timestamp 1625156677
transform 1 0 3212 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_139
timestamp 1625156677
transform 1 0 3244 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_143
timestamp 1625156677
transform -1 0 3308 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_141
timestamp 1625156677
transform 1 0 3308 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_164
timestamp 1625156677
transform 1 0 3340 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_101
timestamp 1625156677
transform 1 0 3364 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_140
timestamp 1625156677
transform -1 0 3428 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_6_0
timestamp 1625156677
transform -1 0 3436 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_6_1
timestamp 1625156677
transform -1 0 3444 0 -1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_162
timestamp 1625156677
transform -1 0 3468 0 -1 2105
box -2 -3 26 103
use AND2X2  AND2X2_48
timestamp 1625156677
transform 1 0 3468 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_170
timestamp 1625156677
transform -1 0 3524 0 -1 2105
box -2 -3 26 103
use INVX2  INVX2_34
timestamp 1625156677
transform 1 0 3524 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_137
timestamp 1625156677
transform -1 0 3572 0 -1 2105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_71
timestamp 1625156677
transform -1 0 3628 0 -1 2105
box -2 -3 58 103
use XOR2X1  XOR2X1_146
timestamp 1625156677
transform 1 0 3628 0 -1 2105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_72
timestamp 1625156677
transform -1 0 3740 0 -1 2105
box -2 -3 58 103
use CLKBUF1  CLKBUF1_3
timestamp 1625156677
transform -1 0 3812 0 -1 2105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_211
timestamp 1625156677
transform 1 0 3812 0 -1 2105
box -2 -3 98 103
use FILL  FILL_20_7_0
timestamp 1625156677
transform -1 0 3916 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_7_1
timestamp 1625156677
transform -1 0 3924 0 -1 2105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_36
timestamp 1625156677
transform -1 0 3996 0 -1 2105
box -2 -3 74 103
use XOR2X1  XOR2X1_122
timestamp 1625156677
transform -1 0 4052 0 -1 2105
box -2 -3 58 103
use INVX1  INVX1_163
timestamp 1625156677
transform 1 0 4052 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_245
timestamp 1625156677
transform 1 0 4068 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_256
timestamp 1625156677
transform 1 0 4100 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_164
timestamp 1625156677
transform -1 0 4148 0 -1 2105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_129
timestamp 1625156677
transform 1 0 4148 0 -1 2105
box -2 -3 58 103
use NAND2X1  NAND2X1_281
timestamp 1625156677
transform -1 0 4228 0 -1 2105
box -2 -3 26 103
use OR2X2  OR2X2_111
timestamp 1625156677
transform -1 0 4260 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_280
timestamp 1625156677
transform 1 0 4260 0 -1 2105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1625156677
transform -1 0 4380 0 -1 2105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_210
timestamp 1625156677
transform 1 0 4380 0 -1 2105
box -2 -3 98 103
use FILL  FILL_20_8_0
timestamp 1625156677
transform 1 0 4476 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_8_1
timestamp 1625156677
transform 1 0 4484 0 -1 2105
box -2 -3 10 103
use XOR2X1  XOR2X1_87
timestamp 1625156677
transform 1 0 4492 0 -1 2105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_127
timestamp 1625156677
transform 1 0 4548 0 -1 2105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_103
timestamp 1625156677
transform 1 0 4604 0 -1 2105
box -2 -3 58 103
use XOR2X1  XOR2X1_102
timestamp 1625156677
transform -1 0 4716 0 -1 2105
box -2 -3 58 103
use XOR2X1  XOR2X1_86
timestamp 1625156677
transform 1 0 4716 0 -1 2105
box -2 -3 58 103
use XOR2X1  XOR2X1_127
timestamp 1625156677
transform -1 0 4828 0 -1 2105
box -2 -3 58 103
use XOR2X1  XOR2X1_128
timestamp 1625156677
transform -1 0 4884 0 -1 2105
box -2 -3 58 103
use NOR2X1  NOR2X1_137
timestamp 1625156677
transform 1 0 4884 0 -1 2105
box -2 -3 26 103
use XOR2X1  XOR2X1_103
timestamp 1625156677
transform -1 0 4964 0 -1 2105
box -2 -3 58 103
use FILL  FILL_20_9_0
timestamp 1625156677
transform 1 0 4964 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_9_1
timestamp 1625156677
transform 1 0 4972 0 -1 2105
box -2 -3 10 103
use BUFX2  BUFX2_160
timestamp 1625156677
transform 1 0 4980 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_247
timestamp 1625156677
transform 1 0 5004 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_141
timestamp 1625156677
transform 1 0 5028 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_211
timestamp 1625156677
transform 1 0 5044 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_243
timestamp 1625156677
transform 1 0 5076 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_142
timestamp 1625156677
transform -1 0 5116 0 -1 2105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_111
timestamp 1625156677
transform -1 0 5172 0 -1 2105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_108
timestamp 1625156677
transform -1 0 5228 0 -1 2105
box -2 -3 58 103
use BUFX2  BUFX2_159
timestamp 1625156677
transform 1 0 5228 0 -1 2105
box -2 -3 26 103
use BUFX2  BUFX2_263
timestamp 1625156677
transform 1 0 5252 0 -1 2105
box -2 -3 26 103
use BUFX2  BUFX2_74
timestamp 1625156677
transform 1 0 5276 0 -1 2105
box -2 -3 26 103
use FILL  FILL_21_1
timestamp 1625156677
transform -1 0 5308 0 -1 2105
box -2 -3 10 103
use FILL  FILL_21_2
timestamp 1625156677
transform -1 0 5316 0 -1 2105
box -2 -3 10 103
use INVX1  INVX1_250
timestamp 1625156677
transform -1 0 20 0 1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_338
timestamp 1625156677
transform -1 0 52 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_227
timestamp 1625156677
transform -1 0 84 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_220
timestamp 1625156677
transform 1 0 84 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_348
timestamp 1625156677
transform 1 0 108 0 1 1905
box -2 -3 34 103
use XOR2X1  XOR2X1_197
timestamp 1625156677
transform 1 0 140 0 1 1905
box -2 -3 58 103
use NAND2X1  NAND2X1_393
timestamp 1625156677
transform 1 0 196 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_255
timestamp 1625156677
transform 1 0 220 0 1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_340
timestamp 1625156677
transform -1 0 268 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_232
timestamp 1625156677
transform -1 0 300 0 1 1905
box -2 -3 34 103
use AOI22X1  AOI22X1_11
timestamp 1625156677
transform -1 0 340 0 1 1905
box -2 -3 42 103
use FILL  FILL_19_0_0
timestamp 1625156677
transform -1 0 348 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1625156677
transform -1 0 356 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_350
timestamp 1625156677
transform -1 0 388 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_353
timestamp 1625156677
transform 1 0 388 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_260
timestamp 1625156677
transform -1 0 436 0 1 1905
box -2 -3 18 103
use INVX1  INVX1_261
timestamp 1625156677
transform 1 0 436 0 1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_343
timestamp 1625156677
transform -1 0 484 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_234
timestamp 1625156677
transform 1 0 484 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_397
timestamp 1625156677
transform -1 0 540 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_259
timestamp 1625156677
transform -1 0 556 0 1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_344
timestamp 1625156677
transform 1 0 556 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_262
timestamp 1625156677
transform -1 0 604 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_355
timestamp 1625156677
transform 1 0 604 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_399
timestamp 1625156677
transform -1 0 660 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_279
timestamp 1625156677
transform -1 0 756 0 1 1905
box -2 -3 98 103
use AND2X2  AND2X2_104
timestamp 1625156677
transform -1 0 788 0 1 1905
box -2 -3 34 103
use NOR3X1  NOR3X1_60
timestamp 1625156677
transform -1 0 852 0 1 1905
box -2 -3 66 103
use FILL  FILL_19_1_0
timestamp 1625156677
transform -1 0 860 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1625156677
transform -1 0 868 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_301
timestamp 1625156677
transform -1 0 900 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_304
timestamp 1625156677
transform 1 0 900 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_60
timestamp 1625156677
transform -1 0 948 0 1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_214
timestamp 1625156677
transform -1 0 980 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_306
timestamp 1625156677
transform 1 0 980 0 1 1905
box -2 -3 34 103
use AND2X2  AND2X2_103
timestamp 1625156677
transform -1 0 1044 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_345
timestamp 1625156677
transform -1 0 1068 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_207
timestamp 1625156677
transform -1 0 1084 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_191
timestamp 1625156677
transform 1 0 1084 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_300
timestamp 1625156677
transform -1 0 1140 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_540
timestamp 1625156677
transform -1 0 1156 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_259
timestamp 1625156677
transform -1 0 1252 0 1 1905
box -2 -3 98 103
use INVX1  INVX1_511
timestamp 1625156677
transform -1 0 1268 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_590
timestamp 1625156677
transform 1 0 1268 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_351
timestamp 1625156677
transform 1 0 1300 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_494
timestamp 1625156677
transform -1 0 1348 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_412
timestamp 1625156677
transform -1 0 1372 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_2_0
timestamp 1625156677
transform -1 0 1380 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1625156677
transform -1 0 1388 0 1 1905
box -2 -3 10 103
use XNOR2X1  XNOR2X1_241
timestamp 1625156677
transform -1 0 1444 0 1 1905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_227
timestamp 1625156677
transform 1 0 1444 0 1 1905
box -2 -3 58 103
use AOI21X1  AOI21X1_363
timestamp 1625156677
transform -1 0 1532 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_602
timestamp 1625156677
transform 1 0 1532 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_523
timestamp 1625156677
transform -1 0 1596 0 1 1905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_237
timestamp 1625156677
transform -1 0 1652 0 1 1905
box -2 -3 58 103
use NOR3X1  NOR3X1_55
timestamp 1625156677
transform -1 0 1716 0 1 1905
box -2 -3 66 103
use OAI21X1  OAI21X1_263
timestamp 1625156677
transform 1 0 1716 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_168
timestamp 1625156677
transform 1 0 1748 0 1 1905
box -2 -3 26 103
use AND2X2  AND2X2_92
timestamp 1625156677
transform -1 0 1804 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_508
timestamp 1625156677
transform -1 0 1820 0 1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_276
timestamp 1625156677
transform -1 0 1852 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_307
timestamp 1625156677
transform 1 0 1852 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_3_0
timestamp 1625156677
transform -1 0 1884 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1625156677
transform -1 0 1892 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_603
timestamp 1625156677
transform -1 0 1924 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_364
timestamp 1625156677
transform -1 0 1956 0 1 1905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_139
timestamp 1625156677
transform 1 0 1956 0 1 1905
box -2 -3 58 103
use NAND3X1  NAND3X1_279
timestamp 1625156677
transform -1 0 2044 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_278
timestamp 1625156677
transform -1 0 2076 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_309
timestamp 1625156677
transform 1 0 2076 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_266
timestamp 1625156677
transform -1 0 2132 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_264
timestamp 1625156677
transform -1 0 2164 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_195
timestamp 1625156677
transform 1 0 2164 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_173
timestamp 1625156677
transform 1 0 2196 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_191
timestamp 1625156677
transform 1 0 2220 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_277
timestamp 1625156677
transform -1 0 2284 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_265
timestamp 1625156677
transform 1 0 2284 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_193
timestamp 1625156677
transform -1 0 2348 0 1 1905
box -2 -3 34 103
use NOR3X1  NOR3X1_56
timestamp 1625156677
transform 1 0 2348 0 1 1905
box -2 -3 66 103
use FILL  FILL_19_4_0
timestamp 1625156677
transform -1 0 2420 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_4_1
timestamp 1625156677
transform -1 0 2428 0 1 1905
box -2 -3 10 103
use AOI21X1  AOI21X1_192
timestamp 1625156677
transform -1 0 2460 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_169
timestamp 1625156677
transform -1 0 2484 0 1 1905
box -2 -3 26 103
use XOR2X1  XOR2X1_142
timestamp 1625156677
transform -1 0 2540 0 1 1905
box -2 -3 58 103
use BUFX2  BUFX2_172
timestamp 1625156677
transform -1 0 2564 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_315
timestamp 1625156677
transform 1 0 2564 0 1 1905
box -2 -3 26 103
use XOR2X1  XOR2X1_144
timestamp 1625156677
transform -1 0 2644 0 1 1905
box -2 -3 58 103
use INVX2  INVX2_56
timestamp 1625156677
transform -1 0 2660 0 1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_242
timestamp 1625156677
transform -1 0 2756 0 1 1905
box -2 -3 98 103
use BUFX2  BUFX2_173
timestamp 1625156677
transform 1 0 2756 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_614
timestamp 1625156677
transform -1 0 2812 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_416
timestamp 1625156677
transform -1 0 2836 0 1 1905
box -2 -3 26 103
use AND2X2  AND2X2_178
timestamp 1625156677
transform -1 0 2868 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_557
timestamp 1625156677
transform -1 0 2884 0 1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_640
timestamp 1625156677
transform -1 0 2908 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_5_0
timestamp 1625156677
transform -1 0 2916 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_5_1
timestamp 1625156677
transform -1 0 2924 0 1 1905
box -2 -3 10 103
use INVX1  INVX1_501
timestamp 1625156677
transform -1 0 2940 0 1 1905
box -2 -3 18 103
use XOR2X1  XOR2X1_147
timestamp 1625156677
transform -1 0 2996 0 1 1905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_226
timestamp 1625156677
transform 1 0 2996 0 1 1905
box -2 -3 98 103
use OR2X2  OR2X2_60
timestamp 1625156677
transform 1 0 3092 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_145
timestamp 1625156677
transform 1 0 3124 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_100
timestamp 1625156677
transform 1 0 3156 0 1 1905
box -2 -3 34 103
use OR2X2  OR2X2_62
timestamp 1625156677
transform 1 0 3188 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_102
timestamp 1625156677
transform 1 0 3220 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_95
timestamp 1625156677
transform 1 0 3252 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_93
timestamp 1625156677
transform -1 0 3292 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_141
timestamp 1625156677
transform -1 0 3324 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_142
timestamp 1625156677
transform 1 0 3324 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_50
timestamp 1625156677
transform 1 0 3356 0 1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_103
timestamp 1625156677
transform 1 0 3372 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_95
timestamp 1625156677
transform 1 0 3404 0 1 1905
box -2 -3 18 103
use FILL  FILL_19_6_0
timestamp 1625156677
transform 1 0 3420 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_6_1
timestamp 1625156677
transform 1 0 3428 0 1 1905
box -2 -3 10 103
use NOR2X1  NOR2X1_96
timestamp 1625156677
transform 1 0 3436 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_97
timestamp 1625156677
transform -1 0 3484 0 1 1905
box -2 -3 26 103
use XOR2X1  XOR2X1_101
timestamp 1625156677
transform -1 0 3540 0 1 1905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_92
timestamp 1625156677
transform -1 0 3596 0 1 1905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_218
timestamp 1625156677
transform 1 0 3596 0 1 1905
box -2 -3 98 103
use XOR2X1  XOR2X1_88
timestamp 1625156677
transform 1 0 3692 0 1 1905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1625156677
transform -1 0 3844 0 1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_200
timestamp 1625156677
transform 1 0 3844 0 1 1905
box -2 -3 98 103
use FILL  FILL_19_7_0
timestamp 1625156677
transform 1 0 3940 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_7_1
timestamp 1625156677
transform 1 0 3948 0 1 1905
box -2 -3 10 103
use INVX1  INVX1_116
timestamp 1625156677
transform 1 0 3956 0 1 1905
box -2 -3 18 103
use XNOR2X1  XNOR2X1_91
timestamp 1625156677
transform -1 0 4028 0 1 1905
box -2 -3 58 103
use NAND2X1  NAND2X1_204
timestamp 1625156677
transform 1 0 4028 0 1 1905
box -2 -3 26 103
use OR2X2  OR2X2_79
timestamp 1625156677
transform 1 0 4052 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_285
timestamp 1625156677
transform -1 0 4108 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_205
timestamp 1625156677
transform 1 0 4108 0 1 1905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_93
timestamp 1625156677
transform -1 0 4188 0 1 1905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_128
timestamp 1625156677
transform 1 0 4188 0 1 1905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_220
timestamp 1625156677
transform 1 0 4244 0 1 1905
box -2 -3 98 103
use INVX1  INVX1_144
timestamp 1625156677
transform 1 0 4340 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_214
timestamp 1625156677
transform -1 0 4388 0 1 1905
box -2 -3 34 103
use NOR3X1  NOR3X1_50
timestamp 1625156677
transform 1 0 4388 0 1 1905
box -2 -3 66 103
use FILL  FILL_19_8_0
timestamp 1625156677
transform 1 0 4452 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_8_1
timestamp 1625156677
transform 1 0 4460 0 1 1905
box -2 -3 10 103
use NOR2X1  NOR2X1_139
timestamp 1625156677
transform 1 0 4468 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_251
timestamp 1625156677
transform -1 0 4516 0 1 1905
box -2 -3 26 103
use AND2X2  AND2X2_75
timestamp 1625156677
transform -1 0 4548 0 1 1905
box -2 -3 34 103
use XOR2X1  XOR2X1_114
timestamp 1625156677
transform -1 0 4604 0 1 1905
box -2 -3 58 103
use AND2X2  AND2X2_76
timestamp 1625156677
transform -1 0 4636 0 1 1905
box -2 -3 34 103
use XOR2X1  XOR2X1_113
timestamp 1625156677
transform -1 0 4692 0 1 1905
box -2 -3 58 103
use XOR2X1  XOR2X1_115
timestamp 1625156677
transform -1 0 4748 0 1 1905
box -2 -3 58 103
use XOR2X1  XOR2X1_129
timestamp 1625156677
transform -1 0 4804 0 1 1905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_109
timestamp 1625156677
transform 1 0 4804 0 1 1905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_213
timestamp 1625156677
transform 1 0 4860 0 1 1905
box -2 -3 98 103
use FILL  FILL_19_9_0
timestamp 1625156677
transform -1 0 4964 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_9_1
timestamp 1625156677
transform -1 0 4972 0 1 1905
box -2 -3 10 103
use XNOR2X1  XNOR2X1_110
timestamp 1625156677
transform -1 0 5028 0 1 1905
box -2 -3 58 103
use NAND2X1  NAND2X1_242
timestamp 1625156677
transform 1 0 5028 0 1 1905
box -2 -3 26 103
use OR2X2  OR2X2_95
timestamp 1625156677
transform 1 0 5052 0 1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_215
timestamp 1625156677
transform 1 0 5084 0 1 1905
box -2 -3 98 103
use BUFX2  BUFX2_272
timestamp 1625156677
transform -1 0 5204 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_217
timestamp 1625156677
transform -1 0 5228 0 1 1905
box -2 -3 26 103
use AND2X2  AND2X2_65
timestamp 1625156677
transform 1 0 5228 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_197
timestamp 1625156677
transform -1 0 5292 0 1 1905
box -2 -3 34 103
use FILL  FILL_20_1
timestamp 1625156677
transform 1 0 5292 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_2
timestamp 1625156677
transform 1 0 5300 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_3
timestamp 1625156677
transform 1 0 5308 0 1 1905
box -2 -3 10 103
use XOR2X1  XOR2X1_183
timestamp 1625156677
transform -1 0 60 0 -1 1905
box -2 -3 58 103
use AOI21X1  AOI21X1_228
timestamp 1625156677
transform -1 0 92 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_342
timestamp 1625156677
transform -1 0 124 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_398
timestamp 1625156677
transform 1 0 124 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_233
timestamp 1625156677
transform -1 0 180 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_391
timestamp 1625156677
transform 1 0 180 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_339
timestamp 1625156677
transform 1 0 204 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_349
timestamp 1625156677
transform 1 0 236 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_389
timestamp 1625156677
transform -1 0 292 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_254
timestamp 1625156677
transform -1 0 308 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_390
timestamp 1625156677
transform 1 0 308 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_222
timestamp 1625156677
transform 1 0 332 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_0_0
timestamp 1625156677
transform 1 0 356 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1625156677
transform 1 0 364 0 -1 1905
box -2 -3 10 103
use INVX1  INVX1_257
timestamp 1625156677
transform 1 0 372 0 -1 1905
box -2 -3 18 103
use XOR2X1  XOR2X1_182
timestamp 1625156677
transform -1 0 444 0 -1 1905
box -2 -3 58 103
use NAND2X1  NAND2X1_414
timestamp 1625156677
transform 1 0 444 0 -1 1905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_167
timestamp 1625156677
transform -1 0 524 0 -1 1905
box -2 -3 58 103
use NAND2X1  NAND2X1_396
timestamp 1625156677
transform 1 0 524 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_224
timestamp 1625156677
transform -1 0 572 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_278
timestamp 1625156677
transform -1 0 668 0 -1 1905
box -2 -3 98 103
use XNOR2X1  XNOR2X1_152
timestamp 1625156677
transform 1 0 668 0 -1 1905
box -2 -3 58 103
use NAND2X1  NAND2X1_350
timestamp 1625156677
transform -1 0 748 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_218
timestamp 1625156677
transform 1 0 748 0 -1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_215
timestamp 1625156677
transform -1 0 796 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_315
timestamp 1625156677
transform -1 0 828 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_209
timestamp 1625156677
transform -1 0 844 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_193
timestamp 1625156677
transform -1 0 868 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_1_0
timestamp 1625156677
transform -1 0 876 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1625156677
transform -1 0 884 0 -1 1905
box -2 -3 10 103
use NAND2X1  NAND2X1_347
timestamp 1625156677
transform -1 0 908 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_307
timestamp 1625156677
transform 1 0 908 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_346
timestamp 1625156677
transform -1 0 964 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_354
timestamp 1625156677
transform -1 0 988 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_192
timestamp 1625156677
transform 1 0 988 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_313
timestamp 1625156677
transform -1 0 1044 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_208
timestamp 1625156677
transform -1 0 1060 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_302
timestamp 1625156677
transform -1 0 1092 0 -1 1905
box -2 -3 34 103
use XOR2X1  XOR2X1_164
timestamp 1625156677
transform -1 0 1148 0 -1 1905
box -2 -3 58 103
use XOR2X1  XOR2X1_163
timestamp 1625156677
transform 1 0 1148 0 -1 1905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_274
timestamp 1625156677
transform -1 0 1300 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_539
timestamp 1625156677
transform -1 0 1316 0 -1 1905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_260
timestamp 1625156677
transform -1 0 1412 0 -1 1905
box -2 -3 98 103
use FILL  FILL_18_2_0
timestamp 1625156677
transform -1 0 1420 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1625156677
transform -1 0 1428 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_304
timestamp 1625156677
transform -1 0 1524 0 -1 1905
box -2 -3 98 103
use XOR2X1  XOR2X1_301
timestamp 1625156677
transform 1 0 1524 0 -1 1905
box -2 -3 58 103
use NOR2X1  NOR2X1_413
timestamp 1625156677
transform 1 0 1580 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_514
timestamp 1625156677
transform -1 0 1620 0 -1 1905
box -2 -3 18 103
use AND2X2  AND2X2_184
timestamp 1625156677
transform 1 0 1620 0 -1 1905
box -2 -3 34 103
use BUFX2  BUFX2_107
timestamp 1625156677
transform -1 0 1676 0 -1 1905
box -2 -3 26 103
use AND2X2  AND2X2_185
timestamp 1625156677
transform 1 0 1676 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_382
timestamp 1625156677
transform -1 0 1740 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_666
timestamp 1625156677
transform 1 0 1740 0 -1 1905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_140
timestamp 1625156677
transform 1 0 1764 0 -1 1905
box -2 -3 58 103
use NAND2X1  NAND2X1_305
timestamp 1625156677
transform 1 0 1820 0 -1 1905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_141
timestamp 1625156677
transform -1 0 1900 0 -1 1905
box -2 -3 58 103
use FILL  FILL_18_3_0
timestamp 1625156677
transform -1 0 1908 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1625156677
transform -1 0 1916 0 -1 1905
box -2 -3 10 103
use AOI21X1  AOI21X1_201
timestamp 1625156677
transform -1 0 1948 0 -1 1905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_142
timestamp 1625156677
transform -1 0 2004 0 -1 1905
box -2 -3 58 103
use NAND3X1  NAND3X1_291
timestamp 1625156677
transform 1 0 2004 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_267
timestamp 1625156677
transform -1 0 2068 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_310
timestamp 1625156677
transform 1 0 2068 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_184
timestamp 1625156677
transform 1 0 2092 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_272
timestamp 1625156677
transform 1 0 2108 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_200
timestamp 1625156677
transform 1 0 2140 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_429
timestamp 1625156677
transform -1 0 2196 0 -1 1905
box -2 -3 26 103
use OR2X2  OR2X2_122
timestamp 1625156677
transform 1 0 2196 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_308
timestamp 1625156677
transform -1 0 2252 0 -1 1905
box -2 -3 26 103
use AND2X2  AND2X2_93
timestamp 1625156677
transform 1 0 2252 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_689
timestamp 1625156677
transform 1 0 2284 0 -1 1905
box -2 -3 26 103
use INVX2  INVX2_57
timestamp 1625156677
transform -1 0 2324 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_171
timestamp 1625156677
transform -1 0 2348 0 -1 1905
box -2 -3 26 103
use AND2X2  AND2X2_96
timestamp 1625156677
transform -1 0 2380 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_314
timestamp 1625156677
transform 1 0 2380 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_4_0
timestamp 1625156677
transform 1 0 2404 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_4_1
timestamp 1625156677
transform 1 0 2412 0 -1 1905
box -2 -3 10 103
use NAND2X1  NAND2X1_648
timestamp 1625156677
transform 1 0 2420 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_374
timestamp 1625156677
transform 1 0 2444 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_287
timestamp 1625156677
transform -1 0 2508 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_286
timestamp 1625156677
transform -1 0 2540 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_288
timestamp 1625156677
transform -1 0 2572 0 -1 1905
box -2 -3 34 103
use OR2X2  OR2X2_125
timestamp 1625156677
transform -1 0 2604 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_275
timestamp 1625156677
transform -1 0 2636 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_274
timestamp 1625156677
transform -1 0 2668 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_174
timestamp 1625156677
transform -1 0 2692 0 -1 1905
box -2 -3 26 103
use AND2X2  AND2X2_97
timestamp 1625156677
transform -1 0 2724 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_589
timestamp 1625156677
transform -1 0 2756 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_350
timestamp 1625156677
transform -1 0 2788 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_493
timestamp 1625156677
transform -1 0 2804 0 -1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_370
timestamp 1625156677
transform -1 0 2836 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_639
timestamp 1625156677
transform -1 0 2860 0 -1 1905
box -2 -3 26 103
use AND2X2  AND2X2_49
timestamp 1625156677
transform 1 0 2860 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_94
timestamp 1625156677
transform -1 0 2916 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_5_0
timestamp 1625156677
transform 1 0 2916 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_5_1
timestamp 1625156677
transform 1 0 2924 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_138
timestamp 1625156677
transform 1 0 2932 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_139
timestamp 1625156677
transform 1 0 2964 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1625156677
transform -1 0 3092 0 -1 1905
box -2 -3 98 103
use NAND2X1  NAND2X1_160
timestamp 1625156677
transform 1 0 3092 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_165
timestamp 1625156677
transform 1 0 3116 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_168
timestamp 1625156677
transform 1 0 3140 0 -1 1905
box -2 -3 26 103
use OR2X2  OR2X2_64
timestamp 1625156677
transform 1 0 3164 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_169
timestamp 1625156677
transform 1 0 3196 0 -1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1625156677
transform -1 0 3316 0 -1 1905
box -2 -3 98 103
use NAND3X1  NAND3X1_148
timestamp 1625156677
transform -1 0 3348 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_97
timestamp 1625156677
transform 1 0 3348 0 -1 1905
box -2 -3 18 103
use INVX1  INVX1_98
timestamp 1625156677
transform 1 0 3364 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_143
timestamp 1625156677
transform -1 0 3412 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_6_0
timestamp 1625156677
transform 1 0 3412 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_6_1
timestamp 1625156677
transform 1 0 3420 0 -1 1905
box -2 -3 10 103
use NAND2X1  NAND2X1_171
timestamp 1625156677
transform 1 0 3428 0 -1 1905
box -2 -3 26 103
use XOR2X1  XOR2X1_89
timestamp 1625156677
transform 1 0 3452 0 -1 1905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1625156677
transform 1 0 3508 0 -1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1625156677
transform -1 0 3700 0 -1 1905
box -2 -3 98 103
use INVX2  INVX2_47
timestamp 1625156677
transform 1 0 3700 0 -1 1905
box -2 -3 18 103
use AND2X2  AND2X2_166
timestamp 1625156677
transform 1 0 3716 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_219
timestamp 1625156677
transform 1 0 3748 0 -1 1905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_233
timestamp 1625156677
transform 1 0 3844 0 -1 1905
box -2 -3 98 103
use FILL  FILL_18_7_0
timestamp 1625156677
transform 1 0 3940 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_7_1
timestamp 1625156677
transform 1 0 3948 0 -1 1905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_221
timestamp 1625156677
transform 1 0 3956 0 -1 1905
box -2 -3 98 103
use XNOR2X1  XNOR2X1_113
timestamp 1625156677
transform -1 0 4108 0 -1 1905
box -2 -3 58 103
use XOR2X1  XOR2X1_141
timestamp 1625156677
transform -1 0 4164 0 -1 1905
box -2 -3 58 103
use NAND2X1  NAND2X1_249
timestamp 1625156677
transform 1 0 4164 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_221
timestamp 1625156677
transform 1 0 4188 0 -1 1905
box -2 -3 34 103
use OR2X2  OR2X2_97
timestamp 1625156677
transform -1 0 4252 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_143
timestamp 1625156677
transform 1 0 4252 0 -1 1905
box -2 -3 18 103
use AND2X2  AND2X2_74
timestamp 1625156677
transform 1 0 4268 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_212
timestamp 1625156677
transform 1 0 4300 0 -1 1905
box -2 -3 34 103
use NOR3X1  NOR3X1_49
timestamp 1625156677
transform 1 0 4332 0 -1 1905
box -2 -3 66 103
use NOR2X1  NOR2X1_138
timestamp 1625156677
transform -1 0 4420 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_155
timestamp 1625156677
transform -1 0 4452 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_8_0
timestamp 1625156677
transform 1 0 4452 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_8_1
timestamp 1625156677
transform 1 0 4460 0 -1 1905
box -2 -3 10 103
use NAND3X1  NAND3X1_223
timestamp 1625156677
transform 1 0 4468 0 -1 1905
box -2 -3 34 103
use OR2X2  OR2X2_98
timestamp 1625156677
transform -1 0 4532 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_145
timestamp 1625156677
transform 1 0 4532 0 -1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_227
timestamp 1625156677
transform 1 0 4548 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_226
timestamp 1625156677
transform 1 0 4580 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_140
timestamp 1625156677
transform 1 0 4612 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_158
timestamp 1625156677
transform -1 0 4668 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_254
timestamp 1625156677
transform -1 0 4692 0 -1 1905
box -2 -3 26 103
use OR2X2  OR2X2_99
timestamp 1625156677
transform -1 0 4724 0 -1 1905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_112
timestamp 1625156677
transform 1 0 4724 0 -1 1905
box -2 -3 58 103
use XOR2X1  XOR2X1_112
timestamp 1625156677
transform -1 0 4836 0 -1 1905
box -2 -3 58 103
use XOR2X1  XOR2X1_108
timestamp 1625156677
transform 1 0 4836 0 -1 1905
box -2 -3 58 103
use XOR2X1  XOR2X1_109
timestamp 1625156677
transform 1 0 4892 0 -1 1905
box -2 -3 58 103
use FILL  FILL_18_9_0
timestamp 1625156677
transform -1 0 4956 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_9_1
timestamp 1625156677
transform -1 0 4964 0 -1 1905
box -2 -3 10 103
use XOR2X1  XOR2X1_121
timestamp 1625156677
transform -1 0 5020 0 -1 1905
box -2 -3 58 103
use XOR2X1  XOR2X1_96
timestamp 1625156677
transform -1 0 5076 0 -1 1905
box -2 -3 58 103
use XOR2X1  XOR2X1_116
timestamp 1625156677
transform -1 0 5132 0 -1 1905
box -2 -3 58 103
use BUFX2  BUFX2_274
timestamp 1625156677
transform 1 0 5132 0 -1 1905
box -2 -3 26 103
use OR2X2  OR2X2_84
timestamp 1625156677
transform 1 0 5156 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_136
timestamp 1625156677
transform 1 0 5188 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_194
timestamp 1625156677
transform -1 0 5252 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_192
timestamp 1625156677
transform -1 0 5284 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_124
timestamp 1625156677
transform -1 0 5300 0 -1 1905
box -2 -3 18 103
use FILL  FILL_19_1
timestamp 1625156677
transform -1 0 5308 0 -1 1905
box -2 -3 10 103
use FILL  FILL_19_2
timestamp 1625156677
transform -1 0 5316 0 -1 1905
box -2 -3 10 103
use INVX1  INVX1_253
timestamp 1625156677
transform -1 0 20 0 1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_336
timestamp 1625156677
transform -1 0 52 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_251
timestamp 1625156677
transform -1 0 68 0 1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_337
timestamp 1625156677
transform 1 0 68 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_346
timestamp 1625156677
transform -1 0 132 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_252
timestamp 1625156677
transform -1 0 148 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_345
timestamp 1625156677
transform 1 0 148 0 1 1705
box -2 -3 34 103
use XOR2X1  XOR2X1_194
timestamp 1625156677
transform 1 0 180 0 1 1705
box -2 -3 58 103
use NOR2X1  NOR2X1_202
timestamp 1625156677
transform 1 0 236 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_362
timestamp 1625156677
transform -1 0 284 0 1 1705
box -2 -3 26 103
use AND2X2  AND2X2_106
timestamp 1625156677
transform 1 0 284 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_363
timestamp 1625156677
transform -1 0 340 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_0_0
timestamp 1625156677
transform 1 0 340 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1625156677
transform 1 0 348 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_318
timestamp 1625156677
transform 1 0 356 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_225
timestamp 1625156677
transform -1 0 404 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_235
timestamp 1625156677
transform 1 0 404 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_371
timestamp 1625156677
transform 1 0 428 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_413
timestamp 1625156677
transform -1 0 484 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_277
timestamp 1625156677
transform -1 0 500 0 1 1705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_166
timestamp 1625156677
transform 1 0 500 0 1 1705
box -2 -3 58 103
use XOR2X1  XOR2X1_185
timestamp 1625156677
transform -1 0 612 0 1 1705
box -2 -3 58 103
use CLKBUF1  CLKBUF1_27
timestamp 1625156677
transform 1 0 612 0 1 1705
box -2 -3 74 103
use NOR2X1  NOR2X1_194
timestamp 1625156677
transform 1 0 684 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_216
timestamp 1625156677
transform -1 0 740 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_309
timestamp 1625156677
transform -1 0 772 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_303
timestamp 1625156677
transform -1 0 804 0 1 1705
box -2 -3 34 103
use NOR3X1  NOR3X1_59
timestamp 1625156677
transform 1 0 804 0 1 1705
box -2 -3 66 103
use FILL  FILL_17_1_0
timestamp 1625156677
transform 1 0 868 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1625156677
transform 1 0 876 0 1 1705
box -2 -3 10 103
use NAND3X1  NAND3X1_309
timestamp 1625156677
transform 1 0 884 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_211
timestamp 1625156677
transform 1 0 916 0 1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_213
timestamp 1625156677
transform -1 0 964 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_306
timestamp 1625156677
transform 1 0 964 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_308
timestamp 1625156677
transform 1 0 996 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_305
timestamp 1625156677
transform 1 0 1028 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_210
timestamp 1625156677
transform -1 0 1076 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_349
timestamp 1625156677
transform 1 0 1076 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_195
timestamp 1625156677
transform -1 0 1124 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_348
timestamp 1625156677
transform -1 0 1148 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_289
timestamp 1625156677
transform -1 0 1244 0 1 1705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_17
timestamp 1625156677
transform -1 0 1316 0 1 1705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_298
timestamp 1625156677
transform -1 0 1412 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_2_0
timestamp 1625156677
transform -1 0 1420 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1625156677
transform -1 0 1428 0 1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_288
timestamp 1625156677
transform -1 0 1524 0 1 1705
box -2 -3 98 103
use BUFX2  BUFX2_180
timestamp 1625156677
transform -1 0 1548 0 1 1705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_215
timestamp 1625156677
transform 1 0 1548 0 1 1705
box -2 -3 58 103
use INVX1  INVX1_553
timestamp 1625156677
transform -1 0 1620 0 1 1705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_211
timestamp 1625156677
transform 1 0 1620 0 1 1705
box -2 -3 58 103
use NAND2X1  NAND2X1_653
timestamp 1625156677
transform 1 0 1676 0 1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_506
timestamp 1625156677
transform 1 0 1700 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_667
timestamp 1625156677
transform -1 0 1756 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_562
timestamp 1625156677
transform -1 0 1772 0 1 1705
box -2 -3 18 103
use INVX1  INVX1_545
timestamp 1625156677
transform -1 0 1788 0 1 1705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_222
timestamp 1625156677
transform 1 0 1788 0 1 1705
box -2 -3 58 103
use INVX1  INVX1_576
timestamp 1625156677
transform 1 0 1844 0 1 1705
box -2 -3 18 103
use FILL  FILL_17_3_0
timestamp 1625156677
transform 1 0 1860 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1625156677
transform 1 0 1868 0 1 1705
box -2 -3 10 103
use XNOR2X1  XNOR2X1_216
timestamp 1625156677
transform 1 0 1876 0 1 1705
box -2 -3 58 103
use INVX2  INVX2_88
timestamp 1625156677
transform -1 0 1948 0 1 1705
box -2 -3 18 103
use BUFX2  BUFX2_181
timestamp 1625156677
transform 1 0 1948 0 1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_525
timestamp 1625156677
transform 1 0 1972 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_646
timestamp 1625156677
transform -1 0 2028 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_503
timestamp 1625156677
transform -1 0 2044 0 1 1705
box -2 -3 18 103
use XOR2X1  XOR2X1_160
timestamp 1625156677
transform 1 0 2044 0 1 1705
box -2 -3 58 103
use NAND3X1  NAND3X1_527
timestamp 1625156677
transform -1 0 2132 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_543
timestamp 1625156677
transform -1 0 2148 0 1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_202
timestamp 1625156677
transform 1 0 2148 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_313
timestamp 1625156677
transform -1 0 2204 0 1 1705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_144
timestamp 1625156677
transform 1 0 2204 0 1 1705
box -2 -3 58 103
use NAND3X1  NAND3X1_290
timestamp 1625156677
transform -1 0 2292 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_58
timestamp 1625156677
transform -1 0 2308 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_273
timestamp 1625156677
transform 1 0 2308 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_277
timestamp 1625156677
transform 1 0 2340 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_181
timestamp 1625156677
transform 1 0 2372 0 1 1705
box -2 -3 18 103
use FILL  FILL_17_4_0
timestamp 1625156677
transform -1 0 2396 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_4_1
timestamp 1625156677
transform -1 0 2404 0 1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_175
timestamp 1625156677
transform -1 0 2428 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_197
timestamp 1625156677
transform -1 0 2460 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_316
timestamp 1625156677
transform -1 0 2484 0 1 1705
box -2 -3 26 103
use OR2X2  OR2X2_126
timestamp 1625156677
transform -1 0 2516 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_198
timestamp 1625156677
transform -1 0 2548 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_289
timestamp 1625156677
transform -1 0 2580 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_317
timestamp 1625156677
transform -1 0 2604 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_626
timestamp 1625156677
transform 1 0 2604 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_180
timestamp 1625156677
transform -1 0 2652 0 1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_386
timestamp 1625156677
transform -1 0 2684 0 1 1705
box -2 -3 34 103
use OR2X2  OR2X2_142
timestamp 1625156677
transform -1 0 2716 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_623
timestamp 1625156677
transform -1 0 2748 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_410
timestamp 1625156677
transform 1 0 2748 0 1 1705
box -2 -3 26 103
use XOR2X1  XOR2X1_298
timestamp 1625156677
transform 1 0 2772 0 1 1705
box -2 -3 58 103
use OR2X2  OR2X2_131
timestamp 1625156677
transform -1 0 2860 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_638
timestamp 1625156677
transform -1 0 2884 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_124
timestamp 1625156677
transform -1 0 2908 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_5_0
timestamp 1625156677
transform 1 0 2908 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_5_1
timestamp 1625156677
transform 1 0 2916 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_163
timestamp 1625156677
transform 1 0 2924 0 1 1705
box -2 -3 26 103
use OR2X2  OR2X2_61
timestamp 1625156677
transform 1 0 2948 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_92
timestamp 1625156677
transform 1 0 2980 0 1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_144
timestamp 1625156677
transform 1 0 2996 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_142
timestamp 1625156677
transform 1 0 3028 0 1 1705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_145
timestamp 1625156677
transform 1 0 3060 0 1 1705
box -2 -3 58 103
use XOR2X1  XOR2X1_148
timestamp 1625156677
transform -1 0 3172 0 1 1705
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1625156677
transform -1 0 3268 0 1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1625156677
transform -1 0 3364 0 1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1625156677
transform 1 0 3364 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_6_0
timestamp 1625156677
transform 1 0 3460 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_6_1
timestamp 1625156677
transform 1 0 3468 0 1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_366
timestamp 1625156677
transform 1 0 3476 0 1 1705
box -2 -3 26 103
use INVX2  INVX2_76
timestamp 1625156677
transform 1 0 3500 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_400
timestamp 1625156677
transform 1 0 3516 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_367
timestamp 1625156677
transform 1 0 3540 0 1 1705
box -2 -3 26 103
use BUFX2  BUFX2_266
timestamp 1625156677
transform 1 0 3564 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_625
timestamp 1625156677
transform 1 0 3588 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1625156677
transform -1 0 3708 0 1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_336
timestamp 1625156677
transform 1 0 3708 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_579
timestamp 1625156677
transform -1 0 3772 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_624
timestamp 1625156677
transform -1 0 3796 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_337
timestamp 1625156677
transform -1 0 3828 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_479
timestamp 1625156677
transform 1 0 3828 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_368
timestamp 1625156677
transform -1 0 3868 0 1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1625156677
transform 1 0 3868 0 1 1705
box -2 -3 98 103
use FILL  FILL_17_7_0
timestamp 1625156677
transform 1 0 3964 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_7_1
timestamp 1625156677
transform 1 0 3972 0 1 1705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_14
timestamp 1625156677
transform 1 0 3980 0 1 1705
box -2 -3 74 103
use INVX1  INVX1_160
timestamp 1625156677
transform 1 0 4052 0 1 1705
box -2 -3 18 103
use XOR2X1  XOR2X1_136
timestamp 1625156677
transform -1 0 4124 0 1 1705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_114
timestamp 1625156677
transform 1 0 4124 0 1 1705
box -2 -3 58 103
use NAND2X1  NAND2X1_248
timestamp 1625156677
transform 1 0 4180 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_165
timestamp 1625156677
transform 1 0 4204 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_250
timestamp 1625156677
transform -1 0 4260 0 1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_222
timestamp 1625156677
transform -1 0 4292 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_252
timestamp 1625156677
transform -1 0 4316 0 1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_224
timestamp 1625156677
transform -1 0 4348 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_225
timestamp 1625156677
transform 1 0 4348 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_215
timestamp 1625156677
transform -1 0 4412 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_213
timestamp 1625156677
transform -1 0 4444 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_8_0
timestamp 1625156677
transform -1 0 4452 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_8_1
timestamp 1625156677
transform -1 0 4460 0 1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_159
timestamp 1625156677
transform -1 0 4492 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_143
timestamp 1625156677
transform 1 0 4492 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_157
timestamp 1625156677
transform -1 0 4548 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_156
timestamp 1625156677
transform -1 0 4580 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_217
timestamp 1625156677
transform -1 0 4612 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_218
timestamp 1625156677
transform 1 0 4612 0 1 1705
box -2 -3 34 103
use AND2X2  AND2X2_78
timestamp 1625156677
transform -1 0 4676 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_257
timestamp 1625156677
transform -1 0 4700 0 1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_231
timestamp 1625156677
transform -1 0 4732 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_229
timestamp 1625156677
transform 1 0 4732 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_220
timestamp 1625156677
transform -1 0 4796 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_219
timestamp 1625156677
transform 1 0 4796 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_142
timestamp 1625156677
transform 1 0 4828 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_146
timestamp 1625156677
transform 1 0 4852 0 1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_228
timestamp 1625156677
transform 1 0 4868 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_230
timestamp 1625156677
transform 1 0 4900 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_160
timestamp 1625156677
transform 1 0 4932 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_9_0
timestamp 1625156677
transform -1 0 4972 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_9_1
timestamp 1625156677
transform -1 0 4980 0 1 1705
box -2 -3 10 103
use OR2X2  OR2X2_100
timestamp 1625156677
transform -1 0 5012 0 1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_222
timestamp 1625156677
transform -1 0 5108 0 1 1705
box -2 -3 98 103
use XOR2X1  XOR2X1_117
timestamp 1625156677
transform -1 0 5164 0 1 1705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_99
timestamp 1625156677
transform -1 0 5220 0 1 1705
box -2 -3 58 103
use OAI21X1  OAI21X1_188
timestamp 1625156677
transform -1 0 5252 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_43
timestamp 1625156677
transform -1 0 5268 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_227
timestamp 1625156677
transform 1 0 5268 0 1 1705
box -2 -3 26 103
use FILL  FILL_18_1
timestamp 1625156677
transform 1 0 5292 0 1 1705
box -2 -3 10 103
use FILL  FILL_18_2
timestamp 1625156677
transform 1 0 5300 0 1 1705
box -2 -3 10 103
use FILL  FILL_18_3
timestamp 1625156677
transform 1 0 5308 0 1 1705
box -2 -3 10 103
use BUFX2  BUFX2_194
timestamp 1625156677
transform -1 0 28 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_190
timestamp 1625156677
transform -1 0 52 0 -1 1705
box -2 -3 26 103
use XOR2X1  XOR2X1_193
timestamp 1625156677
transform -1 0 108 0 -1 1705
box -2 -3 58 103
use XOR2X1  XOR2X1_184
timestamp 1625156677
transform -1 0 164 0 -1 1705
box -2 -3 58 103
use XOR2X1  XOR2X1_171
timestamp 1625156677
transform 1 0 164 0 -1 1705
box -2 -3 58 103
use AND2X2  AND2X2_108
timestamp 1625156677
transform -1 0 252 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_319
timestamp 1625156677
transform 1 0 252 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_364
timestamp 1625156677
transform -1 0 308 0 -1 1705
box -2 -3 26 103
use AND2X2  AND2X2_107
timestamp 1625156677
transform 1 0 308 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_0_0
timestamp 1625156677
transform -1 0 348 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1625156677
transform -1 0 356 0 -1 1705
box -2 -3 10 103
use INVX1  INVX1_226
timestamp 1625156677
transform -1 0 372 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_203
timestamp 1625156677
transform 1 0 372 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_319
timestamp 1625156677
transform -1 0 428 0 -1 1705
box -2 -3 34 103
use XOR2X1  XOR2X1_172
timestamp 1625156677
transform -1 0 484 0 -1 1705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_153
timestamp 1625156677
transform 1 0 484 0 -1 1705
box -2 -3 58 103
use NAND2X1  NAND2X1_395
timestamp 1625156677
transform -1 0 564 0 -1 1705
box -2 -3 26 103
use XOR2X1  XOR2X1_179
timestamp 1625156677
transform 1 0 564 0 -1 1705
box -2 -3 58 103
use OAI21X1  OAI21X1_310
timestamp 1625156677
transform 1 0 620 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_355
timestamp 1625156677
transform 1 0 652 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_196
timestamp 1625156677
transform -1 0 700 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_197
timestamp 1625156677
transform 1 0 700 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_182
timestamp 1625156677
transform -1 0 748 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_316
timestamp 1625156677
transform 1 0 748 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_211
timestamp 1625156677
transform -1 0 812 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_212
timestamp 1625156677
transform -1 0 828 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_360
timestamp 1625156677
transform -1 0 852 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_1_0
timestamp 1625156677
transform -1 0 860 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_1
timestamp 1625156677
transform -1 0 868 0 -1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_217
timestamp 1625156677
transform -1 0 900 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_353
timestamp 1625156677
transform -1 0 924 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_212
timestamp 1625156677
transform -1 0 956 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_316
timestamp 1625156677
transform 1 0 956 0 -1 1705
box -2 -3 34 103
use XOR2X1  XOR2X1_165
timestamp 1625156677
transform -1 0 1044 0 -1 1705
box -2 -3 58 103
use INVX1  INVX1_213
timestamp 1625156677
transform 1 0 1044 0 -1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_311
timestamp 1625156677
transform -1 0 1092 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_310
timestamp 1625156677
transform 1 0 1092 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_215
timestamp 1625156677
transform -1 0 1140 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_308
timestamp 1625156677
transform -1 0 1172 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_214
timestamp 1625156677
transform -1 0 1188 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_307
timestamp 1625156677
transform -1 0 1220 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_261
timestamp 1625156677
transform -1 0 1316 0 -1 1705
box -2 -3 98 103
use INVX1  INVX1_517
timestamp 1625156677
transform -1 0 1332 0 -1 1705
box -2 -3 18 103
use XOR2X1  XOR2X1_300
timestamp 1625156677
transform 1 0 1332 0 -1 1705
box -2 -3 58 103
use FILL  FILL_16_2_0
timestamp 1625156677
transform -1 0 1396 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1625156677
transform -1 0 1404 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_250
timestamp 1625156677
transform -1 0 1500 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_297
timestamp 1625156677
transform -1 0 1596 0 -1 1705
box -2 -3 98 103
use XOR2X1  XOR2X1_166
timestamp 1625156677
transform -1 0 1652 0 -1 1705
box -2 -3 58 103
use NOR2X1  NOR2X1_408
timestamp 1625156677
transform 1 0 1652 0 -1 1705
box -2 -3 26 103
use AND2X2  AND2X2_176
timestamp 1625156677
transform 1 0 1676 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_611
timestamp 1625156677
transform 1 0 1708 0 -1 1705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_231
timestamp 1625156677
transform -1 0 1796 0 -1 1705
box -2 -3 58 103
use NOR2X1  NOR2X1_426
timestamp 1625156677
transform -1 0 1820 0 -1 1705
box -2 -3 26 103
use XOR2X1  XOR2X1_304
timestamp 1625156677
transform 1 0 1820 0 -1 1705
box -2 -3 58 103
use FILL  FILL_16_3_0
timestamp 1625156677
transform -1 0 1884 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_1
timestamp 1625156677
transform -1 0 1892 0 -1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_375
timestamp 1625156677
transform -1 0 1924 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_610
timestamp 1625156677
transform 1 0 1924 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_533
timestamp 1625156677
transform -1 0 1972 0 -1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_373
timestamp 1625156677
transform -1 0 2004 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_645
timestamp 1625156677
transform -1 0 2028 0 -1 1705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_230
timestamp 1625156677
transform -1 0 2084 0 -1 1705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_143
timestamp 1625156677
transform 1 0 2084 0 -1 1705
box -2 -3 58 103
use NAND2X1  NAND2X1_322
timestamp 1625156677
transform -1 0 2164 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_276
timestamp 1625156677
transform 1 0 2164 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_176
timestamp 1625156677
transform -1 0 2220 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_278
timestamp 1625156677
transform 1 0 2220 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_183
timestamp 1625156677
transform -1 0 2268 0 -1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_199
timestamp 1625156677
transform 1 0 2268 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_321
timestamp 1625156677
transform -1 0 2324 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_320
timestamp 1625156677
transform -1 0 2348 0 -1 1705
box -2 -3 26 103
use OR2X2  OR2X2_128
timestamp 1625156677
transform -1 0 2380 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_647
timestamp 1625156677
transform -1 0 2404 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_4_0
timestamp 1625156677
transform 1 0 2404 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_4_1
timestamp 1625156677
transform 1 0 2412 0 -1 1705
box -2 -3 10 103
use OR2X2  OR2X2_134
timestamp 1625156677
transform 1 0 2420 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_319
timestamp 1625156677
transform -1 0 2476 0 -1 1705
box -2 -3 26 103
use OR2X2  OR2X2_127
timestamp 1625156677
transform -1 0 2508 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_318
timestamp 1625156677
transform 1 0 2508 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_507
timestamp 1625156677
transform -1 0 2548 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_431
timestamp 1625156677
transform 1 0 2548 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_657
timestamp 1625156677
transform -1 0 2596 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_390
timestamp 1625156677
transform -1 0 2628 0 -1 1705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_214
timestamp 1625156677
transform 1 0 2628 0 -1 1705
box -2 -3 58 103
use NAND3X1  NAND3X1_510
timestamp 1625156677
transform 1 0 2684 0 -1 1705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_183
timestamp 1625156677
transform 1 0 2716 0 -1 1705
box -2 -3 98 103
use XOR2X1  XOR2X1_65
timestamp 1625156677
transform 1 0 2812 0 -1 1705
box -2 -3 58 103
use FILL  FILL_16_5_0
timestamp 1625156677
transform 1 0 2868 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_5_1
timestamp 1625156677
transform 1 0 2876 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_181
timestamp 1625156677
transform 1 0 2884 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1625156677
transform -1 0 3076 0 -1 1705
box -2 -3 98 103
use AND2X2  AND2X2_162
timestamp 1625156677
transform -1 0 3108 0 -1 1705
box -2 -3 34 103
use BUFX2  BUFX2_170
timestamp 1625156677
transform -1 0 3132 0 -1 1705
box -2 -3 26 103
use XOR2X1  XOR2X1_149
timestamp 1625156677
transform -1 0 3188 0 -1 1705
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1625156677
transform -1 0 3284 0 -1 1705
box -2 -3 98 103
use AND2X2  AND2X2_165
timestamp 1625156677
transform -1 0 3316 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_363
timestamp 1625156677
transform -1 0 3340 0 -1 1705
box -2 -3 26 103
use AND2X2  AND2X2_170
timestamp 1625156677
transform -1 0 3372 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_334
timestamp 1625156677
transform -1 0 3404 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_6_0
timestamp 1625156677
transform 1 0 3404 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_6_1
timestamp 1625156677
transform 1 0 3412 0 -1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_335
timestamp 1625156677
transform 1 0 3420 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_401
timestamp 1625156677
transform 1 0 3452 0 -1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_494
timestamp 1625156677
transform -1 0 3508 0 -1 1705
box -2 -3 34 103
use INVX2  INVX2_75
timestamp 1625156677
transform -1 0 3524 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_577
timestamp 1625156677
transform -1 0 3556 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_578
timestamp 1625156677
transform 1 0 3556 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_402
timestamp 1625156677
transform -1 0 3612 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_490
timestamp 1625156677
transform 1 0 3612 0 -1 1705
box -2 -3 18 103
use AND2X2  AND2X2_171
timestamp 1625156677
transform 1 0 3628 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_626
timestamp 1625156677
transform 1 0 3660 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_627
timestamp 1625156677
transform -1 0 3708 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1625156677
transform -1 0 3804 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_223
timestamp 1625156677
transform 1 0 3804 0 -1 1705
box -2 -3 98 103
use FILL  FILL_16_7_0
timestamp 1625156677
transform 1 0 3900 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_7_1
timestamp 1625156677
transform 1 0 3908 0 -1 1705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_232
timestamp 1625156677
transform 1 0 3916 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1625156677
transform -1 0 4108 0 -1 1705
box -2 -3 98 103
use XOR2X1  XOR2X1_130
timestamp 1625156677
transform 1 0 4108 0 -1 1705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_115
timestamp 1625156677
transform 1 0 4164 0 -1 1705
box -2 -3 58 103
use NAND3X1  NAND3X1_237
timestamp 1625156677
transform 1 0 4220 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_216
timestamp 1625156677
transform -1 0 4284 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_253
timestamp 1625156677
transform 1 0 4284 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_221
timestamp 1625156677
transform 1 0 4308 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_151
timestamp 1625156677
transform 1 0 4340 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_141
timestamp 1625156677
transform -1 0 4380 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_164
timestamp 1625156677
transform -1 0 4412 0 -1 1705
box -2 -3 34 103
use INVX2  INVX2_48
timestamp 1625156677
transform -1 0 4428 0 -1 1705
box -2 -3 18 103
use FILL  FILL_16_8_0
timestamp 1625156677
transform 1 0 4428 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_8_1
timestamp 1625156677
transform 1 0 4436 0 -1 1705
box -2 -3 10 103
use XNOR2X1  XNOR2X1_116
timestamp 1625156677
transform 1 0 4444 0 -1 1705
box -2 -3 58 103
use NAND2X1  NAND2X1_256
timestamp 1625156677
transform 1 0 4500 0 -1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_236
timestamp 1625156677
transform 1 0 4524 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_222
timestamp 1625156677
transform -1 0 4588 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_161
timestamp 1625156677
transform -1 0 4620 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_259
timestamp 1625156677
transform -1 0 4644 0 -1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_233
timestamp 1625156677
transform -1 0 4676 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_223
timestamp 1625156677
transform -1 0 4708 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_224
timestamp 1625156677
transform 1 0 4708 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_147
timestamp 1625156677
transform -1 0 4756 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_144
timestamp 1625156677
transform 1 0 4756 0 -1 1705
box -2 -3 26 103
use AND2X2  AND2X2_79
timestamp 1625156677
transform -1 0 4812 0 -1 1705
box -2 -3 34 103
use AND2X2  AND2X2_77
timestamp 1625156677
transform -1 0 4844 0 -1 1705
box -2 -3 34 103
use BUFX2  BUFX2_158
timestamp 1625156677
transform 1 0 4844 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_255
timestamp 1625156677
transform 1 0 4868 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_202
timestamp 1625156677
transform 1 0 4892 0 -1 1705
box -2 -3 98 103
use FILL  FILL_16_9_0
timestamp 1625156677
transform 1 0 4988 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_9_1
timestamp 1625156677
transform 1 0 4996 0 -1 1705
box -2 -3 10 103
use INVX2  INVX2_41
timestamp 1625156677
transform 1 0 5004 0 -1 1705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_95
timestamp 1625156677
transform -1 0 5076 0 -1 1705
box -2 -3 58 103
use OAI21X1  OAI21X1_192
timestamp 1625156677
transform -1 0 5108 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_126
timestamp 1625156677
transform 1 0 5108 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_125
timestamp 1625156677
transform -1 0 5148 0 -1 1705
box -2 -3 26 103
use OR2X2  OR2X2_86
timestamp 1625156677
transform -1 0 5180 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_138
timestamp 1625156677
transform -1 0 5212 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_137
timestamp 1625156677
transform -1 0 5244 0 -1 1705
box -2 -3 34 103
use XOR2X1  XOR2X1_95
timestamp 1625156677
transform 1 0 5244 0 -1 1705
box -2 -3 58 103
use FILL  FILL_17_1
timestamp 1625156677
transform -1 0 5308 0 -1 1705
box -2 -3 10 103
use FILL  FILL_17_2
timestamp 1625156677
transform -1 0 5316 0 -1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_204
timestamp 1625156677
transform 1 0 4 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_321
timestamp 1625156677
transform 1 0 28 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_373
timestamp 1625156677
transform 1 0 60 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_222
timestamp 1625156677
transform 1 0 84 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_332
timestamp 1625156677
transform 1 0 116 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_227
timestamp 1625156677
transform -1 0 164 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_365
timestamp 1625156677
transform 1 0 164 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_366
timestamp 1625156677
transform 1 0 188 0 1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_320
timestamp 1625156677
transform 1 0 212 0 1 1505
box -2 -3 34 103
use NOR3X1  NOR3X1_62
timestamp 1625156677
transform -1 0 308 0 1 1505
box -2 -3 66 103
use OAI21X1  OAI21X1_320
timestamp 1625156677
transform -1 0 340 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_0_0
timestamp 1625156677
transform 1 0 340 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1625156677
transform 1 0 348 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_323
timestamp 1625156677
transform 1 0 356 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_61
timestamp 1625156677
transform 1 0 388 0 1 1505
box -2 -3 18 103
use BUFX2  BUFX2_189
timestamp 1625156677
transform -1 0 428 0 1 1505
box -2 -3 26 103
use XOR2X1  XOR2X1_195
timestamp 1625156677
transform -1 0 484 0 1 1505
box -2 -3 58 103
use XOR2X1  XOR2X1_173
timestamp 1625156677
transform -1 0 540 0 1 1505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_163
timestamp 1625156677
transform 1 0 540 0 1 1505
box -2 -3 58 103
use NOR2X1  NOR2X1_223
timestamp 1625156677
transform -1 0 620 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_394
timestamp 1625156677
transform -1 0 644 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_352
timestamp 1625156677
transform 1 0 644 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_258
timestamp 1625156677
transform -1 0 692 0 1 1505
box -2 -3 18 103
use AND2X2  AND2X2_105
timestamp 1625156677
transform -1 0 724 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_315
timestamp 1625156677
transform 1 0 724 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_222
timestamp 1625156677
transform -1 0 772 0 1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_218
timestamp 1625156677
transform -1 0 804 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_317
timestamp 1625156677
transform 1 0 804 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_223
timestamp 1625156677
transform -1 0 852 0 1 1505
box -2 -3 18 103
use FILL  FILL_15_1_0
timestamp 1625156677
transform -1 0 860 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_1
timestamp 1625156677
transform -1 0 868 0 1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_312
timestamp 1625156677
transform -1 0 900 0 1 1505
box -2 -3 34 103
use AOI22X1  AOI22X1_9
timestamp 1625156677
transform -1 0 940 0 1 1505
box -2 -3 42 103
use NAND3X1  NAND3X1_314
timestamp 1625156677
transform 1 0 940 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_217
timestamp 1625156677
transform -1 0 988 0 1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_313
timestamp 1625156677
transform 1 0 988 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_352
timestamp 1625156677
transform -1 0 1044 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_351
timestamp 1625156677
transform -1 0 1068 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_216
timestamp 1625156677
transform 1 0 1068 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_311
timestamp 1625156677
transform -1 0 1116 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_198
timestamp 1625156677
transform -1 0 1140 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_312
timestamp 1625156677
transform -1 0 1172 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_269
timestamp 1625156677
transform -1 0 1268 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_262
timestamp 1625156677
transform -1 0 1364 0 1 1505
box -2 -3 98 103
use FILL  FILL_15_2_0
timestamp 1625156677
transform -1 0 1372 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1625156677
transform -1 0 1380 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_270
timestamp 1625156677
transform -1 0 1476 0 1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_414
timestamp 1625156677
transform 1 0 1476 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_520
timestamp 1625156677
transform -1 0 1516 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_263
timestamp 1625156677
transform -1 0 1612 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_523
timestamp 1625156677
transform -1 0 1628 0 1 1505
box -2 -3 18 103
use XOR2X1  XOR2X1_167
timestamp 1625156677
transform -1 0 1684 0 1 1505
box -2 -3 58 103
use OAI21X1  OAI21X1_617
timestamp 1625156677
transform -1 0 1716 0 1 1505
box -2 -3 34 103
use AND2X2  AND2X2_180
timestamp 1625156677
transform -1 0 1748 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_420
timestamp 1625156677
transform -1 0 1772 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_678
timestamp 1625156677
transform -1 0 1796 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_619
timestamp 1625156677
transform -1 0 1828 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_389
timestamp 1625156677
transform 1 0 1828 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_629
timestamp 1625156677
transform -1 0 1892 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_3_0
timestamp 1625156677
transform 1 0 1892 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_1
timestamp 1625156677
transform 1 0 1900 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_423
timestamp 1625156677
transform 1 0 1908 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_422
timestamp 1625156677
transform -1 0 1956 0 1 1505
box -2 -3 26 103
use INVX2  INVX2_86
timestamp 1625156677
transform -1 0 1972 0 1 1505
box -2 -3 18 103
use INVX1  INVX1_532
timestamp 1625156677
transform -1 0 1988 0 1 1505
box -2 -3 18 103
use XNOR2X1  XNOR2X1_234
timestamp 1625156677
transform -1 0 2044 0 1 1505
box -2 -3 58 103
use AOI21X1  AOI21X1_359
timestamp 1625156677
transform 1 0 2044 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_598
timestamp 1625156677
transform -1 0 2108 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_618
timestamp 1625156677
transform -1 0 2140 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_421
timestamp 1625156677
transform 1 0 2140 0 1 1505
box -2 -3 26 103
use OR2X2  OR2X2_149
timestamp 1625156677
transform -1 0 2196 0 1 1505
box -2 -3 34 103
use OR2X2  OR2X2_154
timestamp 1625156677
transform 1 0 2196 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_177
timestamp 1625156677
transform -1 0 2252 0 1 1505
box -2 -3 26 103
use OR2X2  OR2X2_133
timestamp 1625156677
transform -1 0 2284 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_526
timestamp 1625156677
transform 1 0 2284 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_323
timestamp 1625156677
transform -1 0 2340 0 1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_292
timestamp 1625156677
transform -1 0 2372 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_185
timestamp 1625156677
transform 1 0 2372 0 1 1505
box -2 -3 18 103
use FILL  FILL_15_4_0
timestamp 1625156677
transform 1 0 2388 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_4_1
timestamp 1625156677
transform 1 0 2396 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_279
timestamp 1625156677
transform 1 0 2404 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_186
timestamp 1625156677
transform -1 0 2452 0 1 1505
box -2 -3 18 103
use XNOR2X1  XNOR2X1_147
timestamp 1625156677
transform -1 0 2508 0 1 1505
box -2 -3 58 103
use INVX1  INVX1_182
timestamp 1625156677
transform -1 0 2524 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_248
timestamp 1625156677
transform -1 0 2620 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_247
timestamp 1625156677
transform -1 0 2716 0 1 1505
box -2 -3 98 103
use XNOR2X1  XNOR2X1_146
timestamp 1625156677
transform 1 0 2716 0 1 1505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_226
timestamp 1625156677
transform -1 0 2828 0 1 1505
box -2 -3 58 103
use XOR2X1  XOR2X1_135
timestamp 1625156677
transform -1 0 2884 0 1 1505
box -2 -3 58 103
use BUFX2  BUFX2_169
timestamp 1625156677
transform -1 0 2908 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_5_0
timestamp 1625156677
transform -1 0 2916 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_5_1
timestamp 1625156677
transform -1 0 2924 0 1 1505
box -2 -3 10 103
use XOR2X1  XOR2X1_151
timestamp 1625156677
transform -1 0 2980 0 1 1505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_137
timestamp 1625156677
transform 1 0 2980 0 1 1505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1625156677
transform -1 0 3132 0 1 1505
box -2 -3 98 103
use AND2X2  AND2X2_161
timestamp 1625156677
transform -1 0 3164 0 1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1625156677
transform 1 0 3164 0 1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_328
timestamp 1625156677
transform 1 0 3260 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_573
timestamp 1625156677
transform -1 0 3324 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_616
timestamp 1625156677
transform -1 0 3348 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_329
timestamp 1625156677
transform -1 0 3380 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_476
timestamp 1625156677
transform -1 0 3396 0 1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_491
timestamp 1625156677
transform -1 0 3428 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_6_0
timestamp 1625156677
transform 1 0 3428 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_6_1
timestamp 1625156677
transform 1 0 3436 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_617
timestamp 1625156677
transform 1 0 3444 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1625156677
transform -1 0 3564 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1625156677
transform -1 0 3660 0 1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_618
timestamp 1625156677
transform -1 0 3684 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_391
timestamp 1625156677
transform -1 0 3708 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_392
timestamp 1625156677
transform 1 0 3708 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1625156677
transform 1 0 3732 0 1 1505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_26
timestamp 1625156677
transform -1 0 3900 0 1 1505
box -2 -3 74 103
use FILL  FILL_15_7_0
timestamp 1625156677
transform -1 0 3908 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_7_1
timestamp 1625156677
transform -1 0 3916 0 1 1505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_30
timestamp 1625156677
transform -1 0 3988 0 1 1505
box -2 -3 74 103
use BUFX4  BUFX4_3
timestamp 1625156677
transform -1 0 4020 0 1 1505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_24
timestamp 1625156677
transform 1 0 4020 0 1 1505
box -2 -3 74 103
use XOR2X1  XOR2X1_137
timestamp 1625156677
transform -1 0 4148 0 1 1505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1625156677
transform -1 0 4244 0 1 1505
box -2 -3 98 103
use XOR2X1  XOR2X1_139
timestamp 1625156677
transform -1 0 4300 0 1 1505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_136
timestamp 1625156677
transform 1 0 4300 0 1 1505
box -2 -3 58 103
use XOR2X1  XOR2X1_138
timestamp 1625156677
transform -1 0 4412 0 1 1505
box -2 -3 58 103
use AOI21X1  AOI21X1_166
timestamp 1625156677
transform 1 0 4412 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_8_0
timestamp 1625156677
transform -1 0 4452 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_8_1
timestamp 1625156677
transform -1 0 4460 0 1 1505
box -2 -3 10 103
use BUFX2  BUFX2_164
timestamp 1625156677
transform -1 0 4484 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_147
timestamp 1625156677
transform 1 0 4484 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_163
timestamp 1625156677
transform -1 0 4540 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_146
timestamp 1625156677
transform 1 0 4540 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_225
timestamp 1625156677
transform -1 0 4596 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_265
timestamp 1625156677
transform -1 0 4620 0 1 1505
box -2 -3 26 103
use INVX2  INVX2_49
timestamp 1625156677
transform 1 0 4620 0 1 1505
box -2 -3 18 103
use XNOR2X1  XNOR2X1_117
timestamp 1625156677
transform -1 0 4692 0 1 1505
box -2 -3 58 103
use NAND3X1  NAND3X1_235
timestamp 1625156677
transform -1 0 4724 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_260
timestamp 1625156677
transform 1 0 4724 0 1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_234
timestamp 1625156677
transform 1 0 4748 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_232
timestamp 1625156677
transform 1 0 4780 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_258
timestamp 1625156677
transform -1 0 4836 0 1 1505
box -2 -3 26 103
use XOR2X1  XOR2X1_119
timestamp 1625156677
transform 1 0 4836 0 1 1505
box -2 -3 58 103
use OR2X2  OR2X2_101
timestamp 1625156677
transform -1 0 4924 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_138
timestamp 1625156677
transform 1 0 4924 0 1 1505
box -2 -3 18 103
use FILL  FILL_15_9_0
timestamp 1625156677
transform 1 0 4940 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_9_1
timestamp 1625156677
transform 1 0 4948 0 1 1505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_96
timestamp 1625156677
transform 1 0 4956 0 1 1505
box -2 -3 58 103
use AOI21X1  AOI21X1_141
timestamp 1625156677
transform -1 0 5044 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_210
timestamp 1625156677
transform 1 0 5044 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_193
timestamp 1625156677
transform -1 0 5100 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_126
timestamp 1625156677
transform 1 0 5100 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_191
timestamp 1625156677
transform -1 0 5156 0 1 1505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_94
timestamp 1625156677
transform 1 0 5156 0 1 1505
box -2 -3 58 103
use NAND3X1  NAND3X1_199
timestamp 1625156677
transform -1 0 5244 0 1 1505
box -2 -3 34 103
use XOR2X1  XOR2X1_92
timestamp 1625156677
transform 1 0 5244 0 1 1505
box -2 -3 58 103
use FILL  FILL_16_1
timestamp 1625156677
transform 1 0 5300 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_2
timestamp 1625156677
transform 1 0 5308 0 1 1505
box -2 -3 10 103
use INVX1  INVX1_237
timestamp 1625156677
transform 1 0 4 0 -1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_223
timestamp 1625156677
transform -1 0 52 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_369
timestamp 1625156677
transform 1 0 52 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_328
timestamp 1625156677
transform -1 0 108 0 -1 1505
box -2 -3 34 103
use NOR3X1  NOR3X1_61
timestamp 1625156677
transform -1 0 172 0 -1 1505
box -2 -3 66 103
use OAI21X1  OAI21X1_322
timestamp 1625156677
transform 1 0 172 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_228
timestamp 1625156677
transform 1 0 204 0 -1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_328
timestamp 1625156677
transform 1 0 220 0 -1 1505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_156
timestamp 1625156677
transform -1 0 308 0 -1 1505
box -2 -3 58 103
use NOR2X1  NOR2X1_206
timestamp 1625156677
transform 1 0 308 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_205
timestamp 1625156677
transform -1 0 356 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_0_0
timestamp 1625156677
transform 1 0 356 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1625156677
transform 1 0 364 0 -1 1505
box -2 -3 10 103
use XOR2X1  XOR2X1_196
timestamp 1625156677
transform 1 0 372 0 -1 1505
box -2 -3 58 103
use BUFX2  BUFX2_184
timestamp 1625156677
transform -1 0 452 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_237
timestamp 1625156677
transform -1 0 476 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_225
timestamp 1625156677
transform 1 0 476 0 -1 1505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_162
timestamp 1625156677
transform 1 0 500 0 -1 1505
box -2 -3 58 103
use XOR2X1  XOR2X1_186
timestamp 1625156677
transform -1 0 612 0 -1 1505
box -2 -3 58 103
use NAND3X1  NAND3X1_318
timestamp 1625156677
transform -1 0 644 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_224
timestamp 1625156677
transform -1 0 660 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_317
timestamp 1625156677
transform -1 0 692 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_221
timestamp 1625156677
transform 1 0 692 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_359
timestamp 1625156677
transform -1 0 732 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_200
timestamp 1625156677
transform 1 0 732 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_358
timestamp 1625156677
transform -1 0 780 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_219
timestamp 1625156677
transform -1 0 796 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_271
timestamp 1625156677
transform -1 0 892 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_1_0
timestamp 1625156677
transform -1 0 900 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1625156677
transform -1 0 908 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_280
timestamp 1625156677
transform -1 0 1004 0 -1 1505
box -2 -3 98 103
use BUFX2  BUFX2_175
timestamp 1625156677
transform -1 0 1028 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_251
timestamp 1625156677
transform -1 0 1124 0 -1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_281
timestamp 1625156677
transform -1 0 1220 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_357
timestamp 1625156677
transform -1 0 1244 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_356
timestamp 1625156677
transform -1 0 1268 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_220
timestamp 1625156677
transform -1 0 1284 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_199
timestamp 1625156677
transform 1 0 1284 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_314
timestamp 1625156677
transform -1 0 1340 0 -1 1505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_155
timestamp 1625156677
transform -1 0 1396 0 -1 1505
box -2 -3 58 103
use FILL  FILL_14_2_0
timestamp 1625156677
transform 1 0 1396 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1625156677
transform 1 0 1404 0 -1 1505
box -2 -3 10 103
use XOR2X1  XOR2X1_302
timestamp 1625156677
transform 1 0 1412 0 -1 1505
box -2 -3 58 103
use OAI21X1  OAI21X1_593
timestamp 1625156677
transform 1 0 1468 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_354
timestamp 1625156677
transform 1 0 1500 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_265
timestamp 1625156677
transform 1 0 1532 0 -1 1505
box -2 -3 98 103
use XNOR2X1  XNOR2X1_154
timestamp 1625156677
transform -1 0 1684 0 -1 1505
box -2 -3 58 103
use NOR2X1  NOR2X1_201
timestamp 1625156677
transform 1 0 1684 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_367
timestamp 1625156677
transform -1 0 1740 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_606
timestamp 1625156677
transform 1 0 1740 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_660
timestamp 1625156677
transform 1 0 1772 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_434
timestamp 1625156677
transform -1 0 1820 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_679
timestamp 1625156677
transform 1 0 1820 0 -1 1505
box -2 -3 26 103
use OR2X2  OR2X2_144
timestamp 1625156677
transform -1 0 1876 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_3_0
timestamp 1625156677
transform 1 0 1876 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1625156677
transform 1 0 1884 0 -1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_430
timestamp 1625156677
transform 1 0 1892 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_622
timestamp 1625156677
transform -1 0 1948 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_187
timestamp 1625156677
transform -1 0 1980 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_644
timestamp 1625156677
transform -1 0 2004 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_366
timestamp 1625156677
transform 1 0 2004 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_605
timestamp 1625156677
transform 1 0 2036 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_181
timestamp 1625156677
transform -1 0 2100 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_384
timestamp 1625156677
transform -1 0 2132 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_671
timestamp 1625156677
transform -1 0 2156 0 -1 1505
box -2 -3 26 103
use OR2X2  OR2X2_140
timestamp 1625156677
transform -1 0 2188 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_249
timestamp 1625156677
transform 1 0 2188 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_688
timestamp 1625156677
transform 1 0 2284 0 -1 1505
box -2 -3 26 103
use XOR2X1  XOR2X1_161
timestamp 1625156677
transform -1 0 2364 0 -1 1505
box -2 -3 58 103
use XOR2X1  XOR2X1_159
timestamp 1625156677
transform -1 0 2420 0 -1 1505
box -2 -3 58 103
use FILL  FILL_14_4_0
timestamp 1625156677
transform -1 0 2428 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_4_1
timestamp 1625156677
transform -1 0 2436 0 -1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_304
timestamp 1625156677
transform -1 0 2460 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_362
timestamp 1625156677
transform 1 0 2460 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_601
timestamp 1625156677
transform 1 0 2492 0 -1 1505
box -2 -3 34 103
use XOR2X1  XOR2X1_134
timestamp 1625156677
transform -1 0 2580 0 -1 1505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_138
timestamp 1625156677
transform 1 0 2580 0 -1 1505
box -2 -3 58 103
use NAND3X1  NAND3X1_274
timestamp 1625156677
transform -1 0 2668 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_175
timestamp 1625156677
transform 1 0 2668 0 -1 1505
box -2 -3 18 103
use OR2X2  OR2X2_119
timestamp 1625156677
transform -1 0 2716 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_300
timestamp 1625156677
transform -1 0 2740 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_299
timestamp 1625156677
transform -1 0 2764 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_171
timestamp 1625156677
transform -1 0 2780 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_240
timestamp 1625156677
transform -1 0 2876 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_5_0
timestamp 1625156677
transform -1 0 2884 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_5_1
timestamp 1625156677
transform -1 0 2892 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_241
timestamp 1625156677
transform -1 0 2988 0 -1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_330
timestamp 1625156677
transform 1 0 2988 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_575
timestamp 1625156677
transform 1 0 3020 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1625156677
transform 1 0 3052 0 -1 1505
box -2 -3 98 103
use BUFX4  BUFX4_31
timestamp 1625156677
transform -1 0 3180 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_389
timestamp 1625156677
transform 1 0 3180 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_574
timestamp 1625156677
transform 1 0 3204 0 -1 1505
box -2 -3 34 103
use INVX2  INVX2_82
timestamp 1625156677
transform 1 0 3236 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1625156677
transform 1 0 3252 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_369
timestamp 1625156677
transform 1 0 3348 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_493
timestamp 1625156677
transform -1 0 3404 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_390
timestamp 1625156677
transform -1 0 3428 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_6_0
timestamp 1625156677
transform 1 0 3428 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_6_1
timestamp 1625156677
transform 1 0 3436 0 -1 1505
box -2 -3 10 103
use INVX1  INVX1_488
timestamp 1625156677
transform 1 0 3444 0 -1 1505
box -2 -3 18 103
use NAND3X1  NAND3X1_492
timestamp 1625156677
transform -1 0 3492 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_331
timestamp 1625156677
transform 1 0 3492 0 -1 1505
box -2 -3 34 103
use NOR3X1  NOR3X1_87
timestamp 1625156677
transform 1 0 3524 0 -1 1505
box -2 -3 66 103
use INVX1  INVX1_477
timestamp 1625156677
transform 1 0 3588 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_393
timestamp 1625156677
transform 1 0 3604 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_370
timestamp 1625156677
transform 1 0 3628 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_29
timestamp 1625156677
transform 1 0 3652 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_32
timestamp 1625156677
transform 1 0 3684 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_619
timestamp 1625156677
transform -1 0 3740 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_16
timestamp 1625156677
transform -1 0 3772 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_364
timestamp 1625156677
transform -1 0 3796 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1625156677
transform 1 0 3796 0 -1 1505
box -2 -3 98 103
use BUFX2  BUFX2_269
timestamp 1625156677
transform 1 0 3892 0 -1 1505
box -2 -3 26 103
use BUFX2  BUFX2_94
timestamp 1625156677
transform 1 0 3916 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_7_0
timestamp 1625156677
transform 1 0 3940 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_7_1
timestamp 1625156677
transform 1 0 3948 0 -1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_374
timestamp 1625156677
transform 1 0 3956 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1625156677
transform 1 0 3980 0 -1 1505
box -2 -3 98 103
use INVX2  INVX2_79
timestamp 1625156677
transform -1 0 4092 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_373
timestamp 1625156677
transform 1 0 4092 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_499
timestamp 1625156677
transform -1 0 4148 0 -1 1505
box -2 -3 34 103
use INVX2  INVX2_78
timestamp 1625156677
transform -1 0 4164 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_217
timestamp 1625156677
transform 1 0 4164 0 -1 1505
box -2 -3 98 103
use AND2X2  AND2X2_167
timestamp 1625156677
transform 1 0 4260 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_266
timestamp 1625156677
transform -1 0 4316 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_228
timestamp 1625156677
transform -1 0 4348 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_152
timestamp 1625156677
transform -1 0 4364 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_264
timestamp 1625156677
transform -1 0 4388 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_263
timestamp 1625156677
transform -1 0 4412 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_150
timestamp 1625156677
transform 1 0 4412 0 -1 1505
box -2 -3 18 103
use FILL  FILL_14_8_0
timestamp 1625156677
transform 1 0 4428 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_8_1
timestamp 1625156677
transform 1 0 4436 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_227
timestamp 1625156677
transform 1 0 4444 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_226
timestamp 1625156677
transform -1 0 4508 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_148
timestamp 1625156677
transform 1 0 4508 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_145
timestamp 1625156677
transform -1 0 4548 0 -1 1505
box -2 -3 26 103
use OR2X2  OR2X2_102
timestamp 1625156677
transform -1 0 4580 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_162
timestamp 1625156677
transform -1 0 4612 0 -1 1505
box -2 -3 34 103
use XOR2X1  XOR2X1_97
timestamp 1625156677
transform -1 0 4668 0 -1 1505
box -2 -3 58 103
use BUFX2  BUFX2_157
timestamp 1625156677
transform 1 0 4668 0 -1 1505
box -2 -3 26 103
use XOR2X1  XOR2X1_118
timestamp 1625156677
transform -1 0 4748 0 -1 1505
box -2 -3 58 103
use NOR2X1  NOR2X1_127
timestamp 1625156677
transform 1 0 4748 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_194
timestamp 1625156677
transform 1 0 4772 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_130
timestamp 1625156677
transform -1 0 4820 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_228
timestamp 1625156677
transform -1 0 4844 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_226
timestamp 1625156677
transform -1 0 4868 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_225
timestamp 1625156677
transform -1 0 4892 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_139
timestamp 1625156677
transform -1 0 4924 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_128
timestamp 1625156677
transform 1 0 4924 0 -1 1505
box -2 -3 18 103
use FILL  FILL_14_9_0
timestamp 1625156677
transform -1 0 4948 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_9_1
timestamp 1625156677
transform -1 0 4956 0 -1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_200
timestamp 1625156677
transform -1 0 4988 0 -1 1505
box -2 -3 34 103
use INVX2  INVX2_42
timestamp 1625156677
transform -1 0 5004 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_218
timestamp 1625156677
transform -1 0 5028 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_140
timestamp 1625156677
transform 1 0 5028 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_142
timestamp 1625156677
transform 1 0 5060 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_67
timestamp 1625156677
transform 1 0 5092 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_124
timestamp 1625156677
transform -1 0 5148 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_189
timestamp 1625156677
transform 1 0 5148 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_190
timestamp 1625156677
transform 1 0 5180 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_207
timestamp 1625156677
transform -1 0 5308 0 -1 1505
box -2 -3 98 103
use FILL  FILL_15_1
timestamp 1625156677
transform -1 0 5316 0 -1 1505
box -2 -3 10 103
use NAND3X1  NAND3X1_321
timestamp 1625156677
transform -1 0 36 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_230
timestamp 1625156677
transform 1 0 36 0 1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_322
timestamp 1625156677
transform -1 0 84 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_221
timestamp 1625156677
transform -1 0 116 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_209
timestamp 1625156677
transform 1 0 116 0 1 1305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_157
timestamp 1625156677
transform 1 0 140 0 1 1305
box -2 -3 58 103
use NOR2X1  NOR2X1_208
timestamp 1625156677
transform -1 0 220 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_224
timestamp 1625156677
transform 1 0 220 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_374
timestamp 1625156677
transform -1 0 276 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_335
timestamp 1625156677
transform 1 0 276 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_372
timestamp 1625156677
transform -1 0 332 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_0_0
timestamp 1625156677
transform 1 0 332 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1625156677
transform 1 0 340 0 1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_225
timestamp 1625156677
transform 1 0 348 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_326
timestamp 1625156677
transform -1 0 412 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_236
timestamp 1625156677
transform 1 0 412 0 1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_327
timestamp 1625156677
transform -1 0 460 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_370
timestamp 1625156677
transform -1 0 484 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_371
timestamp 1625156677
transform -1 0 508 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_235
timestamp 1625156677
transform -1 0 524 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_330
timestamp 1625156677
transform -1 0 556 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_331
timestamp 1625156677
transform -1 0 588 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_210
timestamp 1625156677
transform 1 0 588 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_361
timestamp 1625156677
transform -1 0 636 0 1 1305
box -2 -3 26 103
use XOR2X1  XOR2X1_176
timestamp 1625156677
transform 1 0 636 0 1 1305
box -2 -3 58 103
use XOR2X1  XOR2X1_177
timestamp 1625156677
transform 1 0 692 0 1 1305
box -2 -3 58 103
use XOR2X1  XOR2X1_178
timestamp 1625156677
transform -1 0 804 0 1 1305
box -2 -3 58 103
use NAND2X1  NAND2X1_342
timestamp 1625156677
transform -1 0 828 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_305
timestamp 1625156677
transform -1 0 860 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_1_0
timestamp 1625156677
transform -1 0 868 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1625156677
transform -1 0 876 0 1 1305
box -2 -3 10 103
use INVX1  INVX1_205
timestamp 1625156677
transform -1 0 892 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_334
timestamp 1625156677
transform -1 0 916 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_209
timestamp 1625156677
transform 1 0 916 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_198
timestamp 1625156677
transform 1 0 948 0 1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_301
timestamp 1625156677
transform -1 0 996 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_300
timestamp 1625156677
transform 1 0 996 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_333
timestamp 1625156677
transform -1 0 1052 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_332
timestamp 1625156677
transform -1 0 1076 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_197
timestamp 1625156677
transform -1 0 1092 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_292
timestamp 1625156677
transform -1 0 1124 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_186
timestamp 1625156677
transform -1 0 1148 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_293
timestamp 1625156677
transform -1 0 1180 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_541
timestamp 1625156677
transform -1 0 1196 0 1 1305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_31
timestamp 1625156677
transform -1 0 1268 0 1 1305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_254
timestamp 1625156677
transform -1 0 1364 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_2_0
timestamp 1625156677
transform -1 0 1372 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1625156677
transform -1 0 1380 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_255
timestamp 1625156677
transform -1 0 1476 0 1 1305
box -2 -3 98 103
use CLKBUF1  CLKBUF1_11
timestamp 1625156677
transform 1 0 1476 0 1 1305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_256
timestamp 1625156677
transform -1 0 1644 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_264
timestamp 1625156677
transform -1 0 1740 0 1 1305
box -2 -3 98 103
use XNOR2X1  XNOR2X1_229
timestamp 1625156677
transform -1 0 1796 0 1 1305
box -2 -3 58 103
use INVX1  INVX1_529
timestamp 1625156677
transform -1 0 1812 0 1 1305
box -2 -3 18 103
use XOR2X1  XOR2X1_168
timestamp 1625156677
transform -1 0 1868 0 1 1305
box -2 -3 58 103
use FILL  FILL_13_3_0
timestamp 1625156677
transform 1 0 1868 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1625156677
transform 1 0 1876 0 1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_393
timestamp 1625156677
transform 1 0 1884 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_513
timestamp 1625156677
transform 1 0 1916 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_526
timestamp 1625156677
transform -1 0 1964 0 1 1305
box -2 -3 18 103
use XOR2X1  XOR2X1_169
timestamp 1625156677
transform -1 0 2020 0 1 1305
box -2 -3 58 103
use NAND3X1  NAND3X1_519
timestamp 1625156677
transform -1 0 2052 0 1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_233
timestamp 1625156677
transform -1 0 2108 0 1 1305
box -2 -3 58 103
use OAI21X1  OAI21X1_613
timestamp 1625156677
transform -1 0 2140 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_424
timestamp 1625156677
transform -1 0 2164 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_620
timestamp 1625156677
transform 1 0 2164 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_425
timestamp 1625156677
transform 1 0 2196 0 1 1305
box -2 -3 26 103
use INVX2  INVX2_89
timestamp 1625156677
transform -1 0 2236 0 1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_508
timestamp 1625156677
transform -1 0 2268 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_577
timestamp 1625156677
transform 1 0 2268 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_625
timestamp 1625156677
transform -1 0 2316 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_549
timestamp 1625156677
transform 1 0 2316 0 1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_515
timestamp 1625156677
transform -1 0 2364 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_575
timestamp 1625156677
transform -1 0 2380 0 1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_189
timestamp 1625156677
transform 1 0 2380 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_4_0
timestamp 1625156677
transform -1 0 2412 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_4_1
timestamp 1625156677
transform -1 0 2420 0 1 1305
box -2 -3 10 103
use XOR2X1  XOR2X1_157
timestamp 1625156677
transform -1 0 2476 0 1 1305
box -2 -3 58 103
use XOR2X1  XOR2X1_133
timestamp 1625156677
transform -1 0 2532 0 1 1305
box -2 -3 58 103
use INVX1  INVX1_519
timestamp 1625156677
transform -1 0 2548 0 1 1305
box -2 -3 18 103
use XOR2X1  XOR2X1_156
timestamp 1625156677
transform -1 0 2604 0 1 1305
box -2 -3 58 103
use XOR2X1  XOR2X1_158
timestamp 1625156677
transform -1 0 2660 0 1 1305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_135
timestamp 1625156677
transform 1 0 2660 0 1 1305
box -2 -3 58 103
use INVX2  INVX2_55
timestamp 1625156677
transform -1 0 2732 0 1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_166
timestamp 1625156677
transform -1 0 2756 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_167
timestamp 1625156677
transform -1 0 2780 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_261
timestamp 1625156677
transform 1 0 2780 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_172
timestamp 1625156677
transform -1 0 2828 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_260
timestamp 1625156677
transform 1 0 2828 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_262
timestamp 1625156677
transform -1 0 2892 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_174
timestamp 1625156677
transform -1 0 2908 0 1 1305
box -2 -3 18 103
use FILL  FILL_13_5_0
timestamp 1625156677
transform -1 0 2916 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_5_1
timestamp 1625156677
transform -1 0 2924 0 1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_302
timestamp 1625156677
transform -1 0 2948 0 1 1305
box -2 -3 26 103
use OR2X2  OR2X2_120
timestamp 1625156677
transform -1 0 2980 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_301
timestamp 1625156677
transform -1 0 3004 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_525
timestamp 1625156677
transform -1 0 3020 0 1 1305
box -2 -3 18 103
use BUFX2  BUFX2_171
timestamp 1625156677
transform 1 0 3020 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_296
timestamp 1625156677
transform 1 0 3044 0 1 1305
box -2 -3 26 103
use OR2X2  OR2X2_117
timestamp 1625156677
transform -1 0 3100 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_164
timestamp 1625156677
transform -1 0 3124 0 1 1305
box -2 -3 26 103
use AND2X2  AND2X2_91
timestamp 1625156677
transform -1 0 3156 0 1 1305
box -2 -3 34 103
use BUFX2  BUFX2_168
timestamp 1625156677
transform -1 0 3180 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_522
timestamp 1625156677
transform -1 0 3196 0 1 1305
box -2 -3 18 103
use BUFX2  BUFX2_259
timestamp 1625156677
transform 1 0 3196 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_201
timestamp 1625156677
transform 1 0 3220 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_224
timestamp 1625156677
transform 1 0 3316 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_6_0
timestamp 1625156677
transform 1 0 3412 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_6_1
timestamp 1625156677
transform 1 0 3420 0 1 1305
box -2 -3 10 103
use INVX1  INVX1_149
timestamp 1625156677
transform 1 0 3428 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1625156677
transform 1 0 3444 0 1 1305
box -2 -3 98 103
use INVX2  INVX2_83
timestamp 1625156677
transform -1 0 3556 0 1 1305
box -2 -3 18 103
use INVX1  INVX1_480
timestamp 1625156677
transform -1 0 3572 0 1 1305
box -2 -3 18 103
use AND2X2  AND2X2_172
timestamp 1625156677
transform -1 0 3604 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_403
timestamp 1625156677
transform 1 0 3604 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_629
timestamp 1625156677
transform 1 0 3628 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1625156677
transform -1 0 3748 0 1 1305
box -2 -3 98 103
use AND2X2  AND2X2_163
timestamp 1625156677
transform -1 0 3780 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_576
timestamp 1625156677
transform 1 0 3780 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_333
timestamp 1625156677
transform -1 0 3844 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1625156677
transform -1 0 3940 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_7_0
timestamp 1625156677
transform 1 0 3940 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_7_1
timestamp 1625156677
transform 1 0 3948 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_216
timestamp 1625156677
transform 1 0 3956 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1625156677
transform 1 0 4052 0 1 1305
box -2 -3 98 103
use AND2X2  AND2X2_175
timestamp 1625156677
transform -1 0 4180 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_585
timestamp 1625156677
transform -1 0 4212 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_404
timestamp 1625156677
transform -1 0 4236 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_343
timestamp 1625156677
transform -1 0 4268 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_586
timestamp 1625156677
transform 1 0 4268 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_344
timestamp 1625156677
transform 1 0 4300 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_405
timestamp 1625156677
transform 1 0 4332 0 1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1625156677
transform -1 0 4452 0 1 1305
box -2 -3 98 103
use FILL  FILL_13_8_0
timestamp 1625156677
transform -1 0 4460 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_8_1
timestamp 1625156677
transform -1 0 4468 0 1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_238
timestamp 1625156677
transform -1 0 4500 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_153
timestamp 1625156677
transform -1 0 4516 0 1 1305
box -2 -3 18 103
use OR2X2  OR2X2_104
timestamp 1625156677
transform -1 0 4548 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_262
timestamp 1625156677
transform -1 0 4572 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_261
timestamp 1625156677
transform 1 0 4572 0 1 1305
box -2 -3 26 103
use OR2X2  OR2X2_103
timestamp 1625156677
transform 1 0 4596 0 1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_120
timestamp 1625156677
transform -1 0 4684 0 1 1305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_118
timestamp 1625156677
transform 1 0 4684 0 1 1305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_119
timestamp 1625156677
transform 1 0 4740 0 1 1305
box -2 -3 58 103
use BUFX2  BUFX2_162
timestamp 1625156677
transform 1 0 4796 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_131
timestamp 1625156677
transform -1 0 4836 0 1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_202
timestamp 1625156677
transform 1 0 4836 0 1 1305
box -2 -3 34 103
use OR2X2  OR2X2_88
timestamp 1625156677
transform -1 0 4900 0 1 1305
box -2 -3 34 103
use BUFX2  BUFX2_161
timestamp 1625156677
transform 1 0 4900 0 1 1305
box -2 -3 26 103
use XOR2X1  XOR2X1_110
timestamp 1625156677
transform 1 0 4924 0 1 1305
box -2 -3 58 103
use FILL  FILL_13_9_0
timestamp 1625156677
transform -1 0 4988 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_9_1
timestamp 1625156677
transform -1 0 4996 0 1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_201
timestamp 1625156677
transform -1 0 5028 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_121
timestamp 1625156677
transform -1 0 5052 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_129
timestamp 1625156677
transform -1 0 5068 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_182
timestamp 1625156677
transform -1 0 5100 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_187
timestamp 1625156677
transform 1 0 5100 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_135
timestamp 1625156677
transform -1 0 5164 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_220
timestamp 1625156677
transform 1 0 5164 0 1 1305
box -2 -3 26 103
use OR2X2  OR2X2_85
timestamp 1625156677
transform 1 0 5188 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_125
timestamp 1625156677
transform -1 0 5236 0 1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_198
timestamp 1625156677
transform 1 0 5236 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_196
timestamp 1625156677
transform 1 0 5268 0 1 1305
box -2 -3 34 103
use FILL  FILL_14_1
timestamp 1625156677
transform 1 0 5300 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_2
timestamp 1625156677
transform 1 0 5308 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_324
timestamp 1625156677
transform 1 0 4 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_367
timestamp 1625156677
transform -1 0 60 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_368
timestamp 1625156677
transform -1 0 84 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_229
timestamp 1625156677
transform -1 0 100 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_325
timestamp 1625156677
transform 1 0 100 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_329
timestamp 1625156677
transform 1 0 132 0 -1 1305
box -2 -3 34 103
use XOR2X1  XOR2X1_188
timestamp 1625156677
transform 1 0 164 0 -1 1305
box -2 -3 58 103
use AOI21X1  AOI21X1_219
timestamp 1625156677
transform -1 0 252 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_325
timestamp 1625156677
transform 1 0 252 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_231
timestamp 1625156677
transform -1 0 300 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_220
timestamp 1625156677
transform -1 0 332 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_0_0
timestamp 1625156677
transform 1 0 332 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1625156677
transform 1 0 340 0 -1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_329
timestamp 1625156677
transform 1 0 348 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_379
timestamp 1625156677
transform 1 0 380 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_334
timestamp 1625156677
transform -1 0 436 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_242
timestamp 1625156677
transform -1 0 452 0 -1 1305
box -2 -3 18 103
use AND2X2  AND2X2_109
timestamp 1625156677
transform 1 0 452 0 -1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_10
timestamp 1625156677
transform -1 0 524 0 -1 1305
box -2 -3 42 103
use INVX1  INVX1_238
timestamp 1625156677
transform 1 0 524 0 -1 1305
box -2 -3 18 103
use XOR2X1  XOR2X1_187
timestamp 1625156677
transform -1 0 596 0 -1 1305
box -2 -3 58 103
use BUFX2  BUFX2_179
timestamp 1625156677
transform -1 0 620 0 -1 1305
box -2 -3 26 103
use XOR2X1  XOR2X1_170
timestamp 1625156677
transform -1 0 676 0 -1 1305
box -2 -3 58 103
use AND2X2  AND2X2_101
timestamp 1625156677
transform -1 0 708 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_304
timestamp 1625156677
transform -1 0 740 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_210
timestamp 1625156677
transform 1 0 740 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_204
timestamp 1625156677
transform -1 0 788 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_296
timestamp 1625156677
transform 1 0 788 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_203
timestamp 1625156677
transform -1 0 836 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_298
timestamp 1625156677
transform 1 0 836 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_1_0
timestamp 1625156677
transform 1 0 868 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1625156677
transform 1 0 876 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_202
timestamp 1625156677
transform 1 0 884 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_340
timestamp 1625156677
transform -1 0 924 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_339
timestamp 1625156677
transform -1 0 948 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_188
timestamp 1625156677
transform 1 0 948 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_200
timestamp 1625156677
transform -1 0 988 0 -1 1305
box -2 -3 18 103
use AOI22X1  AOI22X1_8
timestamp 1625156677
transform -1 0 1028 0 -1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_341
timestamp 1625156677
transform -1 0 1052 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_303
timestamp 1625156677
transform 1 0 1052 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_194
timestamp 1625156677
transform 1 0 1084 0 -1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_298
timestamp 1625156677
transform -1 0 1132 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_297
timestamp 1625156677
transform 1 0 1132 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_196
timestamp 1625156677
transform -1 0 1180 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_289
timestamp 1625156677
transform -1 0 1212 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_195
timestamp 1625156677
transform -1 0 1228 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_288
timestamp 1625156677
transform -1 0 1260 0 -1 1305
box -2 -3 34 103
use BUFX2  BUFX2_54
timestamp 1625156677
transform -1 0 1284 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_592
timestamp 1625156677
transform 1 0 1284 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_353
timestamp 1625156677
transform 1 0 1316 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_496
timestamp 1625156677
transform -1 0 1364 0 -1 1305
box -2 -3 18 103
use FILL  FILL_12_2_0
timestamp 1625156677
transform -1 0 1372 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1625156677
transform -1 0 1380 0 -1 1305
box -2 -3 10 103
use BUFX2  BUFX2_176
timestamp 1625156677
transform -1 0 1404 0 -1 1305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_151
timestamp 1625156677
transform 1 0 1404 0 -1 1305
box -2 -3 58 103
use NAND2X1  NAND2X1_338
timestamp 1625156677
transform 1 0 1460 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_1
timestamp 1625156677
transform -1 0 1516 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_337
timestamp 1625156677
transform 1 0 1516 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_201
timestamp 1625156677
transform -1 0 1556 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_295
timestamp 1625156677
transform -1 0 1588 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_187
timestamp 1625156677
transform 1 0 1588 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_594
timestamp 1625156677
transform 1 0 1612 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_355
timestamp 1625156677
transform 1 0 1644 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_498
timestamp 1625156677
transform -1 0 1692 0 -1 1305
box -2 -3 18 103
use AND2X2  AND2X2_186
timestamp 1625156677
transform 1 0 1692 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_365
timestamp 1625156677
transform -1 0 1756 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_604
timestamp 1625156677
transform -1 0 1788 0 -1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_150
timestamp 1625156677
transform 1 0 1788 0 -1 1305
box -2 -3 58 103
use AOI21X1  AOI21X1_385
timestamp 1625156677
transform -1 0 1876 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_3_0
timestamp 1625156677
transform 1 0 1876 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1625156677
transform 1 0 1884 0 -1 1305
box -2 -3 10 103
use AND2X2  AND2X2_182
timestamp 1625156677
transform 1 0 1892 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_528
timestamp 1625156677
transform -1 0 1940 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_257
timestamp 1625156677
transform -1 0 2036 0 -1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_596
timestamp 1625156677
transform -1 0 2068 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_357
timestamp 1625156677
transform 1 0 2068 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_500
timestamp 1625156677
transform -1 0 2116 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_377
timestamp 1625156677
transform -1 0 2148 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_542
timestamp 1625156677
transform -1 0 2164 0 -1 1305
box -2 -3 18 103
use INVX1  INVX1_548
timestamp 1625156677
transform -1 0 2180 0 -1 1305
box -2 -3 18 103
use INVX2  INVX2_87
timestamp 1625156677
transform -1 0 2196 0 -1 1305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_232
timestamp 1625156677
transform 1 0 2196 0 -1 1305
box -2 -3 58 103
use BUFX2  BUFX2_177
timestamp 1625156677
transform 1 0 2252 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_368
timestamp 1625156677
transform 1 0 2276 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_607
timestamp 1625156677
transform 1 0 2308 0 -1 1305
box -2 -3 34 103
use BUFX2  BUFX2_178
timestamp 1625156677
transform 1 0 2340 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_4_0
timestamp 1625156677
transform 1 0 2364 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_4_1
timestamp 1625156677
transform 1 0 2372 0 -1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_208
timestamp 1625156677
transform 1 0 2380 0 -1 1305
box -2 -3 98 103
use INVX2  INVX2_53
timestamp 1625156677
transform -1 0 2492 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_234
timestamp 1625156677
transform -1 0 2588 0 -1 1305
box -2 -3 98 103
use BUFX2  BUFX2_31
timestamp 1625156677
transform 1 0 2588 0 -1 1305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_134
timestamp 1625156677
transform 1 0 2612 0 -1 1305
box -2 -3 58 103
use AOI21X1  AOI21X1_190
timestamp 1625156677
transform 1 0 2668 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_303
timestamp 1625156677
transform -1 0 2724 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_259
timestamp 1625156677
transform 1 0 2724 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_297
timestamp 1625156677
transform -1 0 2780 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_187
timestamp 1625156677
transform 1 0 2780 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_165
timestamp 1625156677
transform 1 0 2812 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_170
timestamp 1625156677
transform -1 0 2852 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_186
timestamp 1625156677
transform -1 0 2884 0 -1 1305
box -2 -3 34 103
use OR2X2  OR2X2_118
timestamp 1625156677
transform -1 0 2916 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_5_0
timestamp 1625156677
transform -1 0 2924 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_5_1
timestamp 1625156677
transform -1 0 2932 0 -1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_271
timestamp 1625156677
transform -1 0 2964 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_298
timestamp 1625156677
transform -1 0 2988 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_269
timestamp 1625156677
transform 1 0 2988 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_270
timestamp 1625156677
transform -1 0 3052 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_268
timestamp 1625156677
transform -1 0 3084 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_169
timestamp 1625156677
transform -1 0 3100 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_258
timestamp 1625156677
transform -1 0 3132 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_257
timestamp 1625156677
transform 1 0 3132 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_239
timestamp 1625156677
transform -1 0 3260 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1625156677
transform -1 0 3356 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1625156677
transform -1 0 3452 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_6_0
timestamp 1625156677
transform 1 0 3452 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_6_1
timestamp 1625156677
transform 1 0 3460 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_489
timestamp 1625156677
transform 1 0 3468 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_394
timestamp 1625156677
transform 1 0 3484 0 -1 1305
box -2 -3 26 103
use BUFX2  BUFX2_270
timestamp 1625156677
transform -1 0 3532 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_580
timestamp 1625156677
transform -1 0 3564 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_338
timestamp 1625156677
transform -1 0 3596 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_628
timestamp 1625156677
transform 1 0 3596 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_14
timestamp 1625156677
transform 1 0 3620 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_339
timestamp 1625156677
transform 1 0 3652 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_581
timestamp 1625156677
transform 1 0 3684 0 -1 1305
box -2 -3 34 103
use INVX2  INVX2_77
timestamp 1625156677
transform -1 0 3732 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1625156677
transform -1 0 3828 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1625156677
transform -1 0 3924 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_7_0
timestamp 1625156677
transform -1 0 3932 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_7_1
timestamp 1625156677
transform -1 0 3940 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_377
timestamp 1625156677
transform -1 0 3964 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1625156677
transform -1 0 4060 0 -1 1305
box -2 -3 98 103
use BUFX4  BUFX4_15
timestamp 1625156677
transform 1 0 4060 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_376
timestamp 1625156677
transform 1 0 4092 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_484
timestamp 1625156677
transform -1 0 4132 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1625156677
transform -1 0 4228 0 -1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_375
timestamp 1625156677
transform 1 0 4228 0 -1 1305
box -2 -3 26 103
use NOR3X1  NOR3X1_92
timestamp 1625156677
transform 1 0 4252 0 -1 1305
box -2 -3 66 103
use OAI21X1  OAI21X1_584
timestamp 1625156677
transform -1 0 4348 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_342
timestamp 1625156677
transform -1 0 4380 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1625156677
transform -1 0 4476 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_8_0
timestamp 1625156677
transform -1 0 4484 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_8_1
timestamp 1625156677
transform -1 0 4492 0 -1 1305
box -2 -3 10 103
use XOR2X1  XOR2X1_98
timestamp 1625156677
transform -1 0 4548 0 -1 1305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_225
timestamp 1625156677
transform 1 0 4548 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_127
timestamp 1625156677
transform 1 0 4644 0 -1 1305
box -2 -3 18 103
use XOR2X1  XOR2X1_131
timestamp 1625156677
transform -1 0 4716 0 -1 1305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_100
timestamp 1625156677
transform -1 0 4772 0 -1 1305
box -2 -3 58 103
use NAND2X1  NAND2X1_223
timestamp 1625156677
transform 1 0 4772 0 -1 1305
box -2 -3 26 103
use OR2X2  OR2X2_87
timestamp 1625156677
transform 1 0 4796 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_224
timestamp 1625156677
transform 1 0 4828 0 -1 1305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_102
timestamp 1625156677
transform -1 0 4908 0 -1 1305
box -2 -3 58 103
use CLKBUF1  CLKBUF1_50
timestamp 1625156677
transform -1 0 4980 0 -1 1305
box -2 -3 74 103
use FILL  FILL_12_9_0
timestamp 1625156677
transform -1 0 4988 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_9_1
timestamp 1625156677
transform -1 0 4996 0 -1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_212
timestamp 1625156677
transform -1 0 5020 0 -1 1305
box -2 -3 26 103
use BUFX2  BUFX2_273
timestamp 1625156677
transform 1 0 5020 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_186
timestamp 1625156677
transform -1 0 5076 0 -1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_97
timestamp 1625156677
transform -1 0 5132 0 -1 1305
box -2 -3 58 103
use NAND2X1  NAND2X1_215
timestamp 1625156677
transform 1 0 5132 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_123
timestamp 1625156677
transform 1 0 5156 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_181
timestamp 1625156677
transform -1 0 5212 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_189
timestamp 1625156677
transform 1 0 5212 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_179
timestamp 1625156677
transform -1 0 5276 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_214
timestamp 1625156677
transform -1 0 5300 0 -1 1305
box -2 -3 26 103
use FILL  FILL_13_1
timestamp 1625156677
transform -1 0 5308 0 -1 1305
box -2 -3 10 103
use FILL  FILL_13_2
timestamp 1625156677
transform -1 0 5316 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_207
timestamp 1625156677
transform 1 0 4 0 1 1105
box -2 -3 26 103
use XOR2X1  XOR2X1_174
timestamp 1625156677
transform -1 0 84 0 1 1105
box -2 -3 58 103
use INVX1  INVX1_232
timestamp 1625156677
transform 1 0 84 0 1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_324
timestamp 1625156677
transform -1 0 132 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_323
timestamp 1625156677
transform 1 0 132 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_233
timestamp 1625156677
transform -1 0 180 0 1 1105
box -2 -3 18 103
use INVX1  INVX1_234
timestamp 1625156677
transform -1 0 196 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_327
timestamp 1625156677
transform -1 0 228 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_326
timestamp 1625156677
transform 1 0 228 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_226
timestamp 1625156677
transform -1 0 292 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_330
timestamp 1625156677
transform -1 0 324 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_241
timestamp 1625156677
transform 1 0 324 0 1 1105
box -2 -3 18 103
use FILL  FILL_11_0_0
timestamp 1625156677
transform 1 0 340 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1625156677
transform 1 0 348 0 1 1105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_158
timestamp 1625156677
transform 1 0 356 0 1 1105
box -2 -3 58 103
use NOR2X1  NOR2X1_213
timestamp 1625156677
transform -1 0 436 0 1 1105
box -2 -3 26 103
use XOR2X1  XOR2X1_175
timestamp 1625156677
transform 1 0 436 0 1 1105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_149
timestamp 1625156677
transform 1 0 492 0 1 1105
box -2 -3 58 103
use NAND2X1  NAND2X1_336
timestamp 1625156677
transform -1 0 572 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_185
timestamp 1625156677
transform -1 0 596 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_297
timestamp 1625156677
transform 1 0 596 0 1 1105
box -2 -3 34 103
use AND2X2  AND2X2_99
timestamp 1625156677
transform -1 0 660 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_326
timestamp 1625156677
transform -1 0 684 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_188
timestamp 1625156677
transform -1 0 700 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_291
timestamp 1625156677
transform 1 0 700 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_184
timestamp 1625156677
transform -1 0 756 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_193
timestamp 1625156677
transform 1 0 756 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_203
timestamp 1625156677
transform -1 0 804 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_299
timestamp 1625156677
transform -1 0 836 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_1_0
timestamp 1625156677
transform -1 0 844 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1625156677
transform -1 0 852 0 1 1105
box -2 -3 10 103
use XOR2X1  XOR2X1_153
timestamp 1625156677
transform -1 0 908 0 1 1105
box -2 -3 58 103
use XOR2X1  XOR2X1_152
timestamp 1625156677
transform -1 0 964 0 1 1105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_253
timestamp 1625156677
transform -1 0 1060 0 1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_204
timestamp 1625156677
transform -1 0 1092 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_121
timestamp 1625156677
transform -1 0 1116 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_70
timestamp 1625156677
transform 1 0 1116 0 1 1105
box -2 -3 26 103
use AND2X2  AND2X2_34
timestamp 1625156677
transform -1 0 1172 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_165
timestamp 1625156677
transform -1 0 1268 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_273
timestamp 1625156677
transform -1 0 1364 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_2_0
timestamp 1625156677
transform -1 0 1372 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1625156677
transform -1 0 1380 0 1 1105
box -2 -3 10 103
use INVX1  INVX1_74
timestamp 1625156677
transform -1 0 1396 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_102
timestamp 1625156677
transform -1 0 1428 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_97
timestamp 1625156677
transform 1 0 1428 0 1 1105
box -2 -3 34 103
use XOR2X1  XOR2X1_60
timestamp 1625156677
transform -1 0 1516 0 1 1105
box -2 -3 58 103
use XOR2X1  XOR2X1_155
timestamp 1625156677
transform -1 0 1572 0 1 1105
box -2 -3 58 103
use OR2X2  OR2X2_42
timestamp 1625156677
transform 1 0 1572 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_97
timestamp 1625156677
transform -1 0 1636 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_71
timestamp 1625156677
transform 1 0 1636 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_118
timestamp 1625156677
transform -1 0 1692 0 1 1105
box -2 -3 26 103
use AND2X2  AND2X2_33
timestamp 1625156677
transform -1 0 1724 0 1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_217
timestamp 1625156677
transform 1 0 1724 0 1 1105
box -2 -3 58 103
use INVX1  INVX1_516
timestamp 1625156677
transform -1 0 1796 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_656
timestamp 1625156677
transform -1 0 1820 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_509
timestamp 1625156677
transform -1 0 1852 0 1 1105
box -2 -3 34 103
use OR2X2  OR2X2_141
timestamp 1625156677
transform -1 0 1884 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_3_0
timestamp 1625156677
transform -1 0 1892 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1625156677
transform -1 0 1900 0 1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_672
timestamp 1625156677
transform -1 0 1924 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_608
timestamp 1625156677
transform -1 0 1956 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_369
timestamp 1625156677
transform -1 0 1988 0 1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_225
timestamp 1625156677
transform -1 0 2044 0 1 1105
box -2 -3 58 103
use OAI21X1  OAI21X1_621
timestamp 1625156677
transform 1 0 2044 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_378
timestamp 1625156677
transform -1 0 2108 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_547
timestamp 1625156677
transform -1 0 2124 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_599
timestamp 1625156677
transform 1 0 2124 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_360
timestamp 1625156677
transform -1 0 2188 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_158
timestamp 1625156677
transform 1 0 2188 0 1 1105
box -2 -3 26 103
use AND2X2  AND2X2_86
timestamp 1625156677
transform -1 0 2244 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_287
timestamp 1625156677
transform 1 0 2244 0 1 1105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_131
timestamp 1625156677
transform 1 0 2268 0 1 1105
box -2 -3 58 103
use NAND2X1  NAND2X1_286
timestamp 1625156677
transform 1 0 2324 0 1 1105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_132
timestamp 1625156677
transform -1 0 2404 0 1 1105
box -2 -3 58 103
use FILL  FILL_11_4_0
timestamp 1625156677
transform -1 0 2412 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_4_1
timestamp 1625156677
transform -1 0 2420 0 1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_189
timestamp 1625156677
transform -1 0 2452 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_506
timestamp 1625156677
transform 1 0 2452 0 1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_273
timestamp 1625156677
transform 1 0 2468 0 1 1105
box -2 -3 34 103
use XOR2X1  XOR2X1_150
timestamp 1625156677
transform -1 0 2556 0 1 1105
box -2 -3 58 103
use OAI21X1  OAI21X1_250
timestamp 1625156677
transform -1 0 2588 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_255
timestamp 1625156677
transform 1 0 2588 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_173
timestamp 1625156677
transform 1 0 2620 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_188
timestamp 1625156677
transform -1 0 2668 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_294
timestamp 1625156677
transform 1 0 2668 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_256
timestamp 1625156677
transform -1 0 2724 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_272
timestamp 1625156677
transform 1 0 2724 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_185
timestamp 1625156677
transform -1 0 2788 0 1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_130
timestamp 1625156677
transform 1 0 2788 0 1 1105
box -2 -3 58 103
use XOR2X1  XOR2X1_132
timestamp 1625156677
transform -1 0 2900 0 1 1105
box -2 -3 58 103
use FILL  FILL_11_5_0
timestamp 1625156677
transform -1 0 2908 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_5_1
timestamp 1625156677
transform -1 0 2916 0 1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_184
timestamp 1625156677
transform -1 0 2948 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_293
timestamp 1625156677
transform -1 0 2972 0 1 1105
box -2 -3 26 103
use OR2X2  OR2X2_116
timestamp 1625156677
transform -1 0 3004 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1625156677
transform -1 0 3100 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1625156677
transform -1 0 3196 0 1 1105
box -2 -3 98 103
use BUFX4  BUFX4_6
timestamp 1625156677
transform 1 0 3196 0 1 1105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_9
timestamp 1625156677
transform 1 0 3228 0 1 1105
box -2 -3 74 103
use BUFX4  BUFX4_28
timestamp 1625156677
transform -1 0 3332 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1625156677
transform -1 0 3428 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_6_0
timestamp 1625156677
transform -1 0 3436 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_6_1
timestamp 1625156677
transform -1 0 3444 0 1 1105
box -2 -3 10 103
use AND2X2  AND2X2_164
timestamp 1625156677
transform -1 0 3476 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_623
timestamp 1625156677
transform 1 0 3476 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_398
timestamp 1625156677
transform 1 0 3500 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_622
timestamp 1625156677
transform -1 0 3548 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_332
timestamp 1625156677
transform 1 0 3548 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_620
timestamp 1625156677
transform 1 0 3580 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_395
timestamp 1625156677
transform -1 0 3628 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1625156677
transform -1 0 3724 0 1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_396
timestamp 1625156677
transform 1 0 3724 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_621
timestamp 1625156677
transform -1 0 3772 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_397
timestamp 1625156677
transform -1 0 3796 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_478
timestamp 1625156677
transform 1 0 3796 0 1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_365
timestamp 1625156677
transform -1 0 3836 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1625156677
transform 1 0 3836 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_7_0
timestamp 1625156677
transform 1 0 3932 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_7_1
timestamp 1625156677
transform 1 0 3940 0 1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_347
timestamp 1625156677
transform 1 0 3948 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_80
timestamp 1625156677
transform -1 0 3996 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_587
timestamp 1625156677
transform 1 0 3996 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_635
timestamp 1625156677
transform 1 0 4028 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_7
timestamp 1625156677
transform 1 0 4052 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_167
timestamp 1625156677
transform -1 0 4108 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_17
timestamp 1625156677
transform 1 0 4108 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_406
timestamp 1625156677
transform -1 0 4164 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_634
timestamp 1625156677
transform -1 0 4188 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_346
timestamp 1625156677
transform -1 0 4220 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_500
timestamp 1625156677
transform 1 0 4220 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_483
timestamp 1625156677
transform -1 0 4268 0 1 1105
box -2 -3 18 103
use INVX1  INVX1_492
timestamp 1625156677
transform -1 0 4284 0 1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_345
timestamp 1625156677
transform 1 0 4284 0 1 1105
box -2 -3 34 103
use NOR3X1  NOR3X1_93
timestamp 1625156677
transform 1 0 4316 0 1 1105
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1625156677
transform -1 0 4476 0 1 1105
box -2 -3 98 103
use FILL  FILL_11_8_0
timestamp 1625156677
transform -1 0 4484 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_8_1
timestamp 1625156677
transform -1 0 4492 0 1 1105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_6
timestamp 1625156677
transform -1 0 4564 0 1 1105
box -2 -3 74 103
use XOR2X1  XOR2X1_99
timestamp 1625156677
transform 1 0 4564 0 1 1105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_190
timestamp 1625156677
transform -1 0 4716 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_203
timestamp 1625156677
transform 1 0 4716 0 1 1105
box -2 -3 98 103
use XNOR2X1  XNOR2X1_101
timestamp 1625156677
transform -1 0 4868 0 1 1105
box -2 -3 58 103
use NAND3X1  NAND3X1_185
timestamp 1625156677
transform -1 0 4900 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_121
timestamp 1625156677
transform 1 0 4900 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_178
timestamp 1625156677
transform -1 0 4948 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_9_0
timestamp 1625156677
transform 1 0 4948 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_9_1
timestamp 1625156677
transform 1 0 4956 0 1 1105
box -2 -3 10 103
use NOR3X1  NOR3X1_45
timestamp 1625156677
transform 1 0 4964 0 1 1105
box -2 -3 66 103
use XOR2X1  XOR2X1_94
timestamp 1625156677
transform 1 0 5028 0 1 1105
box -2 -3 58 103
use NAND3X1  NAND3X1_187
timestamp 1625156677
transform -1 0 5116 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_131
timestamp 1625156677
transform 1 0 5116 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_122
timestamp 1625156677
transform 1 0 5148 0 1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_119
timestamp 1625156677
transform -1 0 5188 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_180
timestamp 1625156677
transform -1 0 5220 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_60
timestamp 1625156677
transform -1 0 5244 0 1 1105
box -2 -3 26 103
use OR2X2  OR2X2_82
timestamp 1625156677
transform -1 0 5276 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_138
timestamp 1625156677
transform -1 0 5300 0 1 1105
box -2 -3 26 103
use FILL  FILL_12_1
timestamp 1625156677
transform 1 0 5300 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1625156677
transform 1 0 5308 0 1 1105
box -2 -3 10 103
use BUFX2  BUFX2_48
timestamp 1625156677
transform 1 0 4 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_243
timestamp 1625156677
transform 1 0 28 0 -1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_331
timestamp 1625156677
transform -1 0 76 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_380
timestamp 1625156677
transform -1 0 100 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_336
timestamp 1625156677
transform -1 0 132 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_240
timestamp 1625156677
transform -1 0 148 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_212
timestamp 1625156677
transform -1 0 172 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_378
timestamp 1625156677
transform -1 0 196 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_377
timestamp 1625156677
transform -1 0 220 0 -1 1105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_159
timestamp 1625156677
transform -1 0 276 0 -1 1105
box -2 -3 58 103
use BUFX2  BUFX2_183
timestamp 1625156677
transform 1 0 276 0 -1 1105
box -2 -3 26 103
use BUFX2  BUFX2_185
timestamp 1625156677
transform 1 0 300 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_0_0
timestamp 1625156677
transform -1 0 332 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1625156677
transform -1 0 340 0 -1 1105
box -2 -3 10 103
use NOR3X1  NOR3X1_58
timestamp 1625156677
transform -1 0 404 0 -1 1105
box -2 -3 66 103
use OAI21X1  OAI21X1_282
timestamp 1625156677
transform 1 0 404 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_100
timestamp 1625156677
transform 1 0 436 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_285
timestamp 1625156677
transform 1 0 468 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_208
timestamp 1625156677
transform 1 0 500 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_293
timestamp 1625156677
transform 1 0 532 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_325
timestamp 1625156677
transform -1 0 588 0 -1 1105
box -2 -3 26 103
use AND2X2  AND2X2_98
timestamp 1625156677
transform -1 0 620 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_324
timestamp 1625156677
transform -1 0 644 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_179
timestamp 1625156677
transform 1 0 644 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_281
timestamp 1625156677
transform 1 0 668 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_187
timestamp 1625156677
transform -1 0 716 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_178
timestamp 1625156677
transform 1 0 716 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_280
timestamp 1625156677
transform -1 0 772 0 -1 1105
box -2 -3 34 103
use XOR2X1  XOR2X1_154
timestamp 1625156677
transform -1 0 828 0 -1 1105
box -2 -3 58 103
use OAI21X1  OAI21X1_287
timestamp 1625156677
transform -1 0 860 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_1_0
timestamp 1625156677
transform -1 0 868 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1625156677
transform -1 0 876 0 -1 1105
box -2 -3 10 103
use XOR2X1  XOR2X1_45
timestamp 1625156677
transform -1 0 932 0 -1 1105
box -2 -3 58 103
use OR2X2  OR2X2_43
timestamp 1625156677
transform 1 0 932 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_74
timestamp 1625156677
transform 1 0 964 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_100
timestamp 1625156677
transform -1 0 1028 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_101
timestamp 1625156677
transform -1 0 1060 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_68
timestamp 1625156677
transform -1 0 1076 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_98
timestamp 1625156677
transform -1 0 1108 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_72
timestamp 1625156677
transform 1 0 1108 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_99
timestamp 1625156677
transform 1 0 1140 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_73
timestamp 1625156677
transform 1 0 1172 0 -1 1105
box -2 -3 34 103
use INVX2  INVX2_27
timestamp 1625156677
transform 1 0 1204 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_71
timestamp 1625156677
transform -1 0 1244 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_80
timestamp 1625156677
transform -1 0 1276 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_75
timestamp 1625156677
transform -1 0 1308 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_73
timestamp 1625156677
transform -1 0 1332 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_96
timestamp 1625156677
transform 1 0 1332 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_2_0
timestamp 1625156677
transform -1 0 1372 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1625156677
transform -1 0 1380 0 -1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_120
timestamp 1625156677
transform -1 0 1404 0 -1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_99
timestamp 1625156677
transform -1 0 1436 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_94
timestamp 1625156677
transform 1 0 1436 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_98
timestamp 1625156677
transform 1 0 1468 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_95
timestamp 1625156677
transform -1 0 1532 0 -1 1105
box -2 -3 34 103
use NOR3X1  NOR3X1_36
timestamp 1625156677
transform 1 0 1532 0 -1 1105
box -2 -3 66 103
use NOR2X1  NOR2X1_69
timestamp 1625156677
transform 1 0 1596 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_67
timestamp 1625156677
transform -1 0 1636 0 -1 1105
box -2 -3 18 103
use BUFX2  BUFX2_261
timestamp 1625156677
transform -1 0 1660 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_164
timestamp 1625156677
transform -1 0 1756 0 -1 1105
box -2 -3 98 103
use XNOR2X1  XNOR2X1_218
timestamp 1625156677
transform 1 0 1756 0 -1 1105
box -2 -3 58 103
use AND2X2  AND2X2_177
timestamp 1625156677
transform -1 0 1844 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_655
timestamp 1625156677
transform 1 0 1844 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_535
timestamp 1625156677
transform -1 0 1884 0 -1 1105
box -2 -3 18 103
use FILL  FILL_10_3_0
timestamp 1625156677
transform -1 0 1892 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1625156677
transform -1 0 1900 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_600
timestamp 1625156677
transform -1 0 1932 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_505
timestamp 1625156677
transform -1 0 1948 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_361
timestamp 1625156677
transform 1 0 1948 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_235
timestamp 1625156677
transform 1 0 1980 0 -1 1105
box -2 -3 98 103
use XNOR2X1  XNOR2X1_224
timestamp 1625156677
transform 1 0 2076 0 -1 1105
box -2 -3 58 103
use INVX1  INVX1_165
timestamp 1625156677
transform 1 0 2132 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_246
timestamp 1625156677
transform -1 0 2180 0 -1 1105
box -2 -3 34 103
use NOR3X1  NOR3X1_53
timestamp 1625156677
transform 1 0 2180 0 -1 1105
box -2 -3 66 103
use NAND3X1  NAND3X1_257
timestamp 1625156677
transform 1 0 2244 0 -1 1105
box -2 -3 34 103
use OR2X2  OR2X2_113
timestamp 1625156677
transform -1 0 2308 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_288
timestamp 1625156677
transform 1 0 2308 0 -1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_258
timestamp 1625156677
transform -1 0 2364 0 -1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_133
timestamp 1625156677
transform -1 0 2420 0 -1 1105
box -2 -3 58 103
use FILL  FILL_10_4_0
timestamp 1625156677
transform 1 0 2420 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_4_1
timestamp 1625156677
transform 1 0 2428 0 -1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_290
timestamp 1625156677
transform 1 0 2436 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_247
timestamp 1625156677
transform -1 0 2492 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_249
timestamp 1625156677
transform -1 0 2524 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_163
timestamp 1625156677
transform -1 0 2548 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_183
timestamp 1625156677
transform 1 0 2548 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_291
timestamp 1625156677
transform -1 0 2604 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_161
timestamp 1625156677
transform 1 0 2604 0 -1 1105
box -2 -3 26 103
use INVX2  INVX2_54
timestamp 1625156677
transform 1 0 2628 0 -1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_267
timestamp 1625156677
transform -1 0 2676 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_90
timestamp 1625156677
transform -1 0 2708 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_295
timestamp 1625156677
transform -1 0 2732 0 -1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_265
timestamp 1625156677
transform 1 0 2732 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_264
timestamp 1625156677
transform -1 0 2796 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_266
timestamp 1625156677
transform -1 0 2828 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_253
timestamp 1625156677
transform -1 0 2860 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_254
timestamp 1625156677
transform -1 0 2892 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_162
timestamp 1625156677
transform 1 0 2892 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_5_0
timestamp 1625156677
transform -1 0 2924 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_5_1
timestamp 1625156677
transform -1 0 2932 0 -1 1105
box -2 -3 10 103
use AND2X2  AND2X2_89
timestamp 1625156677
transform -1 0 2964 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1625156677
transform -1 0 3060 0 -1 1105
box -2 -3 98 103
use BUFX2  BUFX2_145
timestamp 1625156677
transform 1 0 3060 0 -1 1105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_20
timestamp 1625156677
transform -1 0 3156 0 -1 1105
box -2 -3 74 103
use OAI21X1  OAI21X1_568
timestamp 1625156677
transform 1 0 3156 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_324
timestamp 1625156677
transform -1 0 3220 0 -1 1105
box -2 -3 34 103
use INVX2  INVX2_74
timestamp 1625156677
transform -1 0 3236 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1625156677
transform 1 0 3236 0 -1 1105
box -2 -3 98 103
use AND2X2  AND2X2_160
timestamp 1625156677
transform 1 0 3332 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1625156677
transform -1 0 3460 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_6_0
timestamp 1625156677
transform -1 0 3468 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_6_1
timestamp 1625156677
transform -1 0 3476 0 -1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_399
timestamp 1625156677
transform -1 0 3500 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1625156677
transform -1 0 3596 0 -1 1105
box -2 -3 98 103
use NOR3X1  NOR3X1_88
timestamp 1625156677
transform 1 0 3596 0 -1 1105
box -2 -3 66 103
use INVX2  INVX2_84
timestamp 1625156677
transform 1 0 3660 0 -1 1105
box -2 -3 18 103
use NOR3X1  NOR3X1_90
timestamp 1625156677
transform 1 0 3676 0 -1 1105
box -2 -3 66 103
use NOR2X1  NOR2X1_371
timestamp 1625156677
transform 1 0 3740 0 -1 1105
box -2 -3 26 103
use BUFX2  BUFX2_140
timestamp 1625156677
transform 1 0 3764 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1625156677
transform 1 0 3788 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_636
timestamp 1625156677
transform 1 0 3884 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_588
timestamp 1625156677
transform 1 0 3908 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_7_0
timestamp 1625156677
transform -1 0 3948 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_7_1
timestamp 1625156677
transform -1 0 3956 0 -1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_348
timestamp 1625156677
transform -1 0 3988 0 -1 1105
box -2 -3 34 103
use INVX2  INVX2_81
timestamp 1625156677
transform -1 0 4004 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_378
timestamp 1625156677
transform -1 0 4028 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1625156677
transform -1 0 4124 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1625156677
transform 1 0 4124 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_379
timestamp 1625156677
transform -1 0 4244 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1625156677
transform -1 0 4340 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_188
timestamp 1625156677
transform 1 0 4340 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_108
timestamp 1625156677
transform 1 0 4364 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_160
timestamp 1625156677
transform -1 0 4412 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_190
timestamp 1625156677
transform 1 0 4412 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_8_0
timestamp 1625156677
transform 1 0 4436 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_8_1
timestamp 1625156677
transform 1 0 4444 0 -1 1105
box -2 -3 10 103
use BUFX2  BUFX2_71
timestamp 1625156677
transform 1 0 4452 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_106
timestamp 1625156677
transform 1 0 4476 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_115
timestamp 1625156677
transform -1 0 4524 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_107
timestamp 1625156677
transform 1 0 4524 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_106
timestamp 1625156677
transform 1 0 4548 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_157
timestamp 1625156677
transform -1 0 4604 0 -1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_81
timestamp 1625156677
transform -1 0 4660 0 -1 1105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_80
timestamp 1625156677
transform 1 0 4660 0 -1 1105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_209
timestamp 1625156677
transform 1 0 4716 0 -1 1105
box -2 -3 98 103
use XOR2X1  XOR2X1_111
timestamp 1625156677
transform -1 0 4868 0 -1 1105
box -2 -3 58 103
use NAND2X1  NAND2X1_211
timestamp 1625156677
transform 1 0 4868 0 -1 1105
box -2 -3 26 103
use OR2X2  OR2X2_81
timestamp 1625156677
transform -1 0 4924 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_62
timestamp 1625156677
transform 1 0 4924 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_9_0
timestamp 1625156677
transform -1 0 4964 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_9_1
timestamp 1625156677
transform -1 0 4972 0 -1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_118
timestamp 1625156677
transform -1 0 4996 0 -1 1105
box -2 -3 26 103
use XOR2X1  XOR2X1_93
timestamp 1625156677
transform -1 0 5052 0 -1 1105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_204
timestamp 1625156677
transform 1 0 5052 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_213
timestamp 1625156677
transform -1 0 5172 0 -1 1105
box -2 -3 26 103
use NOR3X1  NOR3X1_46
timestamp 1625156677
transform 1 0 5172 0 -1 1105
box -2 -3 66 103
use AND2X2  AND2X2_63
timestamp 1625156677
transform -1 0 5268 0 -1 1105
box -2 -3 34 103
use BUFX2  BUFX2_52
timestamp 1625156677
transform -1 0 5292 0 -1 1105
box -2 -3 26 103
use FILL  FILL_11_1
timestamp 1625156677
transform -1 0 5300 0 -1 1105
box -2 -3 10 103
use FILL  FILL_11_2
timestamp 1625156677
transform -1 0 5308 0 -1 1105
box -2 -3 10 103
use FILL  FILL_11_3
timestamp 1625156677
transform -1 0 5316 0 -1 1105
box -2 -3 10 103
use BUFX2  BUFX2_93
timestamp 1625156677
transform -1 0 28 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_90
timestamp 1625156677
transform -1 0 52 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_148
timestamp 1625156677
transform -1 0 76 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_186
timestamp 1625156677
transform 1 0 76 0 1 905
box -2 -3 26 103
use INVX1  INVX1_239
timestamp 1625156677
transform -1 0 116 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_375
timestamp 1625156677
transform 1 0 116 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_376
timestamp 1625156677
transform -1 0 164 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_211
timestamp 1625156677
transform -1 0 188 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_333
timestamp 1625156677
transform 1 0 188 0 1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_148
timestamp 1625156677
transform 1 0 220 0 1 905
box -2 -3 58 103
use NOR2X1  NOR2X1_182
timestamp 1625156677
transform 1 0 276 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_181
timestamp 1625156677
transform 1 0 300 0 1 905
box -2 -3 26 103
use INVX1  INVX1_190
timestamp 1625156677
transform -1 0 340 0 1 905
box -2 -3 18 103
use FILL  FILL_9_0_0
timestamp 1625156677
transform 1 0 340 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1625156677
transform 1 0 348 0 1 905
box -2 -3 10 103
use NAND3X1  NAND3X1_302
timestamp 1625156677
transform 1 0 356 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_284
timestamp 1625156677
transform -1 0 420 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_290
timestamp 1625156677
transform -1 0 452 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_294
timestamp 1625156677
transform -1 0 484 0 1 905
box -2 -3 34 103
use INVX2  INVX2_59
timestamp 1625156677
transform -1 0 500 0 1 905
box -2 -3 18 103
use INVX1  INVX1_192
timestamp 1625156677
transform 1 0 500 0 1 905
box -2 -3 18 103
use NAND3X1  NAND3X1_296
timestamp 1625156677
transform -1 0 548 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_205
timestamp 1625156677
transform -1 0 580 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_330
timestamp 1625156677
transform -1 0 604 0 1 905
box -2 -3 26 103
use INVX1  INVX1_191
timestamp 1625156677
transform -1 0 620 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_329
timestamp 1625156677
transform 1 0 620 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_295
timestamp 1625156677
transform -1 0 676 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_286
timestamp 1625156677
transform -1 0 708 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_183
timestamp 1625156677
transform -1 0 732 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_252
timestamp 1625156677
transform -1 0 828 0 1 905
box -2 -3 98 103
use OAI21X1  OAI21X1_100
timestamp 1625156677
transform -1 0 860 0 1 905
box -2 -3 34 103
use FILL  FILL_9_1_0
timestamp 1625156677
transform 1 0 860 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1625156677
transform 1 0 868 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_101
timestamp 1625156677
transform 1 0 876 0 1 905
box -2 -3 34 103
use INVX1  INVX1_69
timestamp 1625156677
transform -1 0 924 0 1 905
box -2 -3 18 103
use NAND3X1  NAND3X1_102
timestamp 1625156677
transform 1 0 924 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_104
timestamp 1625156677
transform -1 0 988 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_105
timestamp 1625156677
transform 1 0 988 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_103
timestamp 1625156677
transform -1 0 1052 0 1 905
box -2 -3 34 103
use BUFX2  BUFX2_254
timestamp 1625156677
transform 1 0 1052 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_124
timestamp 1625156677
transform 1 0 1076 0 1 905
box -2 -3 26 103
use AND2X2  AND2X2_36
timestamp 1625156677
transform 1 0 1100 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_75
timestamp 1625156677
transform 1 0 1132 0 1 905
box -2 -3 26 103
use INVX1  INVX1_71
timestamp 1625156677
transform -1 0 1172 0 1 905
box -2 -3 18 103
use XNOR2X1  XNOR2X1_53
timestamp 1625156677
transform -1 0 1228 0 1 905
box -2 -3 58 103
use NAND2X1  NAND2X1_132
timestamp 1625156677
transform -1 0 1252 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_82
timestamp 1625156677
transform 1 0 1252 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_123
timestamp 1625156677
transform 1 0 1284 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_163
timestamp 1625156677
transform -1 0 1404 0 1 905
box -2 -3 98 103
use FILL  FILL_9_2_0
timestamp 1625156677
transform -1 0 1412 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1625156677
transform -1 0 1420 0 1 905
box -2 -3 10 103
use NAND3X1  NAND3X1_111
timestamp 1625156677
transform -1 0 1452 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_119
timestamp 1625156677
transform -1 0 1476 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_415
timestamp 1625156677
transform 1 0 1476 0 1 905
box -2 -3 26 103
use OR2X2  OR2X2_41
timestamp 1625156677
transform 1 0 1500 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_95
timestamp 1625156677
transform -1 0 1564 0 1 905
box -2 -3 34 103
use INVX1  INVX1_66
timestamp 1625156677
transform 1 0 1564 0 1 905
box -2 -3 18 103
use NOR3X1  NOR3X1_35
timestamp 1625156677
transform -1 0 1644 0 1 905
box -2 -3 66 103
use NOR2X1  NOR2X1_68
timestamp 1625156677
transform -1 0 1668 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_93
timestamp 1625156677
transform 1 0 1668 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_96
timestamp 1625156677
transform 1 0 1700 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_117
timestamp 1625156677
transform 1 0 1732 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_81
timestamp 1625156677
transform -1 0 1788 0 1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_51
timestamp 1625156677
transform 1 0 1788 0 1 905
box -2 -3 58 103
use NAND2X1  NAND2X1_115
timestamp 1625156677
transform -1 0 1868 0 1 905
box -2 -3 26 103
use FILL  FILL_9_3_0
timestamp 1625156677
transform 1 0 1868 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1625156677
transform 1 0 1876 0 1 905
box -2 -3 10 103
use XNOR2X1  XNOR2X1_50
timestamp 1625156677
transform 1 0 1884 0 1 905
box -2 -3 58 103
use INVX2  INVX2_26
timestamp 1625156677
transform -1 0 1956 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_162
timestamp 1625156677
transform -1 0 2052 0 1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_409
timestamp 1625156677
transform -1 0 2076 0 1 905
box -2 -3 26 103
use INVX1  INVX1_499
timestamp 1625156677
transform 1 0 2076 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_595
timestamp 1625156677
transform 1 0 2092 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_356
timestamp 1625156677
transform 1 0 2124 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_236
timestamp 1625156677
transform 1 0 2156 0 1 905
box -2 -3 98 103
use INVX1  INVX1_166
timestamp 1625156677
transform 1 0 2252 0 1 905
box -2 -3 18 103
use CLKBUF1  CLKBUF1_47
timestamp 1625156677
transform -1 0 2340 0 1 905
box -2 -3 74 103
use NAND3X1  NAND3X1_261
timestamp 1625156677
transform -1 0 2372 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_260
timestamp 1625156677
transform -1 0 2404 0 1 905
box -2 -3 34 103
use FILL  FILL_9_4_0
timestamp 1625156677
transform -1 0 2412 0 1 905
box -2 -3 10 103
use FILL  FILL_9_4_1
timestamp 1625156677
transform -1 0 2420 0 1 905
box -2 -3 10 103
use INVX1  INVX1_167
timestamp 1625156677
transform -1 0 2436 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_248
timestamp 1625156677
transform -1 0 2468 0 1 905
box -2 -3 34 103
use NOR3X1  NOR3X1_54
timestamp 1625156677
transform 1 0 2468 0 1 905
box -2 -3 66 103
use NOR2X1  NOR2X1_159
timestamp 1625156677
transform -1 0 2556 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_292
timestamp 1625156677
transform -1 0 2580 0 1 905
box -2 -3 26 103
use AND2X2  AND2X2_88
timestamp 1625156677
transform -1 0 2612 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_237
timestamp 1625156677
transform -1 0 2708 0 1 905
box -2 -3 98 103
use XOR2X1  XOR2X1_66
timestamp 1625156677
transform 1 0 2708 0 1 905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_238
timestamp 1625156677
transform 1 0 2764 0 1 905
box -2 -3 98 103
use INVX1  INVX1_168
timestamp 1625156677
transform -1 0 2876 0 1 905
box -2 -3 18 103
use FILL  FILL_9_5_0
timestamp 1625156677
transform -1 0 2884 0 1 905
box -2 -3 10 103
use FILL  FILL_9_5_1
timestamp 1625156677
transform -1 0 2892 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1625156677
transform -1 0 2988 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1625156677
transform -1 0 3084 0 1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_359
timestamp 1625156677
transform 1 0 3084 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_360
timestamp 1625156677
transform 1 0 3108 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_358
timestamp 1625156677
transform 1 0 3132 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_612
timestamp 1625156677
transform 1 0 3156 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_569
timestamp 1625156677
transform -1 0 3212 0 1 905
box -2 -3 34 103
use INVX1  INVX1_473
timestamp 1625156677
transform -1 0 3228 0 1 905
box -2 -3 18 103
use AND2X2  AND2X2_168
timestamp 1625156677
transform -1 0 3260 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_13
timestamp 1625156677
transform -1 0 3292 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_361
timestamp 1625156677
transform 1 0 3292 0 1 905
box -2 -3 26 103
use INVX1  INVX1_474
timestamp 1625156677
transform -1 0 3332 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_615
timestamp 1625156677
transform 1 0 3332 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_388
timestamp 1625156677
transform 1 0 3356 0 1 905
box -2 -3 26 103
use INVX8  INVX8_2
timestamp 1625156677
transform -1 0 3420 0 1 905
box -2 -3 42 103
use FILL  FILL_9_6_0
timestamp 1625156677
transform 1 0 3420 0 1 905
box -2 -3 10 103
use FILL  FILL_9_6_1
timestamp 1625156677
transform 1 0 3428 0 1 905
box -2 -3 10 103
use INVX1  INVX1_472
timestamp 1625156677
transform 1 0 3436 0 1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_380
timestamp 1625156677
transform 1 0 3452 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_490
timestamp 1625156677
transform -1 0 3508 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_382
timestamp 1625156677
transform 1 0 3508 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_565
timestamp 1625156677
transform 1 0 3532 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_30
timestamp 1625156677
transform -1 0 3596 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_633
timestamp 1625156677
transform 1 0 3596 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_496
timestamp 1625156677
transform 1 0 3620 0 1 905
box -2 -3 34 103
use INVX1  INVX1_491
timestamp 1625156677
transform 1 0 3652 0 1 905
box -2 -3 18 103
use NAND3X1  NAND3X1_498
timestamp 1625156677
transform 1 0 3668 0 1 905
box -2 -3 34 103
use NOR3X1  NOR3X1_94
timestamp 1625156677
transform 1 0 3700 0 1 905
box -2 -3 66 103
use BUFX2  BUFX2_113
timestamp 1625156677
transform -1 0 3788 0 1 905
box -2 -3 26 103
use AND2X2  AND2X2_173
timestamp 1625156677
transform -1 0 3820 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_630
timestamp 1625156677
transform 1 0 3820 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_501
timestamp 1625156677
transform 1 0 3844 0 1 905
box -2 -3 34 103
use INVX1  INVX1_481
timestamp 1625156677
transform 1 0 3876 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_582
timestamp 1625156677
transform 1 0 3892 0 1 905
box -2 -3 34 103
use FILL  FILL_9_7_0
timestamp 1625156677
transform -1 0 3932 0 1 905
box -2 -3 10 103
use FILL  FILL_9_7_1
timestamp 1625156677
transform -1 0 3940 0 1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_340
timestamp 1625156677
transform -1 0 3972 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_502
timestamp 1625156677
transform 1 0 3972 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_637
timestamp 1625156677
transform 1 0 4004 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_407
timestamp 1625156677
transform -1 0 4052 0 1 905
box -2 -3 26 103
use OR2X2  OR2X2_130
timestamp 1625156677
transform 1 0 4052 0 1 905
box -2 -3 34 103
use NOR3X1  NOR3X1_95
timestamp 1625156677
transform -1 0 4148 0 1 905
box -2 -3 66 103
use AOI21X1  AOI21X1_349
timestamp 1625156677
transform 1 0 4148 0 1 905
box -2 -3 34 103
use INVX1  INVX1_485
timestamp 1625156677
transform -1 0 4196 0 1 905
box -2 -3 18 103
use NOR3X1  NOR3X1_96
timestamp 1625156677
transform 1 0 4196 0 1 905
box -2 -3 66 103
use OR2X2  OR2X2_72
timestamp 1625156677
transform 1 0 4260 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_166
timestamp 1625156677
transform 1 0 4292 0 1 905
box -2 -3 34 103
use INVX1  INVX1_109
timestamp 1625156677
transform 1 0 4324 0 1 905
box -2 -3 18 103
use OR2X2  OR2X2_70
timestamp 1625156677
transform -1 0 4372 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_114
timestamp 1625156677
transform 1 0 4372 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_105
timestamp 1625156677
transform 1 0 4404 0 1 905
box -2 -3 26 103
use INVX1  INVX1_104
timestamp 1625156677
transform -1 0 4444 0 1 905
box -2 -3 18 103
use FILL  FILL_9_8_0
timestamp 1625156677
transform -1 0 4452 0 1 905
box -2 -3 10 103
use FILL  FILL_9_8_1
timestamp 1625156677
transform -1 0 4460 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_158
timestamp 1625156677
transform -1 0 4492 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_159
timestamp 1625156677
transform -1 0 4524 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_164
timestamp 1625156677
transform -1 0 4556 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_180
timestamp 1625156677
transform 1 0 4556 0 1 905
box -2 -3 26 103
use INVX2  INVX2_37
timestamp 1625156677
transform -1 0 4596 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_189
timestamp 1625156677
transform 1 0 4596 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_118
timestamp 1625156677
transform -1 0 4652 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_154
timestamp 1625156677
transform -1 0 4684 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_116
timestamp 1625156677
transform 1 0 4684 0 1 905
box -2 -3 34 103
use INVX1  INVX1_107
timestamp 1625156677
transform -1 0 4732 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_153
timestamp 1625156677
transform -1 0 4764 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_148
timestamp 1625156677
transform 1 0 4764 0 1 905
box -2 -3 34 103
use XOR2X1  XOR2X1_90
timestamp 1625156677
transform 1 0 4796 0 1 905
box -2 -3 58 103
use NAND3X1  NAND3X1_165
timestamp 1625156677
transform -1 0 4884 0 1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_79
timestamp 1625156677
transform 1 0 4884 0 1 905
box -2 -3 58 103
use FILL  FILL_9_9_0
timestamp 1625156677
transform -1 0 4948 0 1 905
box -2 -3 10 103
use FILL  FILL_9_9_1
timestamp 1625156677
transform -1 0 4956 0 1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_117
timestamp 1625156677
transform -1 0 4988 0 1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_78
timestamp 1625156677
transform 1 0 4988 0 1 905
box -2 -3 58 103
use NAND2X1  NAND2X1_172
timestamp 1625156677
transform -1 0 5068 0 1 905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_77
timestamp 1625156677
transform 1 0 5068 0 1 905
box -2 -3 58 103
use INVX2  INVX2_35
timestamp 1625156677
transform -1 0 5140 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_186
timestamp 1625156677
transform -1 0 5236 0 1 905
box -2 -3 98 103
use BUFX2  BUFX2_271
timestamp 1625156677
transform 1 0 5236 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_222
timestamp 1625156677
transform -1 0 5284 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_101
timestamp 1625156677
transform 1 0 5284 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1625156677
transform 1 0 5308 0 1 905
box -2 -3 10 103
use BUFX2  BUFX2_126
timestamp 1625156677
transform -1 0 28 0 -1 905
box -2 -3 26 103
use BUFX2  BUFX2_39
timestamp 1625156677
transform -1 0 52 0 -1 905
box -2 -3 26 103
use BUFX2  BUFX2_45
timestamp 1625156677
transform -1 0 76 0 -1 905
box -2 -3 26 103
use BUFX2  BUFX2_144
timestamp 1625156677
transform 1 0 76 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_155
timestamp 1625156677
transform 1 0 100 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_272
timestamp 1625156677
transform -1 0 292 0 -1 905
box -2 -3 98 103
use CLKBUF1  CLKBUF1_33
timestamp 1625156677
transform -1 0 364 0 -1 905
box -2 -3 74 103
use FILL  FILL_8_0_0
timestamp 1625156677
transform 1 0 364 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1625156677
transform 1 0 372 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_331
timestamp 1625156677
transform 1 0 380 0 -1 905
box -2 -3 26 103
use NOR3X1  NOR3X1_57
timestamp 1625156677
transform -1 0 468 0 -1 905
box -2 -3 66 103
use NAND2X1  NAND2X1_328
timestamp 1625156677
transform -1 0 492 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_207
timestamp 1625156677
transform 1 0 492 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_199
timestamp 1625156677
transform -1 0 540 0 -1 905
box -2 -3 18 103
use INVX1  INVX1_534
timestamp 1625156677
transform -1 0 556 0 -1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_206
timestamp 1625156677
transform -1 0 588 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_335
timestamp 1625156677
transform -1 0 612 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_327
timestamp 1625156677
transform -1 0 636 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_189
timestamp 1625156677
transform -1 0 652 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_294
timestamp 1625156677
transform -1 0 684 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_180
timestamp 1625156677
transform -1 0 708 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_283
timestamp 1625156677
transform -1 0 740 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_166
timestamp 1625156677
transform 1 0 740 0 -1 905
box -2 -3 98 103
use AND2X2  AND2X2_35
timestamp 1625156677
transform -1 0 868 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_1_0
timestamp 1625156677
transform -1 0 876 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1625156677
transform -1 0 884 0 -1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_72
timestamp 1625156677
transform -1 0 908 0 -1 905
box -2 -3 26 103
use OR2X2  OR2X2_44
timestamp 1625156677
transform 1 0 908 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_122
timestamp 1625156677
transform -1 0 964 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_76
timestamp 1625156677
transform 1 0 964 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_107
timestamp 1625156677
transform 1 0 996 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_109
timestamp 1625156677
transform -1 0 1060 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_127
timestamp 1625156677
transform 1 0 1060 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_126
timestamp 1625156677
transform 1 0 1084 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_77
timestamp 1625156677
transform 1 0 1108 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_78
timestamp 1625156677
transform -1 0 1172 0 -1 905
box -2 -3 34 103
use OR2X2  OR2X2_46
timestamp 1625156677
transform 1 0 1172 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_103
timestamp 1625156677
transform 1 0 1204 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_107
timestamp 1625156677
transform -1 0 1268 0 -1 905
box -2 -3 34 103
use INVX2  INVX2_28
timestamp 1625156677
transform 1 0 1268 0 -1 905
box -2 -3 18 103
use NAND3X1  NAND3X1_110
timestamp 1625156677
transform 1 0 1284 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_106
timestamp 1625156677
transform 1 0 1316 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_2_0
timestamp 1625156677
transform -1 0 1356 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1625156677
transform -1 0 1364 0 -1 905
box -2 -3 10 103
use XNOR2X1  XNOR2X1_54
timestamp 1625156677
transform -1 0 1420 0 -1 905
box -2 -3 58 103
use OAI21X1  OAI21X1_108
timestamp 1625156677
transform 1 0 1420 0 -1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_52
timestamp 1625156677
transform 1 0 1452 0 -1 905
box -2 -3 58 103
use BUFX2  BUFX2_262
timestamp 1625156677
transform 1 0 1508 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_116
timestamp 1625156677
transform 1 0 1532 0 -1 905
box -2 -3 26 103
use XOR2X1  XOR2X1_67
timestamp 1625156677
transform 1 0 1556 0 -1 905
box -2 -3 58 103
use AND2X2  AND2X2_32
timestamp 1625156677
transform -1 0 1644 0 -1 905
box -2 -3 34 103
use XOR2X1  XOR2X1_42
timestamp 1625156677
transform 1 0 1644 0 -1 905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_49
timestamp 1625156677
transform -1 0 1756 0 -1 905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_185
timestamp 1625156677
transform 1 0 1756 0 -1 905
box -2 -3 98 103
use XOR2X1  XOR2X1_81
timestamp 1625156677
transform -1 0 1908 0 -1 905
box -2 -3 58 103
use FILL  FILL_8_3_0
timestamp 1625156677
transform -1 0 1916 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1625156677
transform -1 0 1924 0 -1 905
box -2 -3 10 103
use XNOR2X1  XNOR2X1_74
timestamp 1625156677
transform -1 0 1980 0 -1 905
box -2 -3 58 103
use NAND2X1  NAND2X1_166
timestamp 1625156677
transform -1 0 2004 0 -1 905
box -2 -3 26 103
use OR2X2  OR2X2_63
timestamp 1625156677
transform 1 0 2004 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_167
timestamp 1625156677
transform 1 0 2036 0 -1 905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_75
timestamp 1625156677
transform -1 0 2116 0 -1 905
box -2 -3 58 103
use NAND3X1  NAND3X1_259
timestamp 1625156677
transform -1 0 2148 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_179
timestamp 1625156677
transform 1 0 2148 0 -1 905
box -2 -3 34 103
use OR2X2  OR2X2_114
timestamp 1625156677
transform -1 0 2212 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_289
timestamp 1625156677
transform -1 0 2236 0 -1 905
box -2 -3 26 103
use AND2X2  AND2X2_87
timestamp 1625156677
transform 1 0 2236 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_152
timestamp 1625156677
transform 1 0 2268 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_180
timestamp 1625156677
transform -1 0 2324 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_251
timestamp 1625156677
transform -1 0 2356 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_252
timestamp 1625156677
transform 1 0 2356 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_4_0
timestamp 1625156677
transform 1 0 2388 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_4_1
timestamp 1625156677
transform 1 0 2396 0 -1 905
box -2 -3 10 103
use NAND3X1  NAND3X1_262
timestamp 1625156677
transform 1 0 2404 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_263
timestamp 1625156677
transform 1 0 2436 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_181
timestamp 1625156677
transform 1 0 2468 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_160
timestamp 1625156677
transform 1 0 2500 0 -1 905
box -2 -3 26 103
use OR2X2  OR2X2_115
timestamp 1625156677
transform -1 0 2556 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_182
timestamp 1625156677
transform 1 0 2556 0 -1 905
box -2 -3 34 103
use XOR2X1  XOR2X1_79
timestamp 1625156677
transform 1 0 2588 0 -1 905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1625156677
transform -1 0 2740 0 -1 905
box -2 -3 98 103
use XOR2X1  XOR2X1_76
timestamp 1625156677
transform -1 0 2796 0 -1 905
box -2 -3 58 103
use AND2X2  AND2X2_159
timestamp 1625156677
transform -1 0 2828 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1625156677
transform -1 0 2924 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_5_0
timestamp 1625156677
transform 1 0 2924 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_5_1
timestamp 1625156677
transform 1 0 2932 0 -1 905
box -2 -3 10 103
use AND2X2  AND2X2_158
timestamp 1625156677
transform 1 0 2940 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_475
timestamp 1625156677
transform 1 0 2972 0 -1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_362
timestamp 1625156677
transform -1 0 3012 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_327
timestamp 1625156677
transform -1 0 3044 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_489
timestamp 1625156677
transform 1 0 3044 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_572
timestamp 1625156677
transform -1 0 3108 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_614
timestamp 1625156677
transform -1 0 3132 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_611
timestamp 1625156677
transform 1 0 3132 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1625156677
transform -1 0 3252 0 -1 905
box -2 -3 98 103
use NAND3X1  NAND3X1_488
timestamp 1625156677
transform 1 0 3252 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_632
timestamp 1625156677
transform 1 0 3284 0 -1 905
box -2 -3 26 103
use AND2X2  AND2X2_169
timestamp 1625156677
transform -1 0 3340 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_384
timestamp 1625156677
transform 1 0 3340 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_566
timestamp 1625156677
transform -1 0 3396 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_610
timestamp 1625156677
transform -1 0 3420 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_6_0
timestamp 1625156677
transform 1 0 3420 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_6_1
timestamp 1625156677
transform 1 0 3428 0 -1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_383
timestamp 1625156677
transform 1 0 3436 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_387
timestamp 1625156677
transform 1 0 3460 0 -1 905
box -2 -3 26 103
use OR2X2  OR2X2_129
timestamp 1625156677
transform 1 0 3484 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1625156677
transform -1 0 3612 0 -1 905
box -2 -3 98 103
use NOR3X1  NOR3X1_91
timestamp 1625156677
transform 1 0 3612 0 -1 905
box -2 -3 66 103
use NAND2X1  NAND2X1_609
timestamp 1625156677
transform -1 0 3700 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_486
timestamp 1625156677
transform -1 0 3716 0 -1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_381
timestamp 1625156677
transform 1 0 3716 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_487
timestamp 1625156677
transform 1 0 3740 0 -1 905
box -2 -3 18 103
use NOR3X1  NOR3X1_89
timestamp 1625156677
transform 1 0 3756 0 -1 905
box -2 -3 66 103
use AND2X2  AND2X2_174
timestamp 1625156677
transform -1 0 3852 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_631
timestamp 1625156677
transform -1 0 3876 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_583
timestamp 1625156677
transform 1 0 3876 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_7_0
timestamp 1625156677
transform -1 0 3916 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_7_1
timestamp 1625156677
transform -1 0 3924 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1625156677
transform -1 0 4020 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_341
timestamp 1625156677
transform 1 0 4020 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_495
timestamp 1625156677
transform -1 0 4084 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_482
timestamp 1625156677
transform 1 0 4084 0 -1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_372
timestamp 1625156677
transform -1 0 4124 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1625156677
transform -1 0 4220 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1625156677
transform -1 0 4316 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_187
timestamp 1625156677
transform -1 0 4340 0 -1 905
box -2 -3 26 103
use BUFX2  BUFX2_127
timestamp 1625156677
transform -1 0 4364 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_184
timestamp 1625156677
transform -1 0 4388 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_163
timestamp 1625156677
transform 1 0 4388 0 -1 905
box -2 -3 34 103
use BUFX2  BUFX2_265
timestamp 1625156677
transform 1 0 4420 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_8_0
timestamp 1625156677
transform 1 0 4444 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_8_1
timestamp 1625156677
transform 1 0 4452 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_179
timestamp 1625156677
transform 1 0 4460 0 -1 905
box -2 -3 26 103
use OR2X2  OR2X2_68
timestamp 1625156677
transform 1 0 4484 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_112
timestamp 1625156677
transform 1 0 4516 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_102
timestamp 1625156677
transform 1 0 4548 0 -1 905
box -2 -3 18 103
use NAND3X1  NAND3X1_156
timestamp 1625156677
transform 1 0 4564 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_158
timestamp 1625156677
transform -1 0 4628 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_183
timestamp 1625156677
transform -1 0 4652 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_113
timestamp 1625156677
transform 1 0 4652 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_181
timestamp 1625156677
transform -1 0 4708 0 -1 905
box -2 -3 26 103
use AND2X2  AND2X2_54
timestamp 1625156677
transform 1 0 4708 0 -1 905
box -2 -3 34 103
use INVX2  INVX2_36
timestamp 1625156677
transform -1 0 4756 0 -1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_109
timestamp 1625156677
transform 1 0 4756 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_101
timestamp 1625156677
transform -1 0 4812 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_111
timestamp 1625156677
transform -1 0 4844 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_103
timestamp 1625156677
transform -1 0 4868 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_177
timestamp 1625156677
transform 1 0 4868 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_147
timestamp 1625156677
transform 1 0 4892 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_145
timestamp 1625156677
transform 1 0 4924 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_9_0
timestamp 1625156677
transform -1 0 4964 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_9_1
timestamp 1625156677
transform -1 0 4972 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_176
timestamp 1625156677
transform -1 0 4996 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_174
timestamp 1625156677
transform -1 0 5020 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_150
timestamp 1625156677
transform 1 0 5020 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_49
timestamp 1625156677
transform 1 0 5052 0 -1 905
box -2 -3 74 103
use XNOR2X1  XNOR2X1_76
timestamp 1625156677
transform 1 0 5124 0 -1 905
box -2 -3 58 103
use XOR2X1  XOR2X1_72
timestamp 1625156677
transform -1 0 5236 0 -1 905
box -2 -3 58 103
use BUFX2  BUFX2_70
timestamp 1625156677
transform -1 0 5260 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_133
timestamp 1625156677
transform -1 0 5292 0 -1 905
box -2 -3 34 103
use FILL  FILL_9_1
timestamp 1625156677
transform -1 0 5300 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_2
timestamp 1625156677
transform -1 0 5308 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_3
timestamp 1625156677
transform -1 0 5316 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_156
timestamp 1625156677
transform 1 0 4 0 1 705
box -2 -3 98 103
use AND2X2  AND2X2_27
timestamp 1625156677
transform 1 0 100 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_59
timestamp 1625156677
transform -1 0 156 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_63
timestamp 1625156677
transform -1 0 180 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_77
timestamp 1625156677
transform 1 0 180 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_63
timestamp 1625156677
transform 1 0 212 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_100
timestamp 1625156677
transform -1 0 268 0 1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_43
timestamp 1625156677
transform 1 0 268 0 1 705
box -2 -3 58 103
use NAND3X1  NAND3X1_78
timestamp 1625156677
transform 1 0 324 0 1 705
box -2 -3 34 103
use FILL  FILL_7_0_0
timestamp 1625156677
transform 1 0 356 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1625156677
transform 1 0 364 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_98
timestamp 1625156677
transform 1 0 372 0 1 705
box -2 -3 26 103
use INVX1  INVX1_63
timestamp 1625156677
transform 1 0 396 0 1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_68
timestamp 1625156677
transform 1 0 412 0 1 705
box -2 -3 34 103
use INVX2  INVX2_24
timestamp 1625156677
transform -1 0 460 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_61
timestamp 1625156677
transform -1 0 484 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_93
timestamp 1625156677
transform -1 0 516 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_70
timestamp 1625156677
transform 1 0 516 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_69
timestamp 1625156677
transform -1 0 580 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_96
timestamp 1625156677
transform 1 0 580 0 1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_42
timestamp 1625156677
transform -1 0 660 0 1 705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_41
timestamp 1625156677
transform 1 0 660 0 1 705
box -2 -3 58 103
use INVX2  INVX2_23
timestamp 1625156677
transform -1 0 732 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_154
timestamp 1625156677
transform -1 0 828 0 1 705
box -2 -3 98 103
use BUFX2  BUFX2_257
timestamp 1625156677
transform 1 0 828 0 1 705
box -2 -3 26 103
use FILL  FILL_7_1_0
timestamp 1625156677
transform 1 0 852 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1625156677
transform 1 0 860 0 1 705
box -2 -3 10 103
use XNOR2X1  XNOR2X1_44
timestamp 1625156677
transform 1 0 868 0 1 705
box -2 -3 58 103
use NAND2X1  NAND2X1_113
timestamp 1625156677
transform -1 0 948 0 1 705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_44
timestamp 1625156677
transform 1 0 948 0 1 705
box -2 -3 74 103
use OR2X2  OR2X2_45
timestamp 1625156677
transform 1 0 1020 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_105
timestamp 1625156677
transform -1 0 1084 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_104
timestamp 1625156677
transform 1 0 1084 0 1 705
box -2 -3 34 103
use INVX1  INVX1_70
timestamp 1625156677
transform 1 0 1116 0 1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_106
timestamp 1625156677
transform 1 0 1132 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_108
timestamp 1625156677
transform -1 0 1196 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_167
timestamp 1625156677
transform -1 0 1292 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_130
timestamp 1625156677
transform 1 0 1292 0 1 705
box -2 -3 26 103
use OR2X2  OR2X2_48
timestamp 1625156677
transform 1 0 1316 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_79
timestamp 1625156677
transform 1 0 1348 0 1 705
box -2 -3 34 103
use FILL  FILL_7_2_0
timestamp 1625156677
transform 1 0 1380 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1625156677
transform 1 0 1388 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_131
timestamp 1625156677
transform 1 0 1396 0 1 705
box -2 -3 26 103
use INVX1  INVX1_73
timestamp 1625156677
transform 1 0 1420 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_76
timestamp 1625156677
transform -1 0 1460 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_112
timestamp 1625156677
transform -1 0 1492 0 1 705
box -2 -3 34 103
use INVX1  INVX1_76
timestamp 1625156677
transform 1 0 1492 0 1 705
box -2 -3 18 103
use INVX1  INVX1_75
timestamp 1625156677
transform 1 0 1508 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_109
timestamp 1625156677
transform -1 0 1556 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_133
timestamp 1625156677
transform 1 0 1556 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_77
timestamp 1625156677
transform 1 0 1580 0 1 705
box -2 -3 26 103
use XOR2X1  XOR2X1_43
timestamp 1625156677
transform 1 0 1604 0 1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_68
timestamp 1625156677
transform 1 0 1660 0 1 705
box -2 -3 58 103
use BUFX2  BUFX2_255
timestamp 1625156677
transform 1 0 1716 0 1 705
box -2 -3 26 103
use INVX1  INVX1_509
timestamp 1625156677
transform -1 0 1756 0 1 705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_64
timestamp 1625156677
transform -1 0 1812 0 1 705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_73
timestamp 1625156677
transform -1 0 1868 0 1 705
box -2 -3 58 103
use INVX1  INVX1_521
timestamp 1625156677
transform -1 0 1884 0 1 705
box -2 -3 18 103
use FILL  FILL_7_3_0
timestamp 1625156677
transform -1 0 1892 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1625156677
transform -1 0 1900 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_147
timestamp 1625156677
transform -1 0 1924 0 1 705
box -2 -3 26 103
use OR2X2  OR2X2_55
timestamp 1625156677
transform 1 0 1924 0 1 705
box -2 -3 34 103
use INVX1  INVX1_83
timestamp 1625156677
transform -1 0 1972 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_176
timestamp 1625156677
transform -1 0 2068 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_148
timestamp 1625156677
transform 1 0 2068 0 1 705
box -2 -3 26 103
use INVX1  INVX1_94
timestamp 1625156677
transform -1 0 2108 0 1 705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_66
timestamp 1625156677
transform -1 0 2164 0 1 705
box -2 -3 58 103
use INVX1  INVX1_512
timestamp 1625156677
transform -1 0 2180 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_149
timestamp 1625156677
transform -1 0 2204 0 1 705
box -2 -3 26 103
use OR2X2  OR2X2_56
timestamp 1625156677
transform 1 0 2204 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_150
timestamp 1625156677
transform 1 0 2236 0 1 705
box -2 -3 26 103
use INVX1  INVX1_524
timestamp 1625156677
transform 1 0 2260 0 1 705
box -2 -3 18 103
use NAND3X1  NAND3X1_130
timestamp 1625156677
transform 1 0 2276 0 1 705
box -2 -3 34 103
use INVX1  INVX1_86
timestamp 1625156677
transform 1 0 2308 0 1 705
box -2 -3 18 103
use INVX1  INVX1_87
timestamp 1625156677
transform 1 0 2324 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_126
timestamp 1625156677
transform -1 0 2372 0 1 705
box -2 -3 34 103
use INVX1  INVX1_82
timestamp 1625156677
transform 1 0 2372 0 1 705
box -2 -3 18 103
use FILL  FILL_7_4_0
timestamp 1625156677
transform -1 0 2396 0 1 705
box -2 -3 10 103
use FILL  FILL_7_4_1
timestamp 1625156677
transform -1 0 2404 0 1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_85
timestamp 1625156677
transform -1 0 2428 0 1 705
box -2 -3 26 103
use INVX1  INVX1_84
timestamp 1625156677
transform 1 0 2428 0 1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_91
timestamp 1625156677
transform -1 0 2476 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_125
timestamp 1625156677
transform -1 0 2508 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_124
timestamp 1625156677
transform -1 0 2540 0 1 705
box -2 -3 34 103
use INVX2  INVX2_31
timestamp 1625156677
transform -1 0 2556 0 1 705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_63
timestamp 1625156677
transform -1 0 2612 0 1 705
box -2 -3 58 103
use OAI21X1  OAI21X1_120
timestamp 1625156677
transform -1 0 2644 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_87
timestamp 1625156677
transform 1 0 2644 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_86
timestamp 1625156677
transform 1 0 2668 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_123
timestamp 1625156677
transform -1 0 2724 0 1 705
box -2 -3 34 103
use XOR2X1  XOR2X1_77
timestamp 1625156677
transform 1 0 2724 0 1 705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_62
timestamp 1625156677
transform 1 0 2780 0 1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_78
timestamp 1625156677
transform 1 0 2836 0 1 705
box -2 -3 58 103
use FILL  FILL_7_5_0
timestamp 1625156677
transform 1 0 2892 0 1 705
box -2 -3 10 103
use FILL  FILL_7_5_1
timestamp 1625156677
transform 1 0 2900 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_193
timestamp 1625156677
transform 1 0 2908 0 1 705
box -2 -3 98 103
use XOR2X1  XOR2X1_91
timestamp 1625156677
transform -1 0 3060 0 1 705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_83
timestamp 1625156677
transform -1 0 3116 0 1 705
box -2 -3 58 103
use OAI21X1  OAI21X1_567
timestamp 1625156677
transform -1 0 3148 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_323
timestamp 1625156677
transform -1 0 3180 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_385
timestamp 1625156677
transform -1 0 3204 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1625156677
transform 1 0 3204 0 1 705
box -2 -3 98 103
use INVX4  INVX4_2
timestamp 1625156677
transform -1 0 3324 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_571
timestamp 1625156677
transform 1 0 3324 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_386
timestamp 1625156677
transform 1 0 3356 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_326
timestamp 1625156677
transform 1 0 3380 0 1 705
box -2 -3 34 103
use FILL  FILL_7_6_0
timestamp 1625156677
transform 1 0 3412 0 1 705
box -2 -3 10 103
use FILL  FILL_7_6_1
timestamp 1625156677
transform 1 0 3420 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_570
timestamp 1625156677
transform 1 0 3428 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_325
timestamp 1625156677
transform 1 0 3460 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_33
timestamp 1625156677
transform -1 0 3524 0 1 705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_82
timestamp 1625156677
transform -1 0 3580 0 1 705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_84
timestamp 1625156677
transform 1 0 3580 0 1 705
box -2 -3 58 103
use OR2X2  OR2X2_71
timestamp 1625156677
transform -1 0 3668 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_185
timestamp 1625156677
transform 1 0 3668 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_186
timestamp 1625156677
transform 1 0 3692 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_497
timestamp 1625156677
transform 1 0 3716 0 1 705
box -2 -3 34 103
use XOR2X1  XOR2X1_314
timestamp 1625156677
transform -1 0 3804 0 1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_313
timestamp 1625156677
transform 1 0 3804 0 1 705
box -2 -3 58 103
use AND2X2  AND2X2_5
timestamp 1625156677
transform 1 0 3860 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_27
timestamp 1625156677
transform 1 0 3892 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_22
timestamp 1625156677
transform -1 0 3940 0 1 705
box -2 -3 26 103
use FILL  FILL_7_7_0
timestamp 1625156677
transform -1 0 3948 0 1 705
box -2 -3 10 103
use FILL  FILL_7_7_1
timestamp 1625156677
transform -1 0 3956 0 1 705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_15
timestamp 1625156677
transform -1 0 4028 0 1 705
box -2 -3 74 103
use XOR2X1  XOR2X1_312
timestamp 1625156677
transform -1 0 4084 0 1 705
box -2 -3 58 103
use NAND2X1  NAND2X1_26
timestamp 1625156677
transform 1 0 4084 0 1 705
box -2 -3 26 103
use OR2X2  OR2X2_3
timestamp 1625156677
transform -1 0 4140 0 1 705
box -2 -3 34 103
use AND2X2  AND2X2_4
timestamp 1625156677
transform 1 0 4140 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_191
timestamp 1625156677
transform 1 0 4172 0 1 705
box -2 -3 98 103
use NAND3X1  NAND3X1_162
timestamp 1625156677
transform 1 0 4268 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_160
timestamp 1625156677
transform -1 0 4332 0 1 705
box -2 -3 34 103
use INVX1  INVX1_103
timestamp 1625156677
transform -1 0 4348 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_156
timestamp 1625156677
transform -1 0 4380 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_155
timestamp 1625156677
transform -1 0 4412 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_161
timestamp 1625156677
transform -1 0 4444 0 1 705
box -2 -3 34 103
use FILL  FILL_7_8_0
timestamp 1625156677
transform 1 0 4444 0 1 705
box -2 -3 10 103
use FILL  FILL_7_8_1
timestamp 1625156677
transform 1 0 4452 0 1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_102
timestamp 1625156677
transform 1 0 4460 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_152
timestamp 1625156677
transform 1 0 4484 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_151
timestamp 1625156677
transform 1 0 4516 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_157
timestamp 1625156677
transform -1 0 4580 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_159
timestamp 1625156677
transform 1 0 4580 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_110
timestamp 1625156677
transform -1 0 4644 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_154
timestamp 1625156677
transform 1 0 4644 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_155
timestamp 1625156677
transform -1 0 4708 0 1 705
box -2 -3 34 103
use INVX1  INVX1_101
timestamp 1625156677
transform 1 0 4708 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_149
timestamp 1625156677
transform -1 0 4756 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_150
timestamp 1625156677
transform 1 0 4756 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_108
timestamp 1625156677
transform 1 0 4788 0 1 705
box -2 -3 34 103
use NOR3X1  NOR3X1_42
timestamp 1625156677
transform -1 0 4884 0 1 705
box -2 -3 66 103
use NOR2X1  NOR2X1_99
timestamp 1625156677
transform -1 0 4908 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_146
timestamp 1625156677
transform 1 0 4908 0 1 705
box -2 -3 34 103
use INVX1  INVX1_100
timestamp 1625156677
transform -1 0 4956 0 1 705
box -2 -3 18 103
use FILL  FILL_7_9_0
timestamp 1625156677
transform 1 0 4956 0 1 705
box -2 -3 10 103
use FILL  FILL_7_9_1
timestamp 1625156677
transform 1 0 4964 0 1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_153
timestamp 1625156677
transform 1 0 4972 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_152
timestamp 1625156677
transform 1 0 5004 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_98
timestamp 1625156677
transform -1 0 5060 0 1 705
box -2 -3 26 103
use AND2X2  AND2X2_50
timestamp 1625156677
transform -1 0 5092 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_173
timestamp 1625156677
transform 1 0 5092 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_149
timestamp 1625156677
transform 1 0 5116 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_187
timestamp 1625156677
transform -1 0 5244 0 1 705
box -2 -3 98 103
use XNOR2X1  XNOR2X1_98
timestamp 1625156677
transform 1 0 5244 0 1 705
box -2 -3 58 103
use FILL  FILL_8_1
timestamp 1625156677
transform 1 0 5300 0 1 705
box -2 -3 10 103
use FILL  FILL_8_2
timestamp 1625156677
transform 1 0 5308 0 1 705
box -2 -3 10 103
use BUFX2  BUFX2_79
timestamp 1625156677
transform -1 0 28 0 -1 705
box -2 -3 26 103
use BUFX2  BUFX2_104
timestamp 1625156677
transform -1 0 52 0 -1 705
box -2 -3 26 103
use BUFX2  BUFX2_72
timestamp 1625156677
transform 1 0 52 0 -1 705
box -2 -3 26 103
use BUFX2  BUFX2_42
timestamp 1625156677
transform 1 0 76 0 -1 705
box -2 -3 26 103
use NOR3X1  NOR3X1_34
timestamp 1625156677
transform -1 0 164 0 -1 705
box -2 -3 66 103
use OAI21X1  OAI21X1_78
timestamp 1625156677
transform 1 0 164 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_56
timestamp 1625156677
transform -1 0 212 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_99
timestamp 1625156677
transform 1 0 212 0 -1 705
box -2 -3 26 103
use OR2X2  OR2X2_34
timestamp 1625156677
transform 1 0 236 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_59
timestamp 1625156677
transform -1 0 300 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_79
timestamp 1625156677
transform 1 0 300 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_0_0
timestamp 1625156677
transform 1 0 332 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1625156677
transform 1 0 340 0 -1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_80
timestamp 1625156677
transform 1 0 348 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_81
timestamp 1625156677
transform -1 0 412 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_79
timestamp 1625156677
transform -1 0 444 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_61
timestamp 1625156677
transform -1 0 476 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_60
timestamp 1625156677
transform -1 0 508 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_101
timestamp 1625156677
transform -1 0 532 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_85
timestamp 1625156677
transform -1 0 564 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_80
timestamp 1625156677
transform 1 0 564 0 -1 705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_40
timestamp 1625156677
transform -1 0 652 0 -1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_50
timestamp 1625156677
transform -1 0 708 0 -1 705
box -2 -3 58 103
use CLKBUF1  CLKBUF1_7
timestamp 1625156677
transform 1 0 708 0 -1 705
box -2 -3 74 103
use NAND2X1  NAND2X1_104
timestamp 1625156677
transform 1 0 780 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_92
timestamp 1625156677
transform 1 0 804 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_65
timestamp 1625156677
transform 1 0 836 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_1_0
timestamp 1625156677
transform 1 0 868 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1625156677
transform 1 0 876 0 -1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_105
timestamp 1625156677
transform 1 0 884 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_30
timestamp 1625156677
transform 1 0 908 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_107
timestamp 1625156677
transform -1 0 964 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_89
timestamp 1625156677
transform -1 0 996 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_86
timestamp 1625156677
transform 1 0 996 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_25
timestamp 1625156677
transform 1 0 1028 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_90
timestamp 1625156677
transform 1 0 1044 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_91
timestamp 1625156677
transform 1 0 1076 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_66
timestamp 1625156677
transform 1 0 1108 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_74
timestamp 1625156677
transform 1 0 1132 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_67
timestamp 1625156677
transform 1 0 1156 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_125
timestamp 1625156677
transform -1 0 1204 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_37
timestamp 1625156677
transform -1 0 1236 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_114
timestamp 1625156677
transform 1 0 1236 0 -1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_45
timestamp 1625156677
transform -1 0 1316 0 -1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_56
timestamp 1625156677
transform 1 0 1316 0 -1 705
box -2 -3 58 103
use FILL  FILL_6_2_0
timestamp 1625156677
transform 1 0 1372 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1625156677
transform 1 0 1380 0 -1 705
box -2 -3 10 103
use XOR2X1  XOR2X1_57
timestamp 1625156677
transform 1 0 1388 0 -1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_303
timestamp 1625156677
transform 1 0 1444 0 -1 705
box -2 -3 58 103
use CLKBUF1  CLKBUF1_12
timestamp 1625156677
transform 1 0 1500 0 -1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_169
timestamp 1625156677
transform -1 0 1668 0 -1 705
box -2 -3 98 103
use XOR2X1  XOR2X1_44
timestamp 1625156677
transform 1 0 1668 0 -1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_58
timestamp 1625156677
transform -1 0 1780 0 -1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_59
timestamp 1625156677
transform -1 0 1836 0 -1 705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_213
timestamp 1625156677
transform 1 0 1836 0 -1 705
box -2 -3 58 103
use FILL  FILL_6_3_0
timestamp 1625156677
transform 1 0 1892 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1625156677
transform 1 0 1900 0 -1 705
box -2 -3 10 103
use XOR2X1  XOR2X1_69
timestamp 1625156677
transform 1 0 1908 0 -1 705
box -2 -3 58 103
use INVX1  INVX1_515
timestamp 1625156677
transform -1 0 1980 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_147
timestamp 1625156677
transform -1 0 2076 0 -1 705
box -2 -3 98 103
use XNOR2X1  XNOR2X1_65
timestamp 1625156677
transform -1 0 2132 0 -1 705
box -2 -3 58 103
use XOR2X1  XOR2X1_297
timestamp 1625156677
transform 1 0 2132 0 -1 705
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_175
timestamp 1625156677
transform 1 0 2188 0 -1 705
box -2 -3 98 103
use OR2X2  OR2X2_53
timestamp 1625156677
transform 1 0 2284 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_126
timestamp 1625156677
transform -1 0 2348 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_144
timestamp 1625156677
transform 1 0 2348 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_124
timestamp 1625156677
transform -1 0 2404 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_4_0
timestamp 1625156677
transform -1 0 2412 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_4_1
timestamp 1625156677
transform -1 0 2420 0 -1 705
box -2 -3 10 103
use INVX1  INVX1_81
timestamp 1625156677
transform -1 0 2436 0 -1 705
box -2 -3 18 103
use AND2X2  AND2X2_43
timestamp 1625156677
transform 1 0 2436 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_84
timestamp 1625156677
transform -1 0 2492 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_121
timestamp 1625156677
transform -1 0 2524 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_122
timestamp 1625156677
transform 1 0 2524 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_125
timestamp 1625156677
transform -1 0 2588 0 -1 705
box -2 -3 34 103
use OR2X2  OR2X2_54
timestamp 1625156677
transform -1 0 2620 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_90
timestamp 1625156677
transform 1 0 2620 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_146
timestamp 1625156677
transform 1 0 2652 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_127
timestamp 1625156677
transform 1 0 2676 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_145
timestamp 1625156677
transform 1 0 2708 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_89
timestamp 1625156677
transform 1 0 2732 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_143
timestamp 1625156677
transform -1 0 2788 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_42
timestamp 1625156677
transform 1 0 2788 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_151
timestamp 1625156677
transform 1 0 2820 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_94
timestamp 1625156677
transform -1 0 2876 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_128
timestamp 1625156677
transform 1 0 2876 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_5_0
timestamp 1625156677
transform 1 0 2908 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_5_1
timestamp 1625156677
transform 1 0 2916 0 -1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_142
timestamp 1625156677
transform 1 0 2924 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_119
timestamp 1625156677
transform -1 0 2980 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_139
timestamp 1625156677
transform -1 0 3004 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_114
timestamp 1625156677
transform 1 0 3004 0 -1 705
box -2 -3 34 103
use XOR2X1  XOR2X1_70
timestamp 1625156677
transform -1 0 3092 0 -1 705
box -2 -3 58 103
use XNOR2X1  XNOR2X1_61
timestamp 1625156677
transform -1 0 3148 0 -1 705
box -2 -3 58 103
use CLKBUF1  CLKBUF1_37
timestamp 1625156677
transform -1 0 3220 0 -1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1625156677
transform 1 0 3220 0 -1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_613
timestamp 1625156677
transform -1 0 3340 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1625156677
transform 1 0 3340 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_6_0
timestamp 1625156677
transform -1 0 3444 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_6_1
timestamp 1625156677
transform -1 0 3452 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1625156677
transform -1 0 3548 0 -1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_192
timestamp 1625156677
transform 1 0 3548 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_105
timestamp 1625156677
transform 1 0 3644 0 -1 705
box -2 -3 18 103
use BUFX2  BUFX2_146
timestamp 1625156677
transform -1 0 3684 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_17
timestamp 1625156677
transform -1 0 3716 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_19
timestamp 1625156677
transform -1 0 3748 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_20
timestamp 1625156677
transform -1 0 3780 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_24
timestamp 1625156677
transform -1 0 3804 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_7
timestamp 1625156677
transform -1 0 3836 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_15
timestamp 1625156677
transform 1 0 3836 0 -1 705
box -2 -3 34 103
use OR2X2  OR2X2_4
timestamp 1625156677
transform 1 0 3868 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_12
timestamp 1625156677
transform -1 0 3932 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_7_0
timestamp 1625156677
transform -1 0 3940 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_7_1
timestamp 1625156677
transform -1 0 3948 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_16
timestamp 1625156677
transform -1 0 3980 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_14
timestamp 1625156677
transform -1 0 3996 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_15
timestamp 1625156677
transform 1 0 3996 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_13
timestamp 1625156677
transform -1 0 4060 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_14
timestamp 1625156677
transform -1 0 4092 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1625156677
transform 1 0 4092 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1625156677
transform -1 0 4156 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_13
timestamp 1625156677
transform 1 0 4156 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_14
timestamp 1625156677
transform -1 0 4204 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_13
timestamp 1625156677
transform -1 0 4236 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_20
timestamp 1625156677
transform -1 0 4260 0 -1 705
box -2 -3 26 103
use XOR2X1  XOR2X1_75
timestamp 1625156677
transform 1 0 4260 0 -1 705
box -2 -3 58 103
use NAND2X1  NAND2X1_182
timestamp 1625156677
transform -1 0 4340 0 -1 705
box -2 -3 26 103
use OR2X2  OR2X2_69
timestamp 1625156677
transform -1 0 4372 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_104
timestamp 1625156677
transform 1 0 4372 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_55
timestamp 1625156677
transform -1 0 4428 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_8_0
timestamp 1625156677
transform 1 0 4428 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_8_1
timestamp 1625156677
transform 1 0 4436 0 -1 705
box -2 -3 10 103
use AND2X2  AND2X2_53
timestamp 1625156677
transform 1 0 4444 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_189
timestamp 1625156677
transform 1 0 4476 0 -1 705
box -2 -3 98 103
use XOR2X1  XOR2X1_74
timestamp 1625156677
transform 1 0 4572 0 -1 705
box -2 -3 58 103
use BUFX2  BUFX2_66
timestamp 1625156677
transform -1 0 4652 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_178
timestamp 1625156677
transform -1 0 4676 0 -1 705
box -2 -3 26 103
use OR2X2  OR2X2_67
timestamp 1625156677
transform -1 0 4708 0 -1 705
box -2 -3 34 103
use AND2X2  AND2X2_52
timestamp 1625156677
transform 1 0 4708 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_100
timestamp 1625156677
transform -1 0 4764 0 -1 705
box -2 -3 26 103
use XOR2X1  XOR2X1_73
timestamp 1625156677
transform 1 0 4764 0 -1 705
box -2 -3 58 103
use AND2X2  AND2X2_51
timestamp 1625156677
transform 1 0 4820 0 -1 705
box -2 -3 34 103
use OR2X2  OR2X2_66
timestamp 1625156677
transform 1 0 4852 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_175
timestamp 1625156677
transform -1 0 4908 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_107
timestamp 1625156677
transform 1 0 4908 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_9_0
timestamp 1625156677
transform -1 0 4948 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_9_1
timestamp 1625156677
transform -1 0 4956 0 -1 705
box -2 -3 10 103
use NAND3X1  NAND3X1_151
timestamp 1625156677
transform -1 0 4988 0 -1 705
box -2 -3 34 103
use NOR3X1  NOR3X1_41
timestamp 1625156677
transform -1 0 5052 0 -1 705
box -2 -3 66 103
use OAI21X1  OAI21X1_144
timestamp 1625156677
transform 1 0 5052 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_99
timestamp 1625156677
transform -1 0 5100 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_188
timestamp 1625156677
transform -1 0 5196 0 -1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_206
timestamp 1625156677
transform -1 0 5292 0 -1 705
box -2 -3 98 103
use FILL  FILL_7_1
timestamp 1625156677
transform -1 0 5300 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_2
timestamp 1625156677
transform -1 0 5308 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_3
timestamp 1625156677
transform -1 0 5316 0 -1 705
box -2 -3 10 103
use BUFX2  BUFX2_125
timestamp 1625156677
transform -1 0 28 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_139
timestamp 1625156677
transform 1 0 28 0 1 505
box -2 -3 98 103
use BUFX2  BUFX2_51
timestamp 1625156677
transform -1 0 148 0 1 505
box -2 -3 26 103
use OR2X2  OR2X2_33
timestamp 1625156677
transform 1 0 148 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_97
timestamp 1625156677
transform 1 0 180 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_77
timestamp 1625156677
transform -1 0 236 0 1 505
box -2 -3 34 103
use INVX1  INVX1_55
timestamp 1625156677
transform 1 0 236 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_76
timestamp 1625156677
transform -1 0 284 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_157
timestamp 1625156677
transform 1 0 284 0 1 505
box -2 -3 98 103
use FILL  FILL_5_0_0
timestamp 1625156677
transform -1 0 388 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1625156677
transform -1 0 396 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_82
timestamp 1625156677
transform -1 0 428 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_81
timestamp 1625156677
transform 1 0 428 0 1 505
box -2 -3 34 103
use INVX1  INVX1_57
timestamp 1625156677
transform 1 0 460 0 1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_83
timestamp 1625156677
transform 1 0 476 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_82
timestamp 1625156677
transform 1 0 508 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_62
timestamp 1625156677
transform 1 0 540 0 1 505
box -2 -3 34 103
use XOR2X1  XOR2X1_32
timestamp 1625156677
transform 1 0 572 0 1 505
box -2 -3 58 103
use NAND3X1  NAND3X1_87
timestamp 1625156677
transform -1 0 660 0 1 505
box -2 -3 34 103
use BUFX2  BUFX2_258
timestamp 1625156677
transform -1 0 684 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_66
timestamp 1625156677
transform 1 0 684 0 1 505
box -2 -3 34 103
use OR2X2  OR2X2_38
timestamp 1625156677
transform 1 0 716 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_108
timestamp 1625156677
transform -1 0 772 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_91
timestamp 1625156677
transform 1 0 772 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_65
timestamp 1625156677
transform 1 0 804 0 1 505
box -2 -3 26 103
use INVX1  INVX1_60
timestamp 1625156677
transform -1 0 844 0 1 505
box -2 -3 18 103
use FILL  FILL_5_1_0
timestamp 1625156677
transform 1 0 844 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1625156677
transform 1 0 852 0 1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_67
timestamp 1625156677
transform 1 0 860 0 1 505
box -2 -3 34 103
use INVX1  INVX1_62
timestamp 1625156677
transform 1 0 892 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_112
timestamp 1625156677
transform -1 0 932 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_111
timestamp 1625156677
transform -1 0 956 0 1 505
box -2 -3 26 103
use OR2X2  OR2X2_40
timestamp 1625156677
transform 1 0 956 0 1 505
box -2 -3 34 103
use BUFX2  BUFX2_251
timestamp 1625156677
transform 1 0 988 0 1 505
box -2 -3 26 103
use INVX1  INVX1_64
timestamp 1625156677
transform 1 0 1012 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_92
timestamp 1625156677
transform 1 0 1028 0 1 505
box -2 -3 34 103
use INVX1  INVX1_65
timestamp 1625156677
transform -1 0 1076 0 1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_94
timestamp 1625156677
transform 1 0 1076 0 1 505
box -2 -3 34 103
use XOR2X1  XOR2X1_46
timestamp 1625156677
transform -1 0 1164 0 1 505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_160
timestamp 1625156677
transform -1 0 1260 0 1 505
box -2 -3 98 103
use XNOR2X1  XNOR2X1_56
timestamp 1625156677
transform -1 0 1316 0 1 505
box -2 -3 58 103
use BUFX2  BUFX2_252
timestamp 1625156677
transform -1 0 1340 0 1 505
box -2 -3 26 103
use XOR2X1  XOR2X1_61
timestamp 1625156677
transform 1 0 1340 0 1 505
box -2 -3 58 103
use FILL  FILL_5_2_0
timestamp 1625156677
transform 1 0 1396 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1625156677
transform 1 0 1404 0 1 505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_57
timestamp 1625156677
transform 1 0 1412 0 1 505
box -2 -3 58 103
use NAND2X1  NAND2X1_129
timestamp 1625156677
transform -1 0 1492 0 1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_55
timestamp 1625156677
transform -1 0 1548 0 1 505
box -2 -3 58 103
use BUFX2  BUFX2_253
timestamp 1625156677
transform 1 0 1548 0 1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_32
timestamp 1625156677
transform 1 0 1572 0 1 505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_34
timestamp 1625156677
transform 1 0 1628 0 1 505
box -2 -3 58 103
use NAND2X1  NAND2X1_77
timestamp 1625156677
transform 1 0 1684 0 1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_33
timestamp 1625156677
transform -1 0 1764 0 1 505
box -2 -3 58 103
use NOR3X1  NOR3X1_31
timestamp 1625156677
transform -1 0 1828 0 1 505
box -2 -3 66 103
use OAI21X1  OAI21X1_59
timestamp 1625156677
transform 1 0 1828 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_48
timestamp 1625156677
transform 1 0 1860 0 1 505
box -2 -3 26 103
use FILL  FILL_5_3_0
timestamp 1625156677
transform -1 0 1892 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1625156677
transform -1 0 1900 0 1 505
box -2 -3 10 103
use AND2X2  AND2X2_20
timestamp 1625156677
transform -1 0 1932 0 1 505
box -2 -3 34 103
use INVX1  INVX1_44
timestamp 1625156677
transform -1 0 1948 0 1 505
box -2 -3 18 103
use BUFX2  BUFX2_256
timestamp 1625156677
transform 1 0 1948 0 1 505
box -2 -3 26 103
use INVX2  INVX2_20
timestamp 1625156677
transform -1 0 1988 0 1 505
box -2 -3 18 103
use INVX1  INVX1_527
timestamp 1625156677
transform -1 0 2004 0 1 505
box -2 -3 18 103
use INVX1  INVX1_518
timestamp 1625156677
transform -1 0 2020 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_146
timestamp 1625156677
transform -1 0 2116 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_184
timestamp 1625156677
transform -1 0 2212 0 1 505
box -2 -3 98 103
use BUFX2  BUFX2_91
timestamp 1625156677
transform -1 0 2236 0 1 505
box -2 -3 26 103
use XOR2X1  XOR2X1_54
timestamp 1625156677
transform 1 0 2236 0 1 505
box -2 -3 58 103
use AND2X2  AND2X2_41
timestamp 1625156677
transform -1 0 2324 0 1 505
box -2 -3 34 103
use OR2X2  OR2X2_52
timestamp 1625156677
transform 1 0 2324 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_141
timestamp 1625156677
transform 1 0 2356 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_82
timestamp 1625156677
transform -1 0 2404 0 1 505
box -2 -3 26 103
use FILL  FILL_5_4_0
timestamp 1625156677
transform 1 0 2404 0 1 505
box -2 -3 10 103
use FILL  FILL_5_4_1
timestamp 1625156677
transform 1 0 2412 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_117
timestamp 1625156677
transform 1 0 2420 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_118
timestamp 1625156677
transform 1 0 2452 0 1 505
box -2 -3 34 103
use INVX1  INVX1_80
timestamp 1625156677
transform 1 0 2484 0 1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_120
timestamp 1625156677
transform 1 0 2500 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_121
timestamp 1625156677
transform -1 0 2564 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_88
timestamp 1625156677
transform 1 0 2564 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_122
timestamp 1625156677
transform 1 0 2596 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_123
timestamp 1625156677
transform 1 0 2628 0 1 505
box -2 -3 34 103
use XOR2X1  XOR2X1_53
timestamp 1625156677
transform 1 0 2660 0 1 505
box -2 -3 58 103
use INVX2  INVX2_30
timestamp 1625156677
transform 1 0 2716 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_81
timestamp 1625156677
transform -1 0 2756 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_92
timestamp 1625156677
transform -1 0 2788 0 1 505
box -2 -3 34 103
use INVX1  INVX1_85
timestamp 1625156677
transform -1 0 2804 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_113
timestamp 1625156677
transform 1 0 2804 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_135
timestamp 1625156677
transform 1 0 2836 0 1 505
box -2 -3 26 103
use NOR3X1  NOR3X1_37
timestamp 1625156677
transform -1 0 2924 0 1 505
box -2 -3 66 103
use FILL  FILL_5_5_0
timestamp 1625156677
transform 1 0 2924 0 1 505
box -2 -3 10 103
use FILL  FILL_5_5_1
timestamp 1625156677
transform 1 0 2932 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_78
timestamp 1625156677
transform 1 0 2940 0 1 505
box -2 -3 26 103
use AND2X2  AND2X2_38
timestamp 1625156677
transform 1 0 2964 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_110
timestamp 1625156677
transform 1 0 2996 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_129
timestamp 1625156677
transform -1 0 3060 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_136
timestamp 1625156677
transform 1 0 3060 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_114
timestamp 1625156677
transform 1 0 3084 0 1 505
box -2 -3 34 103
use XOR2X1  XOR2X1_52
timestamp 1625156677
transform 1 0 3116 0 1 505
box -2 -3 58 103
use AOI21X1  AOI21X1_93
timestamp 1625156677
transform -1 0 3204 0 1 505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_58
timestamp 1625156677
transform -1 0 3260 0 1 505
box -2 -3 58 103
use NAND2X1  NAND2X1_134
timestamp 1625156677
transform 1 0 3260 0 1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_60
timestamp 1625156677
transform -1 0 3340 0 1 505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_59
timestamp 1625156677
transform -1 0 3396 0 1 505
box -2 -3 58 103
use BUFX2  BUFX2_32
timestamp 1625156677
transform 1 0 3396 0 1 505
box -2 -3 26 103
use FILL  FILL_5_6_0
timestamp 1625156677
transform -1 0 3428 0 1 505
box -2 -3 10 103
use FILL  FILL_5_6_1
timestamp 1625156677
transform -1 0 3436 0 1 505
box -2 -3 10 103
use XOR2X1  XOR2X1_16
timestamp 1625156677
transform -1 0 3492 0 1 505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_8
timestamp 1625156677
transform 1 0 3492 0 1 505
box -2 -3 58 103
use AND2X2  AND2X2_6
timestamp 1625156677
transform -1 0 3580 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_29
timestamp 1625156677
transform -1 0 3604 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_17
timestamp 1625156677
transform -1 0 3636 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_31
timestamp 1625156677
transform -1 0 3660 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_16
timestamp 1625156677
transform -1 0 3692 0 1 505
box -2 -3 34 103
use INVX1  INVX1_15
timestamp 1625156677
transform -1 0 3708 0 1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_18
timestamp 1625156677
transform 1 0 3708 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_19
timestamp 1625156677
transform 1 0 3740 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_32
timestamp 1625156677
transform -1 0 3796 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_18
timestamp 1625156677
transform 1 0 3796 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1625156677
transform -1 0 3852 0 1 505
box -2 -3 26 103
use OR2X2  OR2X2_5
timestamp 1625156677
transform -1 0 3884 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_14
timestamp 1625156677
transform -1 0 3916 0 1 505
box -2 -3 34 103
use FILL  FILL_5_7_0
timestamp 1625156677
transform 1 0 3916 0 1 505
box -2 -3 10 103
use FILL  FILL_5_7_1
timestamp 1625156677
transform 1 0 3924 0 1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_16
timestamp 1625156677
transform 1 0 3932 0 1 505
box -2 -3 34 103
use INVX1  INVX1_19
timestamp 1625156677
transform 1 0 3964 0 1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_20
timestamp 1625156677
transform 1 0 3980 0 1 505
box -2 -3 34 103
use INVX2  INVX2_12
timestamp 1625156677
transform -1 0 4028 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_21
timestamp 1625156677
transform -1 0 4052 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_12
timestamp 1625156677
transform -1 0 4084 0 1 505
box -2 -3 34 103
use BUFX2  BUFX2_76
timestamp 1625156677
transform 1 0 4084 0 1 505
box -2 -3 26 103
use BUFX2  BUFX2_264
timestamp 1625156677
transform 1 0 4108 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_13
timestamp 1625156677
transform -1 0 4164 0 1 505
box -2 -3 34 103
use NOR3X1  NOR3X1_26
timestamp 1625156677
transform -1 0 4228 0 1 505
box -2 -3 66 103
use INVX1  INVX1_12
timestamp 1625156677
transform 1 0 4228 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_10
timestamp 1625156677
transform -1 0 4276 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_19
timestamp 1625156677
transform -1 0 4300 0 1 505
box -2 -3 26 103
use AND2X2  AND2X2_3
timestamp 1625156677
transform -1 0 4332 0 1 505
box -2 -3 34 103
use XOR2X1  XOR2X1_311
timestamp 1625156677
transform -1 0 4388 0 1 505
box -2 -3 58 103
use BUFX2  BUFX2_87
timestamp 1625156677
transform 1 0 4388 0 1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_251
timestamp 1625156677
transform 1 0 4412 0 1 505
box -2 -3 58 103
use FILL  FILL_5_8_0
timestamp 1625156677
transform 1 0 4468 0 1 505
box -2 -3 10 103
use FILL  FILL_5_8_1
timestamp 1625156677
transform 1 0 4476 0 1 505
box -2 -3 10 103
use OR2X2  OR2X2_155
timestamp 1625156677
transform 1 0 4484 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_705
timestamp 1625156677
transform 1 0 4516 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_532
timestamp 1625156677
transform -1 0 4572 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_445
timestamp 1625156677
transform -1 0 4596 0 1 505
box -2 -3 26 103
use INVX1  INVX1_590
timestamp 1625156677
transform 1 0 4596 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_635
timestamp 1625156677
transform -1 0 4644 0 1 505
box -2 -3 34 103
use NOR3X1  NOR3X1_97
timestamp 1625156677
transform 1 0 4644 0 1 505
box -2 -3 66 103
use AND2X2  AND2X2_193
timestamp 1625156677
transform -1 0 4740 0 1 505
box -2 -3 34 103
use AND2X2  AND2X2_194
timestamp 1625156677
transform 1 0 4740 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_446
timestamp 1625156677
transform 1 0 4772 0 1 505
box -2 -3 26 103
use INVX1  INVX1_591
timestamp 1625156677
transform -1 0 4812 0 1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_394
timestamp 1625156677
transform -1 0 4844 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_534
timestamp 1625156677
transform -1 0 4876 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_707
timestamp 1625156677
transform -1 0 4900 0 1 505
box -2 -3 26 103
use OR2X2  OR2X2_156
timestamp 1625156677
transform -1 0 4932 0 1 505
box -2 -3 34 103
use FILL  FILL_5_9_0
timestamp 1625156677
transform 1 0 4932 0 1 505
box -2 -3 10 103
use FILL  FILL_5_9_1
timestamp 1625156677
transform 1 0 4940 0 1 505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_25
timestamp 1625156677
transform 1 0 4948 0 1 505
box -2 -3 74 103
use NOR2X1  NOR2X1_447
timestamp 1625156677
transform 1 0 5020 0 1 505
box -2 -3 26 103
use AND2X2  AND2X2_195
timestamp 1625156677
transform 1 0 5044 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1625156677
transform -1 0 5172 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1625156677
transform -1 0 5268 0 1 505
box -2 -3 98 103
use NAND3X1  NAND3X1_193
timestamp 1625156677
transform -1 0 5300 0 1 505
box -2 -3 34 103
use FILL  FILL_6_1
timestamp 1625156677
transform 1 0 5300 0 1 505
box -2 -3 10 103
use FILL  FILL_6_2
timestamp 1625156677
transform 1 0 5308 0 1 505
box -2 -3 10 103
use BUFX2  BUFX2_133
timestamp 1625156677
transform -1 0 28 0 -1 505
box -2 -3 26 103
use BUFX2  BUFX2_134
timestamp 1625156677
transform -1 0 52 0 -1 505
box -2 -3 26 103
use BUFX2  BUFX2_69
timestamp 1625156677
transform 1 0 52 0 -1 505
box -2 -3 26 103
use XOR2X1  XOR2X1_34
timestamp 1625156677
transform 1 0 76 0 -1 505
box -2 -3 58 103
use XOR2X1  XOR2X1_33
timestamp 1625156677
transform -1 0 188 0 -1 505
box -2 -3 58 103
use AND2X2  AND2X2_26
timestamp 1625156677
transform 1 0 188 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_58
timestamp 1625156677
transform -1 0 244 0 -1 505
box -2 -3 26 103
use NOR3X1  NOR3X1_33
timestamp 1625156677
transform 1 0 244 0 -1 505
box -2 -3 66 103
use BUFX2  BUFX2_248
timestamp 1625156677
transform 1 0 308 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_0_0
timestamp 1625156677
transform -1 0 340 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1625156677
transform -1 0 348 0 -1 505
box -2 -3 10 103
use XOR2X1  XOR2X1_35
timestamp 1625156677
transform -1 0 404 0 -1 505
box -2 -3 58 103
use NOR2X1  NOR2X1_60
timestamp 1625156677
transform -1 0 428 0 -1 505
box -2 -3 26 103
use AND2X2  AND2X2_28
timestamp 1625156677
transform -1 0 460 0 -1 505
box -2 -3 34 103
use OR2X2  OR2X2_35
timestamp 1625156677
transform 1 0 460 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_102
timestamp 1625156677
transform -1 0 516 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_158
timestamp 1625156677
transform 1 0 516 0 -1 505
box -2 -3 98 103
use NAND3X1  NAND3X1_86
timestamp 1625156677
transform -1 0 644 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_64
timestamp 1625156677
transform 1 0 644 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_85
timestamp 1625156677
transform 1 0 676 0 -1 505
box -2 -3 34 103
use AND2X2  AND2X2_31
timestamp 1625156677
transform 1 0 708 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_64
timestamp 1625156677
transform -1 0 764 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_88
timestamp 1625156677
transform 1 0 764 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_87
timestamp 1625156677
transform 1 0 796 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_89
timestamp 1625156677
transform 1 0 828 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_1_0
timestamp 1625156677
transform 1 0 860 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1625156677
transform 1 0 868 0 -1 505
box -2 -3 10 103
use INVX1  INVX1_59
timestamp 1625156677
transform 1 0 876 0 -1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_88
timestamp 1625156677
transform 1 0 892 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_106
timestamp 1625156677
transform 1 0 924 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_90
timestamp 1625156677
transform 1 0 948 0 -1 505
box -2 -3 34 103
use OR2X2  OR2X2_37
timestamp 1625156677
transform -1 0 1012 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_159
timestamp 1625156677
transform -1 0 1108 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_142
timestamp 1625156677
transform -1 0 1204 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_61
timestamp 1625156677
transform 1 0 1204 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_110
timestamp 1625156677
transform -1 0 1244 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_109
timestamp 1625156677
transform -1 0 1268 0 -1 505
box -2 -3 26 103
use OR2X2  OR2X2_39
timestamp 1625156677
transform 1 0 1268 0 -1 505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_48
timestamp 1625156677
transform -1 0 1356 0 -1 505
box -2 -3 58 103
use FILL  FILL_4_2_0
timestamp 1625156677
transform -1 0 1364 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1625156677
transform -1 0 1372 0 -1 505
box -2 -3 10 103
use XOR2X1  XOR2X1_48
timestamp 1625156677
transform -1 0 1428 0 -1 505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_168
timestamp 1625156677
transform 1 0 1428 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_72
timestamp 1625156677
transform 1 0 1524 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_128
timestamp 1625156677
transform -1 0 1564 0 -1 505
box -2 -3 26 103
use OR2X2  OR2X2_47
timestamp 1625156677
transform 1 0 1564 0 -1 505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_31
timestamp 1625156677
transform -1 0 1652 0 -1 505
box -2 -3 58 103
use BUFX2  BUFX2_240
timestamp 1625156677
transform 1 0 1652 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_75
timestamp 1625156677
transform -1 0 1708 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_57
timestamp 1625156677
transform 1 0 1708 0 -1 505
box -2 -3 34 103
use XOR2X1  XOR2X1_40
timestamp 1625156677
transform -1 0 1796 0 -1 505
box -2 -3 58 103
use OAI21X1  OAI21X1_63
timestamp 1625156677
transform -1 0 1828 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_60
timestamp 1625156677
transform -1 0 1860 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_79
timestamp 1625156677
transform 1 0 1860 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_3_0
timestamp 1625156677
transform -1 0 1892 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1625156677
transform -1 0 1900 0 -1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_81
timestamp 1625156677
transform -1 0 1924 0 -1 505
box -2 -3 26 103
use OR2X2  OR2X2_25
timestamp 1625156677
transform 1 0 1924 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_59
timestamp 1625156677
transform -1 0 1988 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_78
timestamp 1625156677
transform -1 0 2012 0 -1 505
box -2 -3 26 103
use XOR2X1  XOR2X1_23
timestamp 1625156677
transform 1 0 2012 0 -1 505
box -2 -3 58 103
use XOR2X1  XOR2X1_71
timestamp 1625156677
transform 1 0 2068 0 -1 505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_177
timestamp 1625156677
transform -1 0 2220 0 -1 505
box -2 -3 98 103
use XOR2X1  XOR2X1_55
timestamp 1625156677
transform 1 0 2220 0 -1 505
box -2 -3 58 103
use CLKBUF1  CLKBUF1_29
timestamp 1625156677
transform -1 0 2348 0 -1 505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_1
timestamp 1625156677
transform 1 0 2348 0 -1 505
box -2 -3 74 103
use FILL  FILL_4_4_0
timestamp 1625156677
transform 1 0 2420 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_4_1
timestamp 1625156677
transform 1 0 2428 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_174
timestamp 1625156677
transform 1 0 2436 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_171
timestamp 1625156677
transform 1 0 2532 0 -1 505
box -2 -3 98 103
use OR2X2  OR2X2_51
timestamp 1625156677
transform 1 0 2628 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_86
timestamp 1625156677
transform -1 0 2692 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_85
timestamp 1625156677
transform 1 0 2692 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_84
timestamp 1625156677
transform 1 0 2724 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_83
timestamp 1625156677
transform -1 0 2780 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_87
timestamp 1625156677
transform -1 0 2812 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_111
timestamp 1625156677
transform 1 0 2812 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_138
timestamp 1625156677
transform 1 0 2844 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_113
timestamp 1625156677
transform 1 0 2868 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_5_0
timestamp 1625156677
transform 1 0 2900 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_5_1
timestamp 1625156677
transform 1 0 2908 0 -1 505
box -2 -3 10 103
use INVX1  INVX1_77
timestamp 1625156677
transform 1 0 2916 0 -1 505
box -2 -3 18 103
use OR2X2  OR2X2_49
timestamp 1625156677
transform -1 0 2964 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_130
timestamp 1625156677
transform -1 0 3060 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_170
timestamp 1625156677
transform 1 0 3060 0 -1 505
box -2 -3 98 103
use INVX2  INVX2_29
timestamp 1625156677
transform 1 0 3156 0 -1 505
box -2 -3 18 103
use CLKBUF1  CLKBUF1_38
timestamp 1625156677
transform 1 0 3172 0 -1 505
box -2 -3 74 103
use XOR2X1  XOR2X1_17
timestamp 1625156677
transform -1 0 3300 0 -1 505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1625156677
transform 1 0 3300 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_6_0
timestamp 1625156677
transform 1 0 3396 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_6_1
timestamp 1625156677
transform 1 0 3404 0 -1 505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_9
timestamp 1625156677
transform 1 0 3412 0 -1 505
box -2 -3 58 103
use OAI21X1  OAI21X1_18
timestamp 1625156677
transform -1 0 3500 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_21
timestamp 1625156677
transform 1 0 3500 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_37
timestamp 1625156677
transform -1 0 3556 0 -1 505
box -2 -3 26 103
use INVX2  INVX2_13
timestamp 1625156677
transform 1 0 3556 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_28
timestamp 1625156677
transform -1 0 3596 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_20
timestamp 1625156677
transform 1 0 3596 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_23
timestamp 1625156677
transform -1 0 3660 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_22
timestamp 1625156677
transform 1 0 3660 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_16
timestamp 1625156677
transform 1 0 3692 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_25
timestamp 1625156677
transform -1 0 3732 0 -1 505
box -2 -3 26 103
use OR2X2  OR2X2_6
timestamp 1625156677
transform -1 0 3764 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_22
timestamp 1625156677
transform -1 0 3796 0 -1 505
box -2 -3 34 103
use XOR2X1  XOR2X1_10
timestamp 1625156677
transform -1 0 3852 0 -1 505
box -2 -3 58 103
use OAI21X1  OAI21X1_17
timestamp 1625156677
transform -1 0 3884 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_12
timestamp 1625156677
transform 1 0 3884 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_25
timestamp 1625156677
transform 1 0 3916 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_7_0
timestamp 1625156677
transform 1 0 3940 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_7_1
timestamp 1625156677
transform 1 0 3948 0 -1 505
box -2 -3 10 103
use NAND3X1  NAND3X1_9
timestamp 1625156677
transform 1 0 3956 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_15
timestamp 1625156677
transform -1 0 4020 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_9
timestamp 1625156677
transform -1 0 4052 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_23
timestamp 1625156677
transform 1 0 4052 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_11
timestamp 1625156677
transform -1 0 4108 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_11
timestamp 1625156677
transform -1 0 4140 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_7
timestamp 1625156677
transform 1 0 4140 0 -1 505
box -2 -3 34 103
use OR2X2  OR2X2_2
timestamp 1625156677
transform -1 0 4204 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_23
timestamp 1625156677
transform -1 0 4228 0 -1 505
box -2 -3 26 103
use BUFX2  BUFX2_92
timestamp 1625156677
transform -1 0 4252 0 -1 505
box -2 -3 26 103
use BUFX2  BUFX2_151
timestamp 1625156677
transform -1 0 4276 0 -1 505
box -2 -3 26 103
use BUFX2  BUFX2_152
timestamp 1625156677
transform 1 0 4276 0 -1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_252
timestamp 1625156677
transform 1 0 4300 0 -1 505
box -2 -3 58 103
use NAND2X1  NAND2X1_704
timestamp 1625156677
transform 1 0 4356 0 -1 505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_253
timestamp 1625156677
transform -1 0 4436 0 -1 505
box -2 -3 58 103
use FILL  FILL_4_8_0
timestamp 1625156677
transform 1 0 4436 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_8_1
timestamp 1625156677
transform 1 0 4444 0 -1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_404
timestamp 1625156677
transform 1 0 4452 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_533
timestamp 1625156677
transform -1 0 4516 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_706
timestamp 1625156677
transform -1 0 4540 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_535
timestamp 1625156677
transform -1 0 4572 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_638
timestamp 1625156677
transform -1 0 4604 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_536
timestamp 1625156677
transform 1 0 4604 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_636
timestamp 1625156677
transform -1 0 4668 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_398
timestamp 1625156677
transform 1 0 4668 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_93
timestamp 1625156677
transform -1 0 4716 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_450
timestamp 1625156677
transform -1 0 4740 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_637
timestamp 1625156677
transform -1 0 4772 0 -1 505
box -2 -3 34 103
use NOR3X1  NOR3X1_98
timestamp 1625156677
transform 1 0 4772 0 -1 505
box -2 -3 66 103
use AOI21X1  AOI21X1_396
timestamp 1625156677
transform -1 0 4868 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_395
timestamp 1625156677
transform -1 0 4900 0 -1 505
box -2 -3 34 103
use OR2X2  OR2X2_157
timestamp 1625156677
transform 1 0 4900 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_537
timestamp 1625156677
transform -1 0 4964 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_9_0
timestamp 1625156677
transform -1 0 4972 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_9_1
timestamp 1625156677
transform -1 0 4980 0 -1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_397
timestamp 1625156677
transform -1 0 5012 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_538
timestamp 1625156677
transform -1 0 5044 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_710
timestamp 1625156677
transform 1 0 5044 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_641
timestamp 1625156677
transform -1 0 5100 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_640
timestamp 1625156677
transform 1 0 5100 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_540
timestamp 1625156677
transform 1 0 5132 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_592
timestamp 1625156677
transform -1 0 5180 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1625156677
transform -1 0 5276 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_123
timestamp 1625156677
transform 1 0 5276 0 -1 505
box -2 -3 18 103
use FILL  FILL_5_1
timestamp 1625156677
transform -1 0 5300 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_2
timestamp 1625156677
transform -1 0 5308 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_3
timestamp 1625156677
transform -1 0 5316 0 -1 505
box -2 -3 10 103
use BUFX2  BUFX2_119
timestamp 1625156677
transform -1 0 28 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_138
timestamp 1625156677
transform 1 0 28 0 1 305
box -2 -3 98 103
use INVX2  INVX2_17
timestamp 1625156677
transform 1 0 124 0 1 305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_24
timestamp 1625156677
transform 1 0 140 0 1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_58
timestamp 1625156677
transform 1 0 196 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_45
timestamp 1625156677
transform -1 0 252 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_39
timestamp 1625156677
transform -1 0 276 0 1 305
box -2 -3 26 103
use AND2X2  AND2X2_15
timestamp 1625156677
transform -1 0 308 0 1 305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_23
timestamp 1625156677
transform -1 0 364 0 1 305
box -2 -3 58 103
use FILL  FILL_3_0_0
timestamp 1625156677
transform 1 0 364 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1625156677
transform 1 0 372 0 1 305
box -2 -3 10 103
use XNOR2X1  XNOR2X1_22
timestamp 1625156677
transform 1 0 380 0 1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_140
timestamp 1625156677
transform -1 0 532 0 1 305
box -2 -3 98 103
use OR2X2  OR2X2_36
timestamp 1625156677
transform 1 0 532 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_103
timestamp 1625156677
transform 1 0 564 0 1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_84
timestamp 1625156677
transform -1 0 620 0 1 305
box -2 -3 34 103
use INVX1  INVX1_58
timestamp 1625156677
transform -1 0 636 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_84
timestamp 1625156677
transform -1 0 668 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_83
timestamp 1625156677
transform -1 0 700 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_62
timestamp 1625156677
transform -1 0 724 0 1 305
box -2 -3 26 103
use AND2X2  AND2X2_29
timestamp 1625156677
transform -1 0 756 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_65
timestamp 1625156677
transform 1 0 756 0 1 305
box -2 -3 26 103
use OR2X2  OR2X2_20
timestamp 1625156677
transform -1 0 812 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_42
timestamp 1625156677
transform 1 0 812 0 1 305
box -2 -3 26 103
use AND2X2  AND2X2_17
timestamp 1625156677
transform -1 0 868 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1625156677
transform 1 0 868 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1625156677
transform 1 0 876 0 1 305
box -2 -3 10 103
use BUFX2  BUFX2_247
timestamp 1625156677
transform 1 0 884 0 1 305
box -2 -3 26 103
use BUFX2  BUFX2_198
timestamp 1625156677
transform -1 0 932 0 1 305
box -2 -3 26 103
use XOR2X1  XOR2X1_37
timestamp 1625156677
transform 1 0 932 0 1 305
box -2 -3 58 103
use XOR2X1  XOR2X1_47
timestamp 1625156677
transform -1 0 1044 0 1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_143
timestamp 1625156677
transform -1 0 1140 0 1 305
box -2 -3 98 103
use XNOR2X1  XNOR2X1_46
timestamp 1625156677
transform 1 0 1140 0 1 305
box -2 -3 58 103
use XOR2X1  XOR2X1_49
timestamp 1625156677
transform -1 0 1252 0 1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_95
timestamp 1625156677
transform 1 0 1252 0 1 305
box -2 -3 26 103
use INVX1  INVX1_54
timestamp 1625156677
transform 1 0 1276 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_75
timestamp 1625156677
transform -1 0 1324 0 1 305
box -2 -3 34 103
use INVX1  INVX1_53
timestamp 1625156677
transform -1 0 1340 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_55
timestamp 1625156677
transform -1 0 1372 0 1 305
box -2 -3 34 103
use FILL  FILL_3_2_0
timestamp 1625156677
transform 1 0 1372 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1625156677
transform 1 0 1380 0 1 305
box -2 -3 10 103
use NOR2X1  NOR2X1_57
timestamp 1625156677
transform 1 0 1388 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_56
timestamp 1625156677
transform 1 0 1412 0 1 305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_35
timestamp 1625156677
transform -1 0 1492 0 1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_94
timestamp 1625156677
transform 1 0 1492 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_72
timestamp 1625156677
transform -1 0 1548 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_74
timestamp 1625156677
transform -1 0 1580 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_85
timestamp 1625156677
transform -1 0 1604 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_58
timestamp 1625156677
transform -1 0 1636 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_56
timestamp 1625156677
transform -1 0 1668 0 1 305
box -2 -3 34 103
use INVX2  INVX2_21
timestamp 1625156677
transform -1 0 1684 0 1 305
box -2 -3 18 103
use INVX1  INVX1_52
timestamp 1625156677
transform -1 0 1700 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_51
timestamp 1625156677
transform -1 0 1724 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_68
timestamp 1625156677
transform -1 0 1756 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_51
timestamp 1625156677
transform -1 0 1788 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_53
timestamp 1625156677
transform -1 0 1812 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_82
timestamp 1625156677
transform 1 0 1812 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_62
timestamp 1625156677
transform 1 0 1836 0 1 305
box -2 -3 34 103
use FILL  FILL_3_3_0
timestamp 1625156677
transform 1 0 1868 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1625156677
transform 1 0 1876 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_60
timestamp 1625156677
transform 1 0 1884 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_63
timestamp 1625156677
transform -1 0 1948 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_62
timestamp 1625156677
transform 1 0 1948 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_149
timestamp 1625156677
transform -1 0 2076 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_61
timestamp 1625156677
transform 1 0 2076 0 1 305
box -2 -3 34 103
use NOR3X1  NOR3X1_32
timestamp 1625156677
transform 1 0 2108 0 1 305
box -2 -3 66 103
use INVX1  INVX1_45
timestamp 1625156677
transform -1 0 2188 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_47
timestamp 1625156677
transform -1 0 2220 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_61
timestamp 1625156677
transform 1 0 2220 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_148
timestamp 1625156677
transform -1 0 2348 0 1 305
box -2 -3 98 103
use XOR2X1  XOR2X1_31
timestamp 1625156677
transform -1 0 2404 0 1 305
box -2 -3 58 103
use FILL  FILL_3_4_0
timestamp 1625156677
transform 1 0 2404 0 1 305
box -2 -3 10 103
use FILL  FILL_3_4_1
timestamp 1625156677
transform 1 0 2412 0 1 305
box -2 -3 10 103
use XNOR2X1  XNOR2X1_29
timestamp 1625156677
transform 1 0 2420 0 1 305
box -2 -3 58 103
use AND2X2  AND2X2_40
timestamp 1625156677
transform 1 0 2476 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_80
timestamp 1625156677
transform 1 0 2508 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_116
timestamp 1625156677
transform 1 0 2532 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1625156677
transform 1 0 2564 0 1 305
box -2 -3 34 103
use INVX1  INVX1_79
timestamp 1625156677
transform -1 0 2612 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_140
timestamp 1625156677
transform 1 0 2612 0 1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_119
timestamp 1625156677
transform 1 0 2636 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_118
timestamp 1625156677
transform 1 0 2668 0 1 305
box -2 -3 34 103
use OR2X2  OR2X2_50
timestamp 1625156677
transform 1 0 2700 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_115
timestamp 1625156677
transform -1 0 2764 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_83
timestamp 1625156677
transform -1 0 2796 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_117
timestamp 1625156677
transform 1 0 2796 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_116
timestamp 1625156677
transform 1 0 2828 0 1 305
box -2 -3 34 103
use FILL  FILL_3_5_0
timestamp 1625156677
transform -1 0 2868 0 1 305
box -2 -3 10 103
use FILL  FILL_3_5_1
timestamp 1625156677
transform -1 0 2876 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_132
timestamp 1625156677
transform -1 0 2972 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_133
timestamp 1625156677
transform 1 0 2972 0 1 305
box -2 -3 98 103
use AND2X2  AND2X2_10
timestamp 1625156677
transform -1 0 3100 0 1 305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_28
timestamp 1625156677
transform 1 0 3100 0 1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_134
timestamp 1625156677
transform 1 0 3156 0 1 305
box -2 -3 98 103
use XOR2X1  XOR2X1_5
timestamp 1625156677
transform -1 0 3308 0 1 305
box -2 -3 58 103
use AND2X2  AND2X2_11
timestamp 1625156677
transform -1 0 3340 0 1 305
box -2 -3 34 103
use XOR2X1  XOR2X1_18
timestamp 1625156677
transform -1 0 3396 0 1 305
box -2 -3 58 103
use BUFX2  BUFX2_149
timestamp 1625156677
transform 1 0 3396 0 1 305
box -2 -3 26 103
use FILL  FILL_3_6_0
timestamp 1625156677
transform -1 0 3428 0 1 305
box -2 -3 10 103
use FILL  FILL_3_6_1
timestamp 1625156677
transform -1 0 3436 0 1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_46
timestamp 1625156677
transform -1 0 3460 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_27
timestamp 1625156677
transform -1 0 3484 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_26
timestamp 1625156677
transform -1 0 3508 0 1 305
box -2 -3 26 103
use INVX1  INVX1_18
timestamp 1625156677
transform -1 0 3524 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_19
timestamp 1625156677
transform -1 0 3556 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_36
timestamp 1625156677
transform -1 0 3580 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_35
timestamp 1625156677
transform -1 0 3604 0 1 305
box -2 -3 26 103
use OR2X2  OR2X2_8
timestamp 1625156677
transform 1 0 3604 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_22
timestamp 1625156677
transform 1 0 3636 0 1 305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_6
timestamp 1625156677
transform 1 0 3668 0 1 305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_7
timestamp 1625156677
transform 1 0 3724 0 1 305
box -2 -3 58 103
use NAND3X1  NAND3X1_21
timestamp 1625156677
transform 1 0 3780 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_6
timestamp 1625156677
transform -1 0 3844 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_22
timestamp 1625156677
transform -1 0 3868 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_24
timestamp 1625156677
transform -1 0 3892 0 1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_8
timestamp 1625156677
transform -1 0 3924 0 1 305
box -2 -3 34 103
use FILL  FILL_3_7_0
timestamp 1625156677
transform -1 0 3932 0 1 305
box -2 -3 10 103
use FILL  FILL_3_7_1
timestamp 1625156677
transform -1 0 3940 0 1 305
box -2 -3 10 103
use NOR3X1  NOR3X1_25
timestamp 1625156677
transform -1 0 4004 0 1 305
box -2 -3 66 103
use OAI21X1  OAI21X1_8
timestamp 1625156677
transform -1 0 4036 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_18
timestamp 1625156677
transform 1 0 4036 0 1 305
box -2 -3 26 103
use AND2X2  AND2X2_2
timestamp 1625156677
transform -1 0 4092 0 1 305
box -2 -3 34 103
use INVX1  INVX1_11
timestamp 1625156677
transform -1 0 4108 0 1 305
box -2 -3 18 103
use XOR2X1  XOR2X1_310
timestamp 1625156677
transform -1 0 4164 0 1 305
box -2 -3 58 103
use XOR2X1  XOR2X1_7
timestamp 1625156677
transform -1 0 4220 0 1 305
box -2 -3 58 103
use XOR2X1  XOR2X1_315
timestamp 1625156677
transform -1 0 4276 0 1 305
box -2 -3 58 103
use XNOR2X1  XNOR2X1_10
timestamp 1625156677
transform -1 0 4332 0 1 305
box -2 -3 58 103
use XOR2X1  XOR2X1_317
timestamp 1625156677
transform 1 0 4332 0 1 305
box -2 -3 58 103
use INVX2  INVX2_92
timestamp 1625156677
transform -1 0 4404 0 1 305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_254
timestamp 1625156677
transform 1 0 4404 0 1 305
box -2 -3 58 103
use FILL  FILL_3_8_0
timestamp 1625156677
transform 1 0 4460 0 1 305
box -2 -3 10 103
use FILL  FILL_3_8_1
timestamp 1625156677
transform 1 0 4468 0 1 305
box -2 -3 10 103
use NAND3X1  NAND3X1_548
timestamp 1625156677
transform 1 0 4476 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_639
timestamp 1625156677
transform -1 0 4540 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_708
timestamp 1625156677
transform -1 0 4564 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_709
timestamp 1625156677
transform 1 0 4564 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_644
timestamp 1625156677
transform 1 0 4588 0 1 305
box -2 -3 34 103
use INVX1  INVX1_598
timestamp 1625156677
transform 1 0 4620 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_403
timestamp 1625156677
transform 1 0 4636 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_448
timestamp 1625156677
transform 1 0 4668 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_405
timestamp 1625156677
transform 1 0 4692 0 1 305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_256
timestamp 1625156677
transform 1 0 4724 0 1 305
box -2 -3 58 103
use OAI21X1  OAI21X1_645
timestamp 1625156677
transform 1 0 4780 0 1 305
box -2 -3 34 103
use AND2X2  AND2X2_197
timestamp 1625156677
transform -1 0 4844 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_713
timestamp 1625156677
transform 1 0 4844 0 1 305
box -2 -3 26 103
use OR2X2  OR2X2_158
timestamp 1625156677
transform 1 0 4868 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_542
timestamp 1625156677
transform -1 0 4932 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_541
timestamp 1625156677
transform -1 0 4964 0 1 305
box -2 -3 34 103
use FILL  FILL_3_9_0
timestamp 1625156677
transform 1 0 4964 0 1 305
box -2 -3 10 103
use FILL  FILL_3_9_1
timestamp 1625156677
transform 1 0 4972 0 1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_399
timestamp 1625156677
transform 1 0 4980 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_711
timestamp 1625156677
transform 1 0 5012 0 1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_539
timestamp 1625156677
transform -1 0 5068 0 1 305
box -2 -3 34 103
use INVX1  INVX1_593
timestamp 1625156677
transform -1 0 5084 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_643
timestamp 1625156677
transform -1 0 5116 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_449
timestamp 1625156677
transform -1 0 5140 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_642
timestamp 1625156677
transform 1 0 5140 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1625156677
transform -1 0 5268 0 1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_134
timestamp 1625156677
transform 1 0 5268 0 1 305
box -2 -3 34 103
use FILL  FILL_4_1
timestamp 1625156677
transform 1 0 5300 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1625156677
transform 1 0 5308 0 1 305
box -2 -3 10 103
use BUFX2  BUFX2_249
timestamp 1625156677
transform -1 0 28 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_42
timestamp 1625156677
transform -1 0 60 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_60
timestamp 1625156677
transform 1 0 60 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_44
timestamp 1625156677
transform -1 0 116 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_45
timestamp 1625156677
transform 1 0 116 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_45
timestamp 1625156677
transform -1 0 180 0 -1 305
box -2 -3 34 103
use NOR3X1  NOR3X1_30
timestamp 1625156677
transform -1 0 244 0 -1 305
box -2 -3 66 103
use OAI21X1  OAI21X1_44
timestamp 1625156677
transform -1 0 276 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_34
timestamp 1625156677
transform -1 0 292 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_61
timestamp 1625156677
transform 1 0 292 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_35
timestamp 1625156677
transform -1 0 348 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_0_0
timestamp 1625156677
transform 1 0 348 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1625156677
transform 1 0 356 0 -1 305
box -2 -3 10 103
use NAND3X1  NAND3X1_43
timestamp 1625156677
transform 1 0 364 0 -1 305
box -2 -3 34 103
use OR2X2  OR2X2_18
timestamp 1625156677
transform -1 0 428 0 -1 305
box -2 -3 34 103
use XOR2X1  XOR2X1_12
timestamp 1625156677
transform -1 0 484 0 -1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_141
timestamp 1625156677
transform 1 0 484 0 -1 305
box -2 -3 98 103
use XOR2X1  XOR2X1_36
timestamp 1625156677
transform 1 0 580 0 -1 305
box -2 -3 58 103
use NAND3X1  NAND3X1_51
timestamp 1625156677
transform -1 0 668 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_50
timestamp 1625156677
transform -1 0 700 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_40
timestamp 1625156677
transform 1 0 700 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_48
timestamp 1625156677
transform -1 0 764 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_36
timestamp 1625156677
transform 1 0 764 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_50
timestamp 1625156677
transform -1 0 812 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_49
timestamp 1625156677
transform 1 0 812 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1625156677
transform -1 0 852 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1625156677
transform -1 0 860 0 -1 305
box -2 -3 10 103
use XOR2X1  XOR2X1_14
timestamp 1625156677
transform -1 0 916 0 -1 305
box -2 -3 58 103
use NAND3X1  NAND3X1_53
timestamp 1625156677
transform 1 0 916 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_53
timestamp 1625156677
transform -1 0 980 0 -1 305
box -2 -3 34 103
use AND2X2  AND2X2_19
timestamp 1625156677
transform -1 0 1012 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_44
timestamp 1625156677
transform 1 0 1012 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_54
timestamp 1625156677
transform 1 0 1036 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_37
timestamp 1625156677
transform -1 0 1084 0 -1 305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_36
timestamp 1625156677
transform 1 0 1084 0 -1 305
box -2 -3 58 103
use XOR2X1  XOR2X1_38
timestamp 1625156677
transform 1 0 1140 0 -1 305
box -2 -3 58 103
use INVX1  INVX1_51
timestamp 1625156677
transform -1 0 1212 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_74
timestamp 1625156677
transform -1 0 1244 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_76
timestamp 1625156677
transform -1 0 1276 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_73
timestamp 1625156677
transform 1 0 1276 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_22
timestamp 1625156677
transform -1 0 1324 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_69
timestamp 1625156677
transform -1 0 1356 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_86
timestamp 1625156677
transform 1 0 1356 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_2_0
timestamp 1625156677
transform 1 0 1380 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1625156677
transform 1 0 1388 0 -1 305
box -2 -3 10 103
use AND2X2  AND2X2_24
timestamp 1625156677
transform 1 0 1396 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_53
timestamp 1625156677
transform -1 0 1460 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_88
timestamp 1625156677
transform -1 0 1484 0 -1 305
box -2 -3 26 103
use XOR2X1  XOR2X1_22
timestamp 1625156677
transform 1 0 1484 0 -1 305
box -2 -3 58 103
use NAND3X1  NAND3X1_64
timestamp 1625156677
transform -1 0 1572 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_50
timestamp 1625156677
transform 1 0 1572 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_48
timestamp 1625156677
transform 1 0 1604 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_65
timestamp 1625156677
transform -1 0 1668 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_46
timestamp 1625156677
transform -1 0 1684 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_64
timestamp 1625156677
transform -1 0 1716 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_49
timestamp 1625156677
transform 1 0 1716 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_65
timestamp 1625156677
transform -1 0 1780 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_50
timestamp 1625156677
transform 1 0 1780 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_83
timestamp 1625156677
transform -1 0 1828 0 -1 305
box -2 -3 26 103
use AND2X2  AND2X2_22
timestamp 1625156677
transform -1 0 1860 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_197
timestamp 1625156677
transform -1 0 1884 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_3_0
timestamp 1625156677
transform 1 0 1884 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1625156677
transform 1 0 1892 0 -1 305
box -2 -3 10 103
use XOR2X1  XOR2X1_24
timestamp 1625156677
transform 1 0 1900 0 -1 305
box -2 -3 58 103
use OR2X2  OR2X2_26
timestamp 1625156677
transform 1 0 1956 0 -1 305
box -2 -3 34 103
use AND2X2  AND2X2_21
timestamp 1625156677
transform 1 0 1988 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_80
timestamp 1625156677
transform 1 0 2020 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_49
timestamp 1625156677
transform -1 0 2068 0 -1 305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_30
timestamp 1625156677
transform 1 0 2068 0 -1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_145
timestamp 1625156677
transform 1 0 2124 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_172
timestamp 1625156677
transform 1 0 2220 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_173
timestamp 1625156677
transform 1 0 2316 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_4_0
timestamp 1625156677
transform 1 0 2412 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_4_1
timestamp 1625156677
transform 1 0 2420 0 -1 305
box -2 -3 10 103
use AND2X2  AND2X2_39
timestamp 1625156677
transform 1 0 2428 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_79
timestamp 1625156677
transform -1 0 2484 0 -1 305
box -2 -3 26 103
use NOR3X1  NOR3X1_38
timestamp 1625156677
transform -1 0 2548 0 -1 305
box -2 -3 66 103
use OAI21X1  OAI21X1_112
timestamp 1625156677
transform 1 0 2548 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_78
timestamp 1625156677
transform -1 0 2596 0 -1 305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_13
timestamp 1625156677
transform 1 0 2596 0 -1 305
box -2 -3 58 103
use XOR2X1  XOR2X1_2
timestamp 1625156677
transform -1 0 2708 0 -1 305
box -2 -3 58 103
use INVX2  INVX2_14
timestamp 1625156677
transform -1 0 2724 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_137
timestamp 1625156677
transform -1 0 2748 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_25
timestamp 1625156677
transform -1 0 2780 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_23
timestamp 1625156677
transform -1 0 2812 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_42
timestamp 1625156677
transform 1 0 2812 0 -1 305
box -2 -3 26 103
use OR2X2  OR2X2_10
timestamp 1625156677
transform -1 0 2868 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_23
timestamp 1625156677
transform 1 0 2868 0 -1 305
box -2 -3 18 103
use NAND3X1  NAND3X1_28
timestamp 1625156677
transform -1 0 2916 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_5_0
timestamp 1625156677
transform -1 0 2924 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_5_1
timestamp 1625156677
transform -1 0 2932 0 -1 305
box -2 -3 10 103
use NAND3X1  NAND3X1_29
timestamp 1625156677
transform -1 0 2964 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_24
timestamp 1625156677
transform -1 0 2980 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_30
timestamp 1625156677
transform -1 0 3012 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_31
timestamp 1625156677
transform -1 0 3044 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_30
timestamp 1625156677
transform 1 0 3044 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_26
timestamp 1625156677
transform -1 0 3100 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_45
timestamp 1625156677
transform -1 0 3124 0 -1 305
box -2 -3 26 103
use OR2X2  OR2X2_11
timestamp 1625156677
transform -1 0 3156 0 -1 305
box -2 -3 34 103
use XOR2X1  XOR2X1_4
timestamp 1625156677
transform -1 0 3212 0 -1 305
box -2 -3 58 103
use NAND3X1  NAND3X1_33
timestamp 1625156677
transform -1 0 3244 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_25
timestamp 1625156677
transform 1 0 3244 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_33
timestamp 1625156677
transform -1 0 3292 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_32
timestamp 1625156677
transform 1 0 3292 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_32
timestamp 1625156677
transform 1 0 3316 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_31
timestamp 1625156677
transform 1 0 3348 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_30
timestamp 1625156677
transform 1 0 3380 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_6_0
timestamp 1625156677
transform 1 0 3412 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_6_1
timestamp 1625156677
transform 1 0 3420 0 -1 305
box -2 -3 10 103
use NAND3X1  NAND3X1_32
timestamp 1625156677
transform 1 0 3428 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_28
timestamp 1625156677
transform 1 0 3460 0 -1 305
box -2 -3 34 103
use OR2X2  OR2X2_12
timestamp 1625156677
transform -1 0 3524 0 -1 305
box -2 -3 34 103
use XOR2X1  XOR2X1_19
timestamp 1625156677
transform -1 0 3580 0 -1 305
box -2 -3 58 103
use INVX1  INVX1_20
timestamp 1625156677
transform 1 0 3580 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_24
timestamp 1625156677
transform 1 0 3596 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_38
timestamp 1625156677
transform -1 0 3652 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_21
timestamp 1625156677
transform -1 0 3668 0 -1 305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_5
timestamp 1625156677
transform 1 0 3668 0 -1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_20
timestamp 1625156677
transform -1 0 3748 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1625156677
transform 1 0 3748 0 -1 305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_4
timestamp 1625156677
transform 1 0 3780 0 -1 305
box -2 -3 58 103
use XOR2X1  XOR2X1_309
timestamp 1625156677
transform 1 0 3836 0 -1 305
box -2 -3 58 103
use BUFX2  BUFX2_154
timestamp 1625156677
transform -1 0 3916 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_7_0
timestamp 1625156677
transform -1 0 3924 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_7_1
timestamp 1625156677
transform -1 0 3932 0 -1 305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_16
timestamp 1625156677
transform -1 0 4004 0 -1 305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1625156677
transform -1 0 4100 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_21
timestamp 1625156677
transform 1 0 4100 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_5
timestamp 1625156677
transform 1 0 4124 0 -1 305
box -2 -3 34 103
use OR2X2  OR2X2_1
timestamp 1625156677
transform -1 0 4188 0 -1 305
box -2 -3 34 103
use XOR2X1  XOR2X1_6
timestamp 1625156677
transform -1 0 4244 0 -1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_34
timestamp 1625156677
transform -1 0 4268 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_33
timestamp 1625156677
transform -1 0 4292 0 -1 305
box -2 -3 26 103
use OR2X2  OR2X2_7
timestamp 1625156677
transform 1 0 4292 0 -1 305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_12
timestamp 1625156677
transform -1 0 4380 0 -1 305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1625156677
transform -1 0 4476 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_8_0
timestamp 1625156677
transform 1 0 4476 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_8_1
timestamp 1625156677
transform 1 0 4484 0 -1 305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_5
timestamp 1625156677
transform 1 0 4492 0 -1 305
box -2 -3 74 103
use BUFX2  BUFX2_118
timestamp 1625156677
transform -1 0 4588 0 -1 305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_255
timestamp 1625156677
transform 1 0 4588 0 -1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_712
timestamp 1625156677
transform 1 0 4644 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_547
timestamp 1625156677
transform -1 0 4700 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_648
timestamp 1625156677
transform 1 0 4700 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_721
timestamp 1625156677
transform -1 0 4756 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_650
timestamp 1625156677
transform 1 0 4756 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_94
timestamp 1625156677
transform 1 0 4788 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_649
timestamp 1625156677
transform 1 0 4804 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_595
timestamp 1625156677
transform 1 0 4836 0 -1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_452
timestamp 1625156677
transform -1 0 4876 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_400
timestamp 1625156677
transform -1 0 4908 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_715
timestamp 1625156677
transform -1 0 4932 0 -1 305
box -2 -3 26 103
use OR2X2  OR2X2_160
timestamp 1625156677
transform -1 0 4964 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_9_0
timestamp 1625156677
transform -1 0 4972 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_9_1
timestamp 1625156677
transform -1 0 4980 0 -1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_401
timestamp 1625156677
transform -1 0 5012 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_546
timestamp 1625156677
transform -1 0 5044 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_716
timestamp 1625156677
transform -1 0 5068 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_544
timestamp 1625156677
transform 1 0 5068 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_646
timestamp 1625156677
transform -1 0 5132 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_647
timestamp 1625156677
transform -1 0 5164 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_451
timestamp 1625156677
transform 1 0 5164 0 -1 305
box -2 -3 26 103
use AND2X2  AND2X2_196
timestamp 1625156677
transform -1 0 5220 0 -1 305
box -2 -3 34 103
use AND2X2  AND2X2_198
timestamp 1625156677
transform -1 0 5252 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_122
timestamp 1625156677
transform -1 0 5276 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_190
timestamp 1625156677
transform -1 0 5308 0 -1 305
box -2 -3 34 103
use FILL  FILL_3_1
timestamp 1625156677
transform -1 0 5316 0 -1 305
box -2 -3 10 103
use BUFX2  BUFX2_147
timestamp 1625156677
transform 1 0 4 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_131
timestamp 1625156677
transform 1 0 28 0 1 105
box -2 -3 26 103
use OR2X2  OR2X2_17
timestamp 1625156677
transform 1 0 52 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_41
timestamp 1625156677
transform -1 0 116 0 1 105
box -2 -3 34 103
use INVX1  INVX1_33
timestamp 1625156677
transform 1 0 116 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_42
timestamp 1625156677
transform -1 0 164 0 1 105
box -2 -3 34 103
use NOR3X1  NOR3X1_29
timestamp 1625156677
transform 1 0 164 0 1 105
box -2 -3 66 103
use NAND2X1  NAND2X1_63
timestamp 1625156677
transform -1 0 252 0 1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_25
timestamp 1625156677
transform -1 0 308 0 1 105
box -2 -3 58 103
use NAND2X1  NAND2X1_62
timestamp 1625156677
transform 1 0 308 0 1 105
box -2 -3 26 103
use FILL  FILL_1_0_0
timestamp 1625156677
transform -1 0 340 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1625156677
transform -1 0 348 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_43
timestamp 1625156677
transform -1 0 380 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_43
timestamp 1625156677
transform 1 0 380 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_39
timestamp 1625156677
transform 1 0 404 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_57
timestamp 1625156677
transform 1 0 436 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_36
timestamp 1625156677
transform -1 0 500 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_37
timestamp 1625156677
transform -1 0 532 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_46
timestamp 1625156677
transform -1 0 564 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_47
timestamp 1625156677
transform -1 0 596 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_38
timestamp 1625156677
transform 1 0 596 0 1 105
box -2 -3 34 103
use INVX1  INVX1_35
timestamp 1625156677
transform 1 0 628 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_48
timestamp 1625156677
transform -1 0 676 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_47
timestamp 1625156677
transform 1 0 676 0 1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_26
timestamp 1625156677
transform 1 0 708 0 1 105
box -2 -3 58 103
use AND2X2  AND2X2_18
timestamp 1625156677
transform -1 0 796 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_49
timestamp 1625156677
transform 1 0 796 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_67
timestamp 1625156677
transform -1 0 852 0 1 105
box -2 -3 26 103
use FILL  FILL_1_1_0
timestamp 1625156677
transform -1 0 860 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1625156677
transform -1 0 868 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_41
timestamp 1625156677
transform -1 0 900 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_69
timestamp 1625156677
transform -1 0 924 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_42
timestamp 1625156677
transform -1 0 956 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_45
timestamp 1625156677
transform 1 0 956 0 1 105
box -2 -3 26 103
use INVX1  INVX1_38
timestamp 1625156677
transform -1 0 996 0 1 105
box -2 -3 18 103
use OR2X2  OR2X2_22
timestamp 1625156677
transform -1 0 1028 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_55
timestamp 1625156677
transform -1 0 1060 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_70
timestamp 1625156677
transform 1 0 1060 0 1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_52
timestamp 1625156677
transform 1 0 1084 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_54
timestamp 1625156677
transform 1 0 1116 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_47
timestamp 1625156677
transform -1 0 1172 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_68
timestamp 1625156677
transform -1 0 1196 0 1 105
box -2 -3 26 103
use OR2X2  OR2X2_21
timestamp 1625156677
transform -1 0 1228 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_161
timestamp 1625156677
transform -1 0 1324 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_241
timestamp 1625156677
transform 1 0 1324 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_195
timestamp 1625156677
transform 1 0 1348 0 1 105
box -2 -3 26 103
use FILL  FILL_1_2_0
timestamp 1625156677
transform -1 0 1380 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1625156677
transform -1 0 1388 0 1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_93
timestamp 1625156677
transform -1 0 1412 0 1 105
box -2 -3 26 103
use OR2X2  OR2X2_32
timestamp 1625156677
transform -1 0 1444 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_92
timestamp 1625156677
transform -1 0 1468 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_55
timestamp 1625156677
transform -1 0 1492 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_54
timestamp 1625156677
transform -1 0 1524 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_73
timestamp 1625156677
transform -1 0 1556 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_89
timestamp 1625156677
transform -1 0 1580 0 1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_69
timestamp 1625156677
transform -1 0 1612 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_67
timestamp 1625156677
transform 1 0 1612 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_71
timestamp 1625156677
transform 1 0 1644 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_72
timestamp 1625156677
transform -1 0 1708 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_70
timestamp 1625156677
transform -1 0 1740 0 1 105
box -2 -3 34 103
use INVX1  INVX1_48
timestamp 1625156677
transform 1 0 1740 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_71
timestamp 1625156677
transform -1 0 1788 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_70
timestamp 1625156677
transform -1 0 1820 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_54
timestamp 1625156677
transform 1 0 1820 0 1 105
box -2 -3 26 103
use AND2X2  AND2X2_25
timestamp 1625156677
transform -1 0 1876 0 1 105
box -2 -3 34 103
use FILL  FILL_1_3_0
timestamp 1625156677
transform -1 0 1884 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_1
timestamp 1625156677
transform -1 0 1892 0 1 105
box -2 -3 10 103
use OR2X2  OR2X2_29
timestamp 1625156677
transform -1 0 1924 0 1 105
box -2 -3 34 103
use OR2X2  OR2X2_27
timestamp 1625156677
transform -1 0 1956 0 1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_25
timestamp 1625156677
transform 1 0 1956 0 1 105
box -2 -3 58 103
use BUFX2  BUFX2_117
timestamp 1625156677
transform 1 0 2012 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_91
timestamp 1625156677
transform -1 0 2060 0 1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_39
timestamp 1625156677
transform -1 0 2116 0 1 105
box -2 -3 58 103
use NAND2X1  NAND2X1_72
timestamp 1625156677
transform -1 0 2140 0 1 105
box -2 -3 26 103
use OR2X2  OR2X2_23
timestamp 1625156677
transform -1 0 2172 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_71
timestamp 1625156677
transform -1 0 2196 0 1 105
box -2 -3 26 103
use INVX1  INVX1_39
timestamp 1625156677
transform -1 0 2212 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_144
timestamp 1625156677
transform -1 0 2308 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_239
timestamp 1625156677
transform -1 0 2332 0 1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_38
timestamp 1625156677
transform 1 0 2332 0 1 105
box -2 -3 58 103
use FILL  FILL_1_4_0
timestamp 1625156677
transform 1 0 2388 0 1 105
box -2 -3 10 103
use FILL  FILL_1_4_1
timestamp 1625156677
transform 1 0 2396 0 1 105
box -2 -3 10 103
use BUFX2  BUFX2_86
timestamp 1625156677
transform 1 0 2404 0 1 105
box -2 -3 26 103
use XOR2X1  XOR2X1_26
timestamp 1625156677
transform -1 0 2484 0 1 105
box -2 -3 58 103
use XOR2X1  XOR2X1_28
timestamp 1625156677
transform -1 0 2540 0 1 105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_14
timestamp 1625156677
transform 1 0 2540 0 1 105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_15
timestamp 1625156677
transform 1 0 2596 0 1 105
box -2 -3 58 103
use NAND2X1  NAND2X1_39
timestamp 1625156677
transform -1 0 2676 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_33
timestamp 1625156677
transform 1 0 2676 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_26
timestamp 1625156677
transform -1 0 2740 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_43
timestamp 1625156677
transform 1 0 2740 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_26
timestamp 1625156677
transform -1 0 2796 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_28
timestamp 1625156677
transform -1 0 2828 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_33
timestamp 1625156677
transform 1 0 2828 0 1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_27
timestamp 1625156677
transform -1 0 2884 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_27
timestamp 1625156677
transform 1 0 2884 0 1 105
box -2 -3 34 103
use FILL  FILL_1_5_0
timestamp 1625156677
transform -1 0 2924 0 1 105
box -2 -3 10 103
use FILL  FILL_1_5_1
timestamp 1625156677
transform -1 0 2932 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_24
timestamp 1625156677
transform -1 0 2964 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_44
timestamp 1625156677
transform -1 0 2988 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_25
timestamp 1625156677
transform -1 0 3020 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_27
timestamp 1625156677
transform -1 0 3052 0 1 105
box -2 -3 34 103
use NOR3X1  NOR3X1_28
timestamp 1625156677
transform 1 0 3052 0 1 105
box -2 -3 66 103
use NOR2X1  NOR2X1_29
timestamp 1625156677
transform 1 0 3116 0 1 105
box -2 -3 26 103
use AND2X2  AND2X2_9
timestamp 1625156677
transform -1 0 3172 0 1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_17
timestamp 1625156677
transform 1 0 3172 0 1 105
box -2 -3 58 103
use NOR2X1  NOR2X1_37
timestamp 1625156677
transform -1 0 3252 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_36
timestamp 1625156677
transform 1 0 3252 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_38
timestamp 1625156677
transform -1 0 3308 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_56
timestamp 1625156677
transform -1 0 3332 0 1 105
box -2 -3 26 103
use AND2X2  AND2X2_12
timestamp 1625156677
transform -1 0 3364 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_48
timestamp 1625156677
transform -1 0 3388 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_29
timestamp 1625156677
transform -1 0 3420 0 1 105
box -2 -3 34 103
use FILL  FILL_1_6_0
timestamp 1625156677
transform 1 0 3420 0 1 105
box -2 -3 10 103
use FILL  FILL_1_6_1
timestamp 1625156677
transform 1 0 3428 0 1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_50
timestamp 1625156677
transform 1 0 3436 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_30
timestamp 1625156677
transform -1 0 3492 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_35
timestamp 1625156677
transform 1 0 3492 0 1 105
box -2 -3 26 103
use INVX1  INVX1_27
timestamp 1625156677
transform -1 0 3532 0 1 105
box -2 -3 18 103
use OR2X2  OR2X2_14
timestamp 1625156677
transform 1 0 3532 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_37
timestamp 1625156677
transform -1 0 3596 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1625156677
transform -1 0 3620 0 1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_35
timestamp 1625156677
transform 1 0 3620 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_37
timestamp 1625156677
transform -1 0 3684 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_36
timestamp 1625156677
transform 1 0 3684 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_34
timestamp 1625156677
transform 1 0 3716 0 1 105
box -2 -3 26 103
use INVX1  INVX1_26
timestamp 1625156677
transform 1 0 3740 0 1 105
box -2 -3 18 103
use INVX2  INVX2_11
timestamp 1625156677
transform -1 0 3772 0 1 105
box -2 -3 18 103
use NAND3X1  NAND3X1_34
timestamp 1625156677
transform 1 0 3772 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_36
timestamp 1625156677
transform -1 0 3836 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_135
timestamp 1625156677
transform -1 0 3932 0 1 105
box -2 -3 98 103
use FILL  FILL_1_7_0
timestamp 1625156677
transform -1 0 3940 0 1 105
box -2 -3 10 103
use FILL  FILL_1_7_1
timestamp 1625156677
transform -1 0 3948 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1625156677
transform -1 0 4044 0 1 105
box -2 -3 98 103
use BUFX2  BUFX2_128
timestamp 1625156677
transform 1 0 4044 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_137
timestamp 1625156677
transform 1 0 4068 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1625156677
transform -1 0 4260 0 1 105
box -2 -3 98 103
use XOR2X1  XOR2X1_21
timestamp 1625156677
transform -1 0 4316 0 1 105
box -2 -3 58 103
use BUFX2  BUFX2_153
timestamp 1625156677
transform -1 0 4340 0 1 105
box -2 -3 26 103
use INVX1  INVX1_17
timestamp 1625156677
transform -1 0 4356 0 1 105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_19
timestamp 1625156677
transform 1 0 4356 0 1 105
box -2 -3 58 103
use XOR2X1  XOR2X1_316
timestamp 1625156677
transform 1 0 4412 0 1 105
box -2 -3 58 103
use FILL  FILL_1_8_0
timestamp 1625156677
transform -1 0 4476 0 1 105
box -2 -3 10 103
use FILL  FILL_1_8_1
timestamp 1625156677
transform -1 0 4484 0 1 105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_11
timestamp 1625156677
transform -1 0 4540 0 1 105
box -2 -3 58 103
use XOR2X1  XOR2X1_9
timestamp 1625156677
transform -1 0 4596 0 1 105
box -2 -3 58 103
use XOR2X1  XOR2X1_8
timestamp 1625156677
transform -1 0 4652 0 1 105
box -2 -3 58 103
use BUFX2  BUFX2_129
timestamp 1625156677
transform 1 0 4652 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_454
timestamp 1625156677
transform -1 0 4700 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_453
timestamp 1625156677
transform -1 0 4724 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_402
timestamp 1625156677
transform 1 0 4724 0 1 105
box -2 -3 34 103
use INVX1  INVX1_597
timestamp 1625156677
transform 1 0 4756 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_722
timestamp 1625156677
transform -1 0 4796 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_651
timestamp 1625156677
transform 1 0 4796 0 1 105
box -2 -3 34 103
use INVX1  INVX1_600
timestamp 1625156677
transform -1 0 4844 0 1 105
box -2 -3 18 103
use NAND3X1  NAND3X1_549
timestamp 1625156677
transform -1 0 4876 0 1 105
box -2 -3 34 103
use INVX1  INVX1_599
timestamp 1625156677
transform -1 0 4892 0 1 105
box -2 -3 18 103
use BUFX2  BUFX2_28
timestamp 1625156677
transform 1 0 4892 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_720
timestamp 1625156677
transform -1 0 4940 0 1 105
box -2 -3 26 103
use FILL  FILL_1_9_0
timestamp 1625156677
transform -1 0 4948 0 1 105
box -2 -3 10 103
use FILL  FILL_1_9_1
timestamp 1625156677
transform -1 0 4956 0 1 105
box -2 -3 10 103
use OR2X2  OR2X2_162
timestamp 1625156677
transform -1 0 4988 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_719
timestamp 1625156677
transform -1 0 5012 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_46
timestamp 1625156677
transform -1 0 5036 0 1 105
box -2 -3 26 103
use OR2X2  OR2X2_159
timestamp 1625156677
transform 1 0 5036 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_545
timestamp 1625156677
transform -1 0 5100 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_543
timestamp 1625156677
transform -1 0 5132 0 1 105
box -2 -3 34 103
use INVX1  INVX1_594
timestamp 1625156677
transform -1 0 5148 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_714
timestamp 1625156677
transform -1 0 5172 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1625156677
transform -1 0 5268 0 1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_216
timestamp 1625156677
transform -1 0 5292 0 1 105
box -2 -3 26 103
use FILL  FILL_2_1
timestamp 1625156677
transform 1 0 5292 0 1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1625156677
transform 1 0 5300 0 1 105
box -2 -3 10 103
use FILL  FILL_2_3
timestamp 1625156677
transform 1 0 5308 0 1 105
box -2 -3 10 103
use BUFX2  BUFX2_85
timestamp 1625156677
transform -1 0 28 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_59
timestamp 1625156677
transform 1 0 28 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_47
timestamp 1625156677
transform -1 0 76 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_59
timestamp 1625156677
transform 1 0 76 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_141
timestamp 1625156677
transform 1 0 100 0 -1 105
box -2 -3 26 103
use AND2X2  AND2X2_14
timestamp 1625156677
transform 1 0 124 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_38
timestamp 1625156677
transform -1 0 180 0 -1 105
box -2 -3 26 103
use XOR2X1  XOR2X1_13
timestamp 1625156677
transform -1 0 236 0 -1 105
box -2 -3 58 103
use OAI21X1  OAI21X1_46
timestamp 1625156677
transform 1 0 236 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_51
timestamp 1625156677
transform 1 0 268 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_41
timestamp 1625156677
transform 1 0 300 0 -1 105
box -2 -3 18 103
use XOR2X1  XOR2X1_30
timestamp 1625156677
transform 1 0 316 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_0_0
timestamp 1625156677
transform 1 0 372 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1625156677
transform 1 0 380 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_250
timestamp 1625156677
transform 1 0 388 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_44
timestamp 1625156677
transform 1 0 412 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_41
timestamp 1625156677
transform 1 0 444 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_18
timestamp 1625156677
transform 1 0 468 0 -1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_46
timestamp 1625156677
transform 1 0 484 0 -1 105
box -2 -3 34 103
use OR2X2  OR2X2_19
timestamp 1625156677
transform 1 0 516 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_64
timestamp 1625156677
transform 1 0 548 0 -1 105
box -2 -3 26 103
use AND2X2  AND2X2_16
timestamp 1625156677
transform 1 0 572 0 -1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_15
timestamp 1625156677
transform -1 0 660 0 -1 105
box -2 -3 58 103
use NOR2X1  NOR2X1_40
timestamp 1625156677
transform -1 0 684 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_66
timestamp 1625156677
transform 1 0 684 0 -1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_56
timestamp 1625156677
transform 1 0 708 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_75
timestamp 1625156677
transform -1 0 764 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_55
timestamp 1625156677
transform 1 0 764 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_52
timestamp 1625156677
transform 1 0 796 0 -1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_27
timestamp 1625156677
transform 1 0 828 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_1_0
timestamp 1625156677
transform 1 0 884 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1625156677
transform 1 0 892 0 -1 105
box -2 -3 10 103
use INVX2  INVX2_19
timestamp 1625156677
transform 1 0 900 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_56
timestamp 1625156677
transform 1 0 916 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_57
timestamp 1625156677
transform 1 0 948 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_43
timestamp 1625156677
transform 1 0 980 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_40
timestamp 1625156677
transform -1 0 1028 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_46
timestamp 1625156677
transform 1 0 1028 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_74
timestamp 1625156677
transform 1 0 1052 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_73
timestamp 1625156677
transform 1 0 1076 0 -1 105
box -2 -3 26 103
use OR2X2  OR2X2_24
timestamp 1625156677
transform -1 0 1132 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_58
timestamp 1625156677
transform -1 0 1164 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_42
timestamp 1625156677
transform 1 0 1164 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_58
timestamp 1625156677
transform 1 0 1180 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_43
timestamp 1625156677
transform -1 0 1228 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_76
timestamp 1625156677
transform 1 0 1228 0 -1 105
box -2 -3 26 103
use XOR2X1  XOR2X1_51
timestamp 1625156677
transform -1 0 1308 0 -1 105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_47
timestamp 1625156677
transform 1 0 1308 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_2_0
timestamp 1625156677
transform 1 0 1364 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1625156677
transform 1 0 1372 0 -1 105
box -2 -3 10 103
use XOR2X1  XOR2X1_39
timestamp 1625156677
transform 1 0 1380 0 -1 105
box -2 -3 58 103
use BUFX2  BUFX2_196
timestamp 1625156677
transform 1 0 1436 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_49
timestamp 1625156677
transform -1 0 1476 0 -1 105
box -2 -3 18 103
use BUFX2  BUFX2_242
timestamp 1625156677
transform 1 0 1476 0 -1 105
box -2 -3 26 103
use OR2X2  OR2X2_30
timestamp 1625156677
transform -1 0 1532 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_52
timestamp 1625156677
transform -1 0 1564 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_68
timestamp 1625156677
transform -1 0 1596 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_66
timestamp 1625156677
transform -1 0 1628 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_84
timestamp 1625156677
transform 1 0 1628 0 -1 105
box -2 -3 26 103
use OR2X2  OR2X2_28
timestamp 1625156677
transform -1 0 1684 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_47
timestamp 1625156677
transform 1 0 1684 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_67
timestamp 1625156677
transform -1 0 1732 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_66
timestamp 1625156677
transform -1 0 1764 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_52
timestamp 1625156677
transform 1 0 1764 0 -1 105
box -2 -3 26 103
use AND2X2  AND2X2_23
timestamp 1625156677
transform -1 0 1820 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_87
timestamp 1625156677
transform 1 0 1820 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_3_0
timestamp 1625156677
transform -1 0 1852 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_1
timestamp 1625156677
transform -1 0 1860 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_151
timestamp 1625156677
transform -1 0 1956 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_150
timestamp 1625156677
transform -1 0 2052 0 -1 105
box -2 -3 98 103
use OR2X2  OR2X2_31
timestamp 1625156677
transform -1 0 2084 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_90
timestamp 1625156677
transform -1 0 2108 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_50
timestamp 1625156677
transform -1 0 2124 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_152
timestamp 1625156677
transform -1 0 2220 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_153
timestamp 1625156677
transform 1 0 2220 0 -1 105
box -2 -3 98 103
use XOR2X1  XOR2X1_41
timestamp 1625156677
transform -1 0 2372 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_4_0
timestamp 1625156677
transform 1 0 2372 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_4_1
timestamp 1625156677
transform 1 0 2380 0 -1 105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_37
timestamp 1625156677
transform 1 0 2388 0 -1 105
box -2 -3 58 103
use XOR2X1  XOR2X1_27
timestamp 1625156677
transform -1 0 2500 0 -1 105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_131
timestamp 1625156677
transform 1 0 2500 0 -1 105
box -2 -3 98 103
use XNOR2X1  XNOR2X1_16
timestamp 1625156677
transform 1 0 2596 0 -1 105
box -2 -3 58 103
use NAND2X1  NAND2X1_40
timestamp 1625156677
transform 1 0 2652 0 -1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_23
timestamp 1625156677
transform 1 0 2676 0 -1 105
box -2 -3 34 103
use OR2X2  OR2X2_9
timestamp 1625156677
transform -1 0 2740 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_41
timestamp 1625156677
transform -1 0 2764 0 -1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_24
timestamp 1625156677
transform -1 0 2796 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_22
timestamp 1625156677
transform 1 0 2796 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_25
timestamp 1625156677
transform -1 0 2844 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_28
timestamp 1625156677
transform -1 0 2868 0 -1 105
box -2 -3 26 103
use NOR3X1  NOR3X1_27
timestamp 1625156677
transform 1 0 2868 0 -1 105
box -2 -3 66 103
use FILL  FILL_0_5_0
timestamp 1625156677
transform -1 0 2940 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_5_1
timestamp 1625156677
transform -1 0 2948 0 -1 105
box -2 -3 10 103
use AND2X2  AND2X2_8
timestamp 1625156677
transform -1 0 2980 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_39
timestamp 1625156677
transform 1 0 2980 0 -1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_20
timestamp 1625156677
transform -1 0 3068 0 -1 105
box -2 -3 58 103
use OAI21X1  OAI21X1_29
timestamp 1625156677
transform -1 0 3100 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_34
timestamp 1625156677
transform 1 0 3100 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_31
timestamp 1625156677
transform -1 0 3156 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_15
timestamp 1625156677
transform 1 0 3156 0 -1 105
box -2 -3 18 103
use INVX1  INVX1_30
timestamp 1625156677
transform 1 0 3172 0 -1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_32
timestamp 1625156677
transform 1 0 3188 0 -1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_3
timestamp 1625156677
transform -1 0 3276 0 -1 105
box -2 -3 58 103
use AOI21X1  AOI21X1_34
timestamp 1625156677
transform 1 0 3276 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_47
timestamp 1625156677
transform -1 0 3332 0 -1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_38
timestamp 1625156677
transform 1 0 3332 0 -1 105
box -2 -3 34 103
use XOR2X1  XOR2X1_29
timestamp 1625156677
transform -1 0 3420 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_6_0
timestamp 1625156677
transform 1 0 3420 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_6_1
timestamp 1625156677
transform 1 0 3428 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_35
timestamp 1625156677
transform 1 0 3436 0 -1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_18
timestamp 1625156677
transform 1 0 3468 0 -1 105
box -2 -3 58 103
use INVX2  INVX2_16
timestamp 1625156677
transform 1 0 3524 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_39
timestamp 1625156677
transform 1 0 3540 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_40
timestamp 1625156677
transform 1 0 3572 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_31
timestamp 1625156677
transform 1 0 3604 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_29
timestamp 1625156677
transform -1 0 3652 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_41
timestamp 1625156677
transform 1 0 3652 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_57
timestamp 1625156677
transform -1 0 3708 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_32
timestamp 1625156677
transform -1 0 3724 0 -1 105
box -2 -3 18 103
use NAND3X1  NAND3X1_40
timestamp 1625156677
transform -1 0 3756 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_31
timestamp 1625156677
transform -1 0 3772 0 -1 105
box -2 -3 18 103
use AND2X2  AND2X2_13
timestamp 1625156677
transform -1 0 3804 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_55
timestamp 1625156677
transform -1 0 3828 0 -1 105
box -2 -3 26 103
use OR2X2  OR2X2_16
timestamp 1625156677
transform -1 0 3860 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_54
timestamp 1625156677
transform 1 0 3860 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_49
timestamp 1625156677
transform -1 0 3908 0 -1 105
box -2 -3 26 103
use OR2X2  OR2X2_13
timestamp 1625156677
transform 1 0 3908 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_7_0
timestamp 1625156677
transform 1 0 3940 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_7_1
timestamp 1625156677
transform 1 0 3948 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_89
timestamp 1625156677
transform 1 0 3956 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1625156677
transform -1 0 4076 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_136
timestamp 1625156677
transform 1 0 4076 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1625156677
transform 1 0 4172 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_28
timestamp 1625156677
transform 1 0 4268 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_53
timestamp 1625156677
transform -1 0 4308 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_52
timestamp 1625156677
transform 1 0 4308 0 -1 105
box -2 -3 26 103
use OR2X2  OR2X2_15
timestamp 1625156677
transform 1 0 4332 0 -1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_21
timestamp 1625156677
transform -1 0 4420 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_8_0
timestamp 1625156677
transform 1 0 4420 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_8_1
timestamp 1625156677
transform 1 0 4428 0 -1 105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_20
timestamp 1625156677
transform 1 0 4436 0 -1 105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1625156677
transform -1 0 4588 0 -1 105
box -2 -3 98 103
use XOR2X1  XOR2X1_11
timestamp 1625156677
transform 1 0 4588 0 -1 105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1625156677
transform 1 0 4644 0 -1 105
box -2 -3 98 103
use XOR2X1  XOR2X1_318
timestamp 1625156677
transform -1 0 4796 0 -1 105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_258
timestamp 1625156677
transform 1 0 4796 0 -1 105
box -2 -3 58 103
use XNOR2X1  XNOR2X1_259
timestamp 1625156677
transform 1 0 4852 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_9_0
timestamp 1625156677
transform -1 0 4916 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_9_1
timestamp 1625156677
transform -1 0 4924 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_129
timestamp 1625156677
transform -1 0 5020 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_718
timestamp 1625156677
transform -1 0 5044 0 -1 105
box -2 -3 26 103
use OR2X2  OR2X2_161
timestamp 1625156677
transform -1 0 5076 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_717
timestamp 1625156677
transform -1 0 5100 0 -1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_257
timestamp 1625156677
transform -1 0 5156 0 -1 105
box -2 -3 58 103
use INVX1  INVX1_596
timestamp 1625156677
transform -1 0 5172 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1625156677
transform -1 0 5268 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_183
timestamp 1625156677
transform -1 0 5300 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_1
timestamp 1625156677
transform -1 0 5308 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1625156677
transform -1 0 5316 0 -1 105
box -2 -3 10 103
<< labels >>
flabel metal6 s 344 -30 360 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 856 -30 872 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 3718 -22 3722 -18 7 FreeSans 24 270 0 0 inicio
port 2 nsew
flabel metal3 s 5342 1658 5346 1662 3 FreeSans 24 0 0 0 bloque_bytes[0]
port 3 nsew
flabel metal3 s 5342 1158 5346 1162 3 FreeSans 24 0 0 0 bloque_bytes[1]
port 4 nsew
flabel metal3 s 5342 1058 5346 1062 3 FreeSans 24 0 0 0 bloque_bytes[2]
port 5 nsew
flabel metal3 s 5342 3648 5346 3652 3 FreeSans 24 90 0 0 bloque_bytes[3]
port 6 nsew
flabel metal3 s 5342 678 5346 682 3 FreeSans 24 0 0 0 bloque_bytes[4]
port 7 nsew
flabel metal3 s 5342 1458 5346 1462 3 FreeSans 24 0 0 0 bloque_bytes[5]
port 8 nsew
flabel metal2 s 1478 -22 1482 -18 7 FreeSans 24 270 0 0 bloque_bytes[6]
port 9 nsew
flabel metal3 s 5342 1078 5346 1082 3 FreeSans 24 0 0 0 bloque_bytes[7]
port 10 nsew
flabel metal2 s 4214 3728 4218 3732 3 FreeSans 24 90 0 0 bloque_bytes[8]
port 11 nsew
flabel metal2 s 4294 3728 4298 3732 3 FreeSans 24 90 0 0 bloque_bytes[9]
port 12 nsew
flabel metal2 s 4374 3728 4378 3732 3 FreeSans 24 90 0 0 bloque_bytes[10]
port 13 nsew
flabel metal3 s 5342 2868 5346 2872 3 FreeSans 24 0 0 0 bloque_bytes[11]
port 14 nsew
flabel metal3 s 5342 2748 5346 2752 3 FreeSans 24 0 0 0 bloque_bytes[12]
port 15 nsew
flabel metal2 s 3998 3728 4002 3732 3 FreeSans 24 90 0 0 bloque_bytes[13]
port 16 nsew
flabel metal2 s 2182 -22 2186 -18 7 FreeSans 24 270 0 0 bloque_bytes[14]
port 17 nsew
flabel metal2 s 1894 -22 1898 -18 7 FreeSans 24 270 0 0 bloque_bytes[15]
port 18 nsew
flabel metal3 s 5342 948 5346 952 3 FreeSans 24 0 0 0 bloque_bytes[16]
port 19 nsew
flabel metal3 s 5342 748 5346 752 3 FreeSans 24 0 0 0 bloque_bytes[17]
port 20 nsew
flabel metal3 s 5342 658 5346 662 3 FreeSans 24 0 0 0 bloque_bytes[18]
port 21 nsew
flabel metal2 s 4486 -22 4490 -18 7 FreeSans 24 270 0 0 bloque_bytes[19]
port 22 nsew
flabel metal3 s 5342 1178 5346 1182 3 FreeSans 24 0 0 0 bloque_bytes[20]
port 23 nsew
flabel metal2 s 4190 -22 4194 -18 7 FreeSans 24 270 0 0 bloque_bytes[21]
port 24 nsew
flabel metal2 s 3558 -22 3562 -18 7 FreeSans 24 270 0 0 bloque_bytes[22]
port 25 nsew
flabel metal2 s 2926 -22 2930 -18 7 FreeSans 24 270 0 0 bloque_bytes[23]
port 26 nsew
flabel metal2 s 2686 3728 2690 3732 3 FreeSans 24 90 0 0 bloque_bytes[24]
port 27 nsew
flabel metal2 s 3286 3728 3290 3732 3 FreeSans 24 90 0 0 bloque_bytes[25]
port 28 nsew
flabel metal2 s 2718 3728 2722 3732 3 FreeSans 24 90 0 0 bloque_bytes[26]
port 29 nsew
flabel metal2 s 1358 -22 1362 -18 7 FreeSans 24 270 0 0 bloque_bytes[27]
port 30 nsew
flabel metal2 s 2206 3728 2210 3732 3 FreeSans 24 90 0 0 bloque_bytes[28]
port 31 nsew
flabel metal2 s 1678 -22 1682 -18 7 FreeSans 24 270 0 0 bloque_bytes[29]
port 32 nsew
flabel metal2 s 2198 -22 2202 -18 7 FreeSans 24 270 0 0 bloque_bytes[30]
port 33 nsew
flabel metal2 s 1798 -22 1802 -18 7 FreeSans 24 270 0 0 bloque_bytes[31]
port 34 nsew
flabel metal2 s 3086 -22 3090 -18 7 FreeSans 24 270 0 0 bloque_bytes[32]
port 35 nsew
flabel metal2 s 2558 -22 2562 -18 7 FreeSans 24 270 0 0 bloque_bytes[33]
port 36 nsew
flabel metal2 s 2278 -22 2282 -18 7 FreeSans 24 270 0 0 bloque_bytes[34]
port 37 nsew
flabel metal2 s 2358 -22 2362 -18 7 FreeSans 24 270 0 0 bloque_bytes[35]
port 38 nsew
flabel metal2 s 2446 -22 2450 -18 7 FreeSans 24 270 0 0 bloque_bytes[36]
port 39 nsew
flabel metal2 s 2262 -22 2266 -18 7 FreeSans 24 270 0 0 bloque_bytes[37]
port 40 nsew
flabel metal2 s 2062 -22 2066 -18 7 FreeSans 24 270 0 0 bloque_bytes[38]
port 41 nsew
flabel metal2 s 2214 -22 2218 -18 7 FreeSans 24 270 0 0 bloque_bytes[39]
port 42 nsew
flabel metal2 s 2046 -22 2050 -18 7 FreeSans 24 270 0 0 bloque_bytes[40]
port 43 nsew
flabel metal2 s 1390 -22 1394 -18 7 FreeSans 24 270 0 0 bloque_bytes[41]
port 44 nsew
flabel metal2 s 1734 -22 1738 -18 7 FreeSans 24 270 0 0 bloque_bytes[42]
port 45 nsew
flabel metal2 s 1254 -22 1258 -18 7 FreeSans 24 270 0 0 bloque_bytes[43]
port 46 nsew
flabel metal3 s -26 878 -22 882 7 FreeSans 24 0 0 0 bloque_bytes[44]
port 47 nsew
flabel metal2 s 1278 -22 1282 -18 7 FreeSans 24 270 0 0 bloque_bytes[45]
port 48 nsew
flabel metal2 s 1462 -22 1466 -18 7 FreeSans 24 270 0 0 bloque_bytes[46]
port 49 nsew
flabel metal2 s 1638 -22 1642 -18 7 FreeSans 24 270 0 0 bloque_bytes[47]
port 50 nsew
flabel metal2 s 798 -22 802 -18 7 FreeSans 24 270 0 0 bloque_bytes[48]
port 51 nsew
flabel metal3 s -26 858 -22 862 7 FreeSans 24 0 0 0 bloque_bytes[49]
port 52 nsew
flabel metal3 s -26 748 -22 752 7 FreeSans 24 0 0 0 bloque_bytes[50]
port 53 nsew
flabel metal3 s -26 548 -22 552 7 FreeSans 24 0 0 0 bloque_bytes[51]
port 54 nsew
flabel metal2 s 558 -22 562 -18 7 FreeSans 24 270 0 0 bloque_bytes[52]
port 55 nsew
flabel metal2 s 1078 -22 1082 -18 7 FreeSans 24 270 0 0 bloque_bytes[53]
port 56 nsew
flabel metal2 s 1230 -22 1234 -18 7 FreeSans 24 270 0 0 bloque_bytes[54]
port 57 nsew
flabel metal2 s 1294 -22 1298 -18 7 FreeSans 24 270 0 0 bloque_bytes[55]
port 58 nsew
flabel metal2 s 2126 -22 2130 -18 7 FreeSans 24 270 0 0 bloque_bytes[56]
port 59 nsew
flabel metal2 s 2078 -22 2082 -18 7 FreeSans 24 270 0 0 bloque_bytes[57]
port 60 nsew
flabel metal2 s 2326 -22 2330 -18 7 FreeSans 24 270 0 0 bloque_bytes[58]
port 61 nsew
flabel metal2 s 2094 -22 2098 -18 7 FreeSans 24 270 0 0 bloque_bytes[59]
port 62 nsew
flabel metal2 s 2006 -22 2010 -18 7 FreeSans 24 270 0 0 bloque_bytes[60]
port 63 nsew
flabel metal2 s 1910 -22 1914 -18 7 FreeSans 24 270 0 0 bloque_bytes[61]
port 64 nsew
flabel metal2 s 2246 -22 2250 -18 7 FreeSans 24 270 0 0 bloque_bytes[62]
port 65 nsew
flabel metal2 s 2310 -22 2314 -18 7 FreeSans 24 270 0 0 bloque_bytes[63]
port 66 nsew
flabel metal3 s -26 348 -22 352 7 FreeSans 24 0 0 0 bloque_bytes[64]
port 67 nsew
flabel metal3 s -26 568 -22 572 7 FreeSans 24 0 0 0 bloque_bytes[65]
port 68 nsew
flabel metal2 s 486 -22 490 -18 7 FreeSans 24 270 0 0 bloque_bytes[66]
port 69 nsew
flabel metal2 s 526 -22 530 -18 7 FreeSans 24 270 0 0 bloque_bytes[67]
port 70 nsew
flabel metal2 s 1174 -22 1178 -18 7 FreeSans 24 270 0 0 bloque_bytes[68]
port 71 nsew
flabel metal2 s 1110 -22 1114 -18 7 FreeSans 24 270 0 0 bloque_bytes[69]
port 72 nsew
flabel metal2 s 2294 -22 2298 -18 7 FreeSans 24 270 0 0 bloque_bytes[70]
port 73 nsew
flabel metal2 s 2150 -22 2154 -18 7 FreeSans 24 270 0 0 bloque_bytes[71]
port 74 nsew
flabel metal2 s 3006 -22 3010 -18 7 FreeSans 24 270 0 0 bloque_bytes[72]
port 75 nsew
flabel metal2 s 2510 -22 2514 -18 7 FreeSans 24 270 0 0 bloque_bytes[73]
port 76 nsew
flabel metal2 s 2942 -22 2946 -18 7 FreeSans 24 270 0 0 bloque_bytes[74]
port 77 nsew
flabel metal2 s 2982 -22 2986 -18 7 FreeSans 24 270 0 0 bloque_bytes[75]
port 78 nsew
flabel metal2 s 3182 -22 3186 -18 7 FreeSans 24 270 0 0 bloque_bytes[76]
port 79 nsew
flabel metal2 s 3878 -22 3882 -18 7 FreeSans 24 270 0 0 bloque_bytes[77]
port 80 nsew
flabel metal2 s 4118 -22 4122 -18 7 FreeSans 24 270 0 0 bloque_bytes[78]
port 81 nsew
flabel metal2 s 4094 -22 4098 -18 7 FreeSans 24 270 0 0 bloque_bytes[79]
port 82 nsew
flabel metal2 s 3990 -22 3994 -18 7 FreeSans 24 270 0 0 bloque_bytes[80]
port 83 nsew
flabel metal2 s 4230 -22 4234 -18 7 FreeSans 24 270 0 0 bloque_bytes[81]
port 84 nsew
flabel metal2 s 4214 -22 4218 -18 7 FreeSans 24 270 0 0 bloque_bytes[82]
port 85 nsew
flabel metal2 s 4046 -22 4050 -18 7 FreeSans 24 270 0 0 bloque_bytes[83]
port 86 nsew
flabel metal2 s 4022 -22 4026 -18 7 FreeSans 24 270 0 0 bloque_bytes[84]
port 87 nsew
flabel metal2 s 3342 -22 3346 -18 7 FreeSans 24 270 0 0 bloque_bytes[85]
port 88 nsew
flabel metal2 s 4534 -22 4538 -18 7 FreeSans 24 270 0 0 bloque_bytes[86]
port 89 nsew
flabel metal2 s 4974 -22 4978 -18 7 FreeSans 24 270 0 0 bloque_bytes[87]
port 90 nsew
flabel metal2 s 4422 -22 4426 -18 7 FreeSans 24 270 0 0 bloque_bytes[88]
port 91 nsew
flabel metal3 s 5342 568 5346 572 3 FreeSans 24 0 0 0 bloque_bytes[89]
port 92 nsew
flabel metal3 s 5342 548 5346 552 3 FreeSans 24 0 0 0 bloque_bytes[90]
port 93 nsew
flabel metal3 s 5342 448 5346 452 3 FreeSans 24 0 0 0 bloque_bytes[91]
port 94 nsew
flabel metal2 s 5230 -22 5234 -18 7 FreeSans 24 270 0 0 bloque_bytes[92]
port 95 nsew
flabel metal2 s 5246 -22 5250 -18 7 FreeSans 24 270 0 0 bloque_bytes[93]
port 96 nsew
flabel metal2 s 5214 -22 5218 -18 7 FreeSans 24 270 0 0 bloque_bytes[94]
port 97 nsew
flabel metal2 s 4686 -22 4690 -18 7 FreeSans 24 270 0 0 bloque_bytes[95]
port 98 nsew
flabel metal2 s 3958 3728 3962 3732 3 FreeSans 24 90 0 0 clk
port 99 nsew
flabel metal2 s 3502 -22 3506 -18 7 FreeSans 24 270 0 0 reset
port 100 nsew
flabel metal3 s 5342 3248 5346 3252 3 FreeSans 24 0 0 0 target[0]
port 101 nsew
flabel metal3 s 5342 3268 5346 3272 3 FreeSans 24 0 0 0 target[1]
port 102 nsew
flabel metal2 s 4886 3728 4890 3732 3 FreeSans 24 90 0 0 target[2]
port 103 nsew
flabel metal2 s 4862 3728 4866 3732 3 FreeSans 24 90 0 0 target[3]
port 104 nsew
flabel metal2 s 4358 3728 4362 3732 3 FreeSans 24 90 0 0 target[4]
port 105 nsew
flabel metal2 s 4342 3728 4346 3732 3 FreeSans 24 90 0 0 target[5]
port 106 nsew
flabel metal2 s 4198 3728 4202 3732 3 FreeSans 24 90 0 0 target[6]
port 107 nsew
flabel metal2 s 4238 3728 4242 3732 3 FreeSans 24 90 0 0 target[7]
port 108 nsew
flabel metal2 s 3654 3728 3658 3732 3 FreeSans 24 90 0 0 terminado
port 109 nsew
flabel metal2 s 2942 3728 2946 3732 3 FreeSans 24 90 0 0 hash[0]
port 110 nsew
flabel metal2 s 3166 3728 3170 3732 3 FreeSans 24 90 0 0 hash[1]
port 111 nsew
flabel metal2 s 3374 3728 3378 3732 3 FreeSans 24 90 0 0 hash[2]
port 112 nsew
flabel metal2 s 2982 3728 2986 3732 3 FreeSans 24 90 0 0 hash[3]
port 113 nsew
flabel metal2 s 3790 3728 3794 3732 3 FreeSans 24 90 0 0 hash[4]
port 114 nsew
flabel metal2 s 3302 3728 3306 3732 3 FreeSans 24 90 0 0 hash[5]
port 115 nsew
flabel metal2 s 3678 3728 3682 3732 3 FreeSans 24 90 0 0 hash[6]
port 116 nsew
flabel metal2 s 2758 3728 2762 3732 3 FreeSans 24 90 0 0 hash[7]
port 117 nsew
flabel metal3 s 5342 2848 5346 2852 3 FreeSans 24 0 0 0 hash[8]
port 118 nsew
flabel metal3 s 5342 2948 5346 2952 3 FreeSans 24 0 0 0 hash[9]
port 119 nsew
flabel metal2 s 5174 3728 5178 3732 3 FreeSans 24 90 0 0 hash[10]
port 120 nsew
flabel metal2 s 5222 3728 5226 3732 3 FreeSans 24 90 0 0 hash[11]
port 121 nsew
flabel metal2 s 4430 3728 4434 3732 3 FreeSans 24 90 0 0 hash[12]
port 122 nsew
flabel metal2 s 4582 3728 4586 3732 3 FreeSans 24 90 0 0 hash[13]
port 123 nsew
flabel metal2 s 4078 3728 4082 3732 3 FreeSans 24 90 0 0 hash[14]
port 124 nsew
flabel metal2 s 5238 3728 5242 3732 3 FreeSans 24 90 0 0 hash[15]
port 125 nsew
flabel metal3 s 5342 3168 5346 3172 3 FreeSans 24 0 0 0 hash[16]
port 126 nsew
flabel metal3 s 5342 3048 5346 3052 3 FreeSans 24 0 0 0 hash[17]
port 127 nsew
flabel metal2 s 4766 3728 4770 3732 3 FreeSans 24 90 0 0 hash[18]
port 128 nsew
flabel metal3 s 5342 3148 5346 3152 3 FreeSans 24 0 0 0 hash[19]
port 129 nsew
flabel metal2 s 3974 3728 3978 3732 3 FreeSans 24 90 0 0 hash[20]
port 130 nsew
flabel metal2 s 3630 3728 3634 3732 3 FreeSans 24 90 0 0 hash[21]
port 131 nsew
flabel metal2 s 4110 3728 4114 3732 3 FreeSans 24 90 0 0 hash[22]
port 132 nsew
flabel metal2 s 3398 3728 3402 3732 3 FreeSans 24 90 0 0 hash[23]
port 133 nsew
<< end >>
