module modulo_rendimiento (inicio, bloque_bytes, clk, reset, target, terminado, hash);

input inicio;
input clk;
input reset;
output terminado;
input [95:0] bloque_bytes;
input [7:0] target;
output [23:0] hash;

wire vdd = 1'b1;
wire gnd = 1'b0;

BUFX4 BUFX4_1 ( .A(_127_), .Y(_127__bF_buf4) );
BUFX4 BUFX4_2 ( .A(_127_), .Y(_127__bF_buf3) );
BUFX4 BUFX4_3 ( .A(_127_), .Y(_127__bF_buf2) );
BUFX4 BUFX4_4 ( .A(_127_), .Y(_127__bF_buf1) );
BUFX4 BUFX4_5 ( .A(_127_), .Y(_127__bF_buf0) );
CLKBUF1 CLKBUF1_1 ( .A(clk), .Y(clk_bF_buf9) );
CLKBUF1 CLKBUF1_2 ( .A(clk), .Y(clk_bF_buf8) );
CLKBUF1 CLKBUF1_3 ( .A(clk), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_4 ( .A(clk), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_5 ( .A(clk), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_6 ( .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_7 ( .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_8 ( .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_9 ( .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_10 ( .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_6 ( .A(_3299_), .Y(_3299__bF_buf4) );
BUFX4 BUFX4_7 ( .A(_3299_), .Y(_3299__bF_buf3) );
BUFX4 BUFX4_8 ( .A(_3299_), .Y(_3299__bF_buf2) );
BUFX4 BUFX4_9 ( .A(_3299_), .Y(_3299__bF_buf1) );
BUFX4 BUFX4_10 ( .A(_3299_), .Y(_3299__bF_buf0) );
BUFX4 BUFX4_11 ( .A(_85_), .Y(_85__bF_buf4) );
BUFX4 BUFX4_12 ( .A(_85_), .Y(_85__bF_buf3) );
BUFX4 BUFX4_13 ( .A(_85_), .Y(_85__bF_buf2) );
BUFX4 BUFX4_14 ( .A(_85_), .Y(_85__bF_buf1) );
BUFX4 BUFX4_15 ( .A(_85_), .Y(_85__bF_buf0) );
BUFX4 BUFX4_16 ( .A(_110_), .Y(_110__bF_buf4) );
BUFX4 BUFX4_17 ( .A(_110_), .Y(_110__bF_buf3) );
BUFX4 BUFX4_18 ( .A(_110_), .Y(_110__bF_buf2) );
BUFX4 BUFX4_19 ( .A(_110_), .Y(_110__bF_buf1) );
BUFX4 BUFX4_20 ( .A(_110_), .Y(_110__bF_buf0) );
BUFX4 BUFX4_21 ( .A(reset), .Y(reset_bF_buf5) );
BUFX4 BUFX4_22 ( .A(reset), .Y(reset_bF_buf4) );
BUFX4 BUFX4_23 ( .A(reset), .Y(reset_bF_buf3) );
BUFX4 BUFX4_24 ( .A(reset), .Y(reset_bF_buf2) );
BUFX4 BUFX4_25 ( .A(reset), .Y(reset_bF_buf1) );
BUFX4 BUFX4_26 ( .A(reset), .Y(reset_bF_buf0) );
INVX8 INVX8_1 ( .A(reset_bF_buf1), .Y(_110_) );
NOR2X1 NOR2X1_1 ( .A(target[7]), .B(micro_ucr_hash1_hash_15_), .Y(_111_) );
NAND2X1 NAND2X1_1 ( .A(target[7]), .B(micro_ucr_hash1_hash_15_), .Y(_112_) );
INVX1 INVX1_1 ( .A(_112_), .Y(_113_) );
XNOR2X1 XNOR2X1_1 ( .A(target[6]), .B(micro_ucr_hash1_hash_14_), .Y(_114_) );
OAI21X1 OAI21X1_1 ( .A(_111_), .B(_113_), .C(_114_), .Y(_115_) );
INVX2 INVX2_1 ( .A(micro_ucr_hash1_hash_13_), .Y(_116_) );
INVX2 INVX2_2 ( .A(micro_ucr_hash1_hash_12_), .Y(_117_) );
AOI22X1 AOI22X1_1 ( .A(_116_), .B(target[5]), .C(target[4]), .D(_117_), .Y(_118_) );
INVX4 INVX4_1 ( .A(target[5]), .Y(_119_) );
INVX2 INVX2_3 ( .A(target[4]), .Y(_120_) );
AOI22X1 AOI22X1_2 ( .A(_119_), .B(micro_ucr_hash1_hash_13_), .C(_120_), .D(micro_ucr_hash1_hash_12_), .Y(_121_) );
NAND2X1 NAND2X1_2 ( .A(_118_), .B(_121_), .Y(_122_) );
NOR2X1 NOR2X1_2 ( .A(_122_), .B(_115_), .Y(_123_) );
XNOR2X1 XNOR2X1_2 ( .A(target[3]), .B(micro_ucr_hash1_hash_11_), .Y(_124_) );
XNOR2X1 XNOR2X1_3 ( .A(target[2]), .B(micro_ucr_hash1_hash_10_), .Y(_125_) );
NAND2X1 NAND2X1_3 ( .A(_124_), .B(_125_), .Y(_2_) );
INVX2 INVX2_4 ( .A(target[1]), .Y(_3_) );
NOR2X1 NOR2X1_3 ( .A(micro_ucr_hash1_hash_9_), .B(_3_), .Y(_4_) );
INVX2 INVX2_5 ( .A(target[0]), .Y(_5_) );
NAND2X1 NAND2X1_4 ( .A(micro_ucr_hash1_hash_8_), .B(_5_), .Y(_6_) );
NAND2X1 NAND2X1_5 ( .A(micro_ucr_hash1_hash_9_), .B(_3_), .Y(_7_) );
AOI21X1 AOI21X1_1 ( .A(_6_), .B(_7_), .C(_4_), .Y(_8_) );
INVX2 INVX2_6 ( .A(target[3]), .Y(_9_) );
NOR2X1 NOR2X1_4 ( .A(micro_ucr_hash1_hash_11_), .B(_9_), .Y(_10_) );
NAND2X1 NAND2X1_6 ( .A(micro_ucr_hash1_hash_11_), .B(_9_), .Y(_11_) );
INVX2 INVX2_7 ( .A(target[2]), .Y(_12_) );
NOR2X1 NOR2X1_5 ( .A(micro_ucr_hash1_hash_10_), .B(_12_), .Y(_13_) );
AOI21X1 AOI21X1_2 ( .A(_11_), .B(_13_), .C(_10_), .Y(_14_) );
OAI21X1 OAI21X1_2 ( .A(_2_), .B(_8_), .C(_14_), .Y(_15_) );
NAND2X1 NAND2X1_7 ( .A(_123_), .B(_15_), .Y(_16_) );
INVX1 INVX1_2 ( .A(_111_), .Y(_17_) );
XOR2X1 XOR2X1_1 ( .A(target[6]), .B(micro_ucr_hash1_hash_14_), .Y(_18_) );
AOI21X1 AOI21X1_3 ( .A(_17_), .B(_112_), .C(_18_), .Y(_19_) );
NAND2X1 NAND2X1_8 ( .A(target[5]), .B(_116_), .Y(_20_) );
NAND2X1 NAND2X1_9 ( .A(target[4]), .B(_117_), .Y(_21_) );
NOR2X1 NOR2X1_6 ( .A(target[5]), .B(_116_), .Y(_22_) );
OAI21X1 OAI21X1_3 ( .A(_22_), .B(_21_), .C(_20_), .Y(_23_) );
INVX2 INVX2_8 ( .A(target[7]), .Y(_24_) );
INVX2 INVX2_9 ( .A(target[6]), .Y(_25_) );
NOR2X1 NOR2X1_7 ( .A(micro_ucr_hash1_hash_14_), .B(_25_), .Y(_26_) );
OAI21X1 OAI21X1_4 ( .A(_113_), .B(_111_), .C(_26_), .Y(_27_) );
OAI21X1 OAI21X1_5 ( .A(_24_), .B(micro_ucr_hash1_hash_15_), .C(_27_), .Y(_28_) );
AOI21X1 AOI21X1_4 ( .A(_23_), .B(_19_), .C(_28_), .Y(_29_) );
OAI22X1 OAI22X1_1 ( .A(_119_), .B(micro_ucr_hash1_hash_13_), .C(_120_), .D(micro_ucr_hash1_hash_12_), .Y(_30_) );
OAI22X1 OAI22X1_2 ( .A(_116_), .B(target[5]), .C(target[4]), .D(_117_), .Y(_31_) );
NOR2X1 NOR2X1_8 ( .A(_30_), .B(_31_), .Y(_32_) );
NAND2X1 NAND2X1_10 ( .A(_32_), .B(_19_), .Y(_33_) );
INVX1 INVX1_3 ( .A(micro_ucr_hash1_hash_9_), .Y(_34_) );
INVX1 INVX1_4 ( .A(micro_ucr_hash1_hash_8_), .Y(_35_) );
OAI22X1 OAI22X1_3 ( .A(_34_), .B(target[1]), .C(target[0]), .D(_35_), .Y(_36_) );
OAI22X1 OAI22X1_4 ( .A(_3_), .B(micro_ucr_hash1_hash_9_), .C(_5_), .D(micro_ucr_hash1_hash_8_), .Y(_37_) );
NOR2X1 NOR2X1_9 ( .A(_36_), .B(_37_), .Y(_38_) );
NAND3X1 NAND3X1_1 ( .A(_124_), .B(_125_), .C(_38_), .Y(_39_) );
NOR2X1 NOR2X1_10 ( .A(_33_), .B(_39_), .Y(_40_) );
AOI21X1 AOI21X1_5 ( .A(_29_), .B(_16_), .C(_40_), .Y(_41_) );
INVX1 INVX1_5 ( .A(micro_ucr_hash1_hash_23_), .Y(_42_) );
INVX1 INVX1_6 ( .A(micro_ucr_hash1_hash_22_), .Y(_43_) );
AOI22X1 AOI22X1_3 ( .A(_42_), .B(target[7]), .C(_43_), .D(target[6]), .Y(_44_) );
NAND2X1 NAND2X1_11 ( .A(micro_ucr_hash1_hash_23_), .B(_24_), .Y(_45_) );
NAND2X1 NAND2X1_12 ( .A(micro_ucr_hash1_hash_22_), .B(_25_), .Y(_46_) );
NAND3X1 NAND3X1_2 ( .A(_45_), .B(_46_), .C(_44_), .Y(_47_) );
INVX1 INVX1_7 ( .A(micro_ucr_hash1_hash_21_), .Y(_48_) );
INVX1 INVX1_8 ( .A(micro_ucr_hash1_hash_20_), .Y(_49_) );
AOI22X1 AOI22X1_4 ( .A(_48_), .B(target[5]), .C(_49_), .D(target[4]), .Y(_50_) );
NAND2X1 NAND2X1_13 ( .A(micro_ucr_hash1_hash_21_), .B(_119_), .Y(_51_) );
NAND2X1 NAND2X1_14 ( .A(micro_ucr_hash1_hash_20_), .B(_120_), .Y(_52_) );
NAND3X1 NAND3X1_3 ( .A(_51_), .B(_52_), .C(_50_), .Y(_53_) );
NOR2X1 NOR2X1_11 ( .A(_47_), .B(_53_), .Y(_54_) );
INVX2 INVX2_10 ( .A(micro_ucr_hash1_hash_19_), .Y(_55_) );
INVX1 INVX1_9 ( .A(micro_ucr_hash1_hash_18_), .Y(_56_) );
AOI22X1 AOI22X1_5 ( .A(_55_), .B(target[3]), .C(_56_), .D(target[2]), .Y(_57_) );
AOI22X1 AOI22X1_6 ( .A(_9_), .B(micro_ucr_hash1_hash_19_), .C(micro_ucr_hash1_hash_18_), .D(_12_), .Y(_58_) );
NAND2X1 NAND2X1_15 ( .A(_57_), .B(_58_), .Y(_59_) );
NOR2X1 NOR2X1_12 ( .A(micro_ucr_hash1_hash_17_), .B(_3_), .Y(_60_) );
NAND2X1 NAND2X1_16 ( .A(micro_ucr_hash1_hash_16_), .B(_5_), .Y(_61_) );
NAND2X1 NAND2X1_17 ( .A(micro_ucr_hash1_hash_17_), .B(_3_), .Y(_62_) );
AOI21X1 AOI21X1_6 ( .A(_61_), .B(_62_), .C(_60_), .Y(_63_) );
OAI22X1 OAI22X1_5 ( .A(_9_), .B(micro_ucr_hash1_hash_19_), .C(micro_ucr_hash1_hash_18_), .D(_12_), .Y(_64_) );
OAI21X1 OAI21X1_6 ( .A(_55_), .B(target[3]), .C(_64_), .Y(_65_) );
OAI21X1 OAI21X1_7 ( .A(_59_), .B(_63_), .C(_65_), .Y(_66_) );
NAND2X1 NAND2X1_18 ( .A(_66_), .B(_54_), .Y(_67_) );
OAI22X1 OAI22X1_6 ( .A(_24_), .B(micro_ucr_hash1_hash_23_), .C(micro_ucr_hash1_hash_22_), .D(_25_), .Y(_68_) );
OAI22X1 OAI22X1_7 ( .A(_42_), .B(target[7]), .C(_43_), .D(target[6]), .Y(_69_) );
NOR2X1 NOR2X1_13 ( .A(_68_), .B(_69_), .Y(_70_) );
AOI21X1 AOI21X1_7 ( .A(micro_ucr_hash1_hash_21_), .B(_119_), .C(_50_), .Y(_71_) );
AOI22X1 AOI22X1_7 ( .A(_68_), .B(_45_), .C(_70_), .D(_71_), .Y(_72_) );
OAI22X1 OAI22X1_8 ( .A(_119_), .B(micro_ucr_hash1_hash_21_), .C(micro_ucr_hash1_hash_20_), .D(_120_), .Y(_73_) );
OAI22X1 OAI22X1_9 ( .A(_48_), .B(target[5]), .C(_49_), .D(target[4]), .Y(_74_) );
NOR2X1 NOR2X1_14 ( .A(_73_), .B(_74_), .Y(_75_) );
NAND2X1 NAND2X1_19 ( .A(_70_), .B(_75_), .Y(_76_) );
OAI22X1 OAI22X1_10 ( .A(_55_), .B(target[3]), .C(_56_), .D(target[2]), .Y(_77_) );
NOR2X1 NOR2X1_15 ( .A(_64_), .B(_77_), .Y(_78_) );
AND2X2 AND2X2_1 ( .A(_61_), .B(_62_), .Y(_79_) );
INVX1 INVX1_10 ( .A(micro_ucr_hash1_hash_16_), .Y(_80_) );
AOI21X1 AOI21X1_8 ( .A(_80_), .B(target[0]), .C(_60_), .Y(_81_) );
NAND3X1 NAND3X1_4 ( .A(_79_), .B(_81_), .C(_78_), .Y(_82_) );
NOR2X1 NOR2X1_16 ( .A(_76_), .B(_82_), .Y(_83_) );
AOI21X1 AOI21X1_9 ( .A(_67_), .B(_72_), .C(_83_), .Y(_84_) );
AOI21X1 AOI21X1_10 ( .A(_84_), .B(_41_), .C(_127__bF_buf4), .Y(_85_) );
NOR2X1 NOR2X1_17 ( .A(_110__bF_buf1), .B(_85__bF_buf2), .Y(_1_) );
MUX2X1 MUX2X1_1 ( .A(_126__0_), .B(micro_ucr_hash1_hash_0_), .S(_127__bF_buf3), .Y(_86_) );
NOR3X1 NOR3X1_1 ( .A(_110__bF_buf4), .B(_86_), .C(_85__bF_buf3), .Y(_0__0_) );
MUX2X1 MUX2X1_2 ( .A(_126__1_), .B(micro_ucr_hash1_hash_1_), .S(_127__bF_buf3), .Y(_87_) );
NOR3X1 NOR3X1_2 ( .A(_110__bF_buf4), .B(_87_), .C(_85__bF_buf3), .Y(_0__1_) );
MUX2X1 MUX2X1_3 ( .A(_126__2_), .B(micro_ucr_hash1_hash_2_), .S(_127__bF_buf3), .Y(_88_) );
NOR3X1 NOR3X1_3 ( .A(_110__bF_buf4), .B(_88_), .C(_85__bF_buf3), .Y(_0__2_) );
MUX2X1 MUX2X1_4 ( .A(_126__3_), .B(micro_ucr_hash1_hash_3_), .S(_127__bF_buf3), .Y(_89_) );
NOR3X1 NOR3X1_4 ( .A(_110__bF_buf3), .B(_89_), .C(_85__bF_buf0), .Y(_0__3_) );
MUX2X1 MUX2X1_5 ( .A(_126__4_), .B(micro_ucr_hash1_hash_4_), .S(_127__bF_buf3), .Y(_90_) );
NOR3X1 NOR3X1_5 ( .A(_110__bF_buf4), .B(_90_), .C(_85__bF_buf3), .Y(_0__4_) );
MUX2X1 MUX2X1_6 ( .A(_126__5_), .B(micro_ucr_hash1_hash_5_), .S(_127__bF_buf2), .Y(_91_) );
NOR3X1 NOR3X1_6 ( .A(_110__bF_buf3), .B(_91_), .C(_85__bF_buf0), .Y(_0__5_) );
MUX2X1 MUX2X1_7 ( .A(_126__6_), .B(micro_ucr_hash1_hash_6_), .S(_127__bF_buf3), .Y(_92_) );
NOR3X1 NOR3X1_7 ( .A(_110__bF_buf4), .B(_92_), .C(_85__bF_buf3), .Y(_0__6_) );
MUX2X1 MUX2X1_8 ( .A(_126__7_), .B(micro_ucr_hash1_hash_7_), .S(_127__bF_buf2), .Y(_93_) );
NOR3X1 NOR3X1_8 ( .A(_110__bF_buf3), .B(_93_), .C(_85__bF_buf0), .Y(_0__7_) );
MUX2X1 MUX2X1_9 ( .A(_126__8_), .B(micro_ucr_hash1_hash_8_), .S(_127__bF_buf1), .Y(_94_) );
NOR3X1 NOR3X1_9 ( .A(_110__bF_buf0), .B(_94_), .C(_85__bF_buf4), .Y(_0__8_) );
MUX2X1 MUX2X1_10 ( .A(_126__9_), .B(micro_ucr_hash1_hash_9_), .S(_127__bF_buf1), .Y(_95_) );
NOR3X1 NOR3X1_10 ( .A(_110__bF_buf0), .B(_95_), .C(_85__bF_buf4), .Y(_0__9_) );
MUX2X1 MUX2X1_11 ( .A(_126__10_), .B(micro_ucr_hash1_hash_10_), .S(_127__bF_buf1), .Y(_96_) );
NOR3X1 NOR3X1_11 ( .A(_110__bF_buf0), .B(_96_), .C(_85__bF_buf4), .Y(_0__10_) );
MUX2X1 MUX2X1_12 ( .A(_126__11_), .B(micro_ucr_hash1_hash_11_), .S(_127__bF_buf4), .Y(_97_) );
NOR3X1 NOR3X1_12 ( .A(_110__bF_buf1), .B(_97_), .C(_85__bF_buf2), .Y(_0__11_) );
MUX2X1 MUX2X1_13 ( .A(_126__12_), .B(micro_ucr_hash1_hash_12_), .S(_127__bF_buf0), .Y(_98_) );
NOR3X1 NOR3X1_13 ( .A(_110__bF_buf1), .B(_98_), .C(_85__bF_buf2), .Y(_0__12_) );
MUX2X1 MUX2X1_14 ( .A(_126__13_), .B(micro_ucr_hash1_hash_13_), .S(_127__bF_buf0), .Y(_99_) );
NOR3X1 NOR3X1_14 ( .A(_110__bF_buf1), .B(_99_), .C(_85__bF_buf2), .Y(_0__13_) );
MUX2X1 MUX2X1_15 ( .A(_126__14_), .B(micro_ucr_hash1_hash_14_), .S(_127__bF_buf4), .Y(_100_) );
NOR3X1 NOR3X1_15 ( .A(_110__bF_buf1), .B(_100_), .C(_85__bF_buf2), .Y(_0__14_) );
MUX2X1 MUX2X1_16 ( .A(_126__15_), .B(micro_ucr_hash1_hash_15_), .S(_127__bF_buf1), .Y(_101_) );
NOR3X1 NOR3X1_16 ( .A(_110__bF_buf0), .B(_101_), .C(_85__bF_buf4), .Y(_0__15_) );
MUX2X1 MUX2X1_17 ( .A(_126__16_), .B(micro_ucr_hash1_hash_16_), .S(_127__bF_buf1), .Y(_102_) );
NOR3X1 NOR3X1_17 ( .A(_110__bF_buf0), .B(_102_), .C(_85__bF_buf4), .Y(_0__16_) );
MUX2X1 MUX2X1_18 ( .A(_126__17_), .B(micro_ucr_hash1_hash_17_), .S(_127__bF_buf4), .Y(_103_) );
NOR3X1 NOR3X1_18 ( .A(_110__bF_buf2), .B(_103_), .C(_85__bF_buf1), .Y(_0__17_) );
MUX2X1 MUX2X1_19 ( .A(_126__18_), .B(micro_ucr_hash1_hash_18_), .S(_127__bF_buf4), .Y(_104_) );
NOR3X1 NOR3X1_19 ( .A(_110__bF_buf2), .B(_104_), .C(_85__bF_buf1), .Y(_0__18_) );
MUX2X1 MUX2X1_20 ( .A(_126__19_), .B(micro_ucr_hash1_hash_19_), .S(_127__bF_buf2), .Y(_105_) );
NOR3X1 NOR3X1_20 ( .A(_110__bF_buf2), .B(_105_), .C(_85__bF_buf1), .Y(_0__19_) );
MUX2X1 MUX2X1_21 ( .A(_126__20_), .B(micro_ucr_hash1_hash_20_), .S(_127__bF_buf2), .Y(_106_) );
NOR3X1 NOR3X1_21 ( .A(_110__bF_buf2), .B(_106_), .C(_85__bF_buf1), .Y(_0__20_) );
MUX2X1 MUX2X1_22 ( .A(_126__21_), .B(micro_ucr_hash1_hash_21_), .S(_127__bF_buf4), .Y(_107_) );
NOR3X1 NOR3X1_22 ( .A(_110__bF_buf2), .B(_107_), .C(_85__bF_buf1), .Y(_0__21_) );
MUX2X1 MUX2X1_23 ( .A(_126__22_), .B(micro_ucr_hash1_hash_22_), .S(_127__bF_buf2), .Y(_108_) );
NOR3X1 NOR3X1_23 ( .A(_110__bF_buf3), .B(_108_), .C(_85__bF_buf0), .Y(_0__22_) );
MUX2X1 MUX2X1_24 ( .A(_126__23_), .B(micro_ucr_hash1_hash_23_), .S(_127__bF_buf2), .Y(_109_) );
NOR3X1 NOR3X1_24 ( .A(_110__bF_buf3), .B(_109_), .C(_85__bF_buf0), .Y(_0__23_) );
BUFX2 BUFX2_1 ( .A(_126__0_), .Y(hash[0]) );
BUFX2 BUFX2_2 ( .A(_126__1_), .Y(hash[1]) );
BUFX2 BUFX2_3 ( .A(_126__2_), .Y(hash[2]) );
BUFX2 BUFX2_4 ( .A(_126__3_), .Y(hash[3]) );
BUFX2 BUFX2_5 ( .A(_126__4_), .Y(hash[4]) );
BUFX2 BUFX2_6 ( .A(_126__5_), .Y(hash[5]) );
BUFX2 BUFX2_7 ( .A(_126__6_), .Y(hash[6]) );
BUFX2 BUFX2_8 ( .A(_126__7_), .Y(hash[7]) );
BUFX2 BUFX2_9 ( .A(_126__8_), .Y(hash[8]) );
BUFX2 BUFX2_10 ( .A(_126__9_), .Y(hash[9]) );
BUFX2 BUFX2_11 ( .A(_126__10_), .Y(hash[10]) );
BUFX2 BUFX2_12 ( .A(_126__11_), .Y(hash[11]) );
BUFX2 BUFX2_13 ( .A(_126__12_), .Y(hash[12]) );
BUFX2 BUFX2_14 ( .A(_126__13_), .Y(hash[13]) );
BUFX2 BUFX2_15 ( .A(_126__14_), .Y(hash[14]) );
BUFX2 BUFX2_16 ( .A(_126__15_), .Y(hash[15]) );
BUFX2 BUFX2_17 ( .A(_126__16_), .Y(hash[16]) );
BUFX2 BUFX2_18 ( .A(_126__17_), .Y(hash[17]) );
BUFX2 BUFX2_19 ( .A(_126__18_), .Y(hash[18]) );
BUFX2 BUFX2_20 ( .A(_126__19_), .Y(hash[19]) );
BUFX2 BUFX2_21 ( .A(_126__20_), .Y(hash[20]) );
BUFX2 BUFX2_22 ( .A(_126__21_), .Y(hash[21]) );
BUFX2 BUFX2_23 ( .A(_126__22_), .Y(hash[22]) );
BUFX2 BUFX2_24 ( .A(_126__23_), .Y(hash[23]) );
BUFX2 BUFX2_25 ( .A(_127__bF_buf1), .Y(terminado) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf0), .D(_1_), .Q(_127_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf6), .D(_0__0_), .Q(_126__0_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf8), .D(_0__1_), .Q(_126__1_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf8), .D(_0__2_), .Q(_126__2_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf8), .D(_0__3_), .Q(_126__3_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf6), .D(_0__4_), .Q(_126__4_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf6), .D(_0__5_), .Q(_126__5_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf6), .D(_0__6_), .Q(_126__6_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf8), .D(_0__7_), .Q(_126__7_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf2), .D(_0__8_), .Q(_126__8_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf2), .D(_0__9_), .Q(_126__9_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf2), .D(_0__10_), .Q(_126__10_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf2), .D(_0__11_), .Q(_126__11_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf4), .D(_0__12_), .Q(_126__12_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf0), .D(_0__13_), .Q(_126__13_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf2), .D(_0__14_), .Q(_126__14_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf2), .D(_0__15_), .Q(_126__15_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf2), .D(_0__16_), .Q(_126__16_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf0), .D(_0__17_), .Q(_126__17_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf0), .D(_0__18_), .Q(_126__18_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf0), .D(_0__19_), .Q(_126__19_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf0), .D(_0__20_), .Q(_126__20_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf0), .D(_0__21_), .Q(_126__21_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf0), .D(_0__22_), .Q(_126__22_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf6), .D(_0__23_), .Q(_126__23_) );
XOR2X1 XOR2X1_2 ( .A(micro_ucr_hash1_b_1__4_), .B(gnd), .Y(micro_ucr_hash1_a_1__0_) );
XOR2X1 XOR2X1_3 ( .A(micro_ucr_hash1_b_1__5_), .B(gnd), .Y(micro_ucr_hash1_a_1__1_) );
XOR2X1 XOR2X1_4 ( .A(micro_ucr_hash1_b_1__6_), .B(gnd), .Y(micro_ucr_hash1_a_1__2_) );
XOR2X1 XOR2X1_5 ( .A(micro_ucr_hash1_b_1__7_), .B(gnd), .Y(micro_ucr_hash1_a_1__3_) );
XOR2X1 XOR2X1_6 ( .A(micro_ucr_hash1_c_0__4_), .B(gnd), .Y(micro_ucr_hash1_a_1__4_) );
XOR2X1 XOR2X1_7 ( .A(micro_ucr_hash1_c_0__5_), .B(vdd), .Y(micro_ucr_hash1_a_1__5_) );
XOR2X1 XOR2X1_8 ( .A(micro_ucr_hash1_c_0__6_), .B(vdd), .Y(micro_ucr_hash1_a_1__6_) );
XOR2X1 XOR2X1_9 ( .A(micro_ucr_hash1_c_0__7_), .B(vdd), .Y(micro_ucr_hash1_a_1__7_) );
INVX2 INVX2_11 ( .A(bloque_bytes[80]), .Y(_197_) );
XNOR2X1 XNOR2X1_4 ( .A(gnd), .B(micro_ucr_hash1_a_0__0_), .Y(_198_) );
XNOR2X1 XNOR2X1_5 ( .A(_198_), .B(_197_), .Y(micro_ucr_hash1_b_2__4_) );
NAND2X1 NAND2X1_20 ( .A(_197_), .B(_198_), .Y(_199_) );
OR2X2 OR2X2_1 ( .A(gnd), .B(micro_ucr_hash1_a_0__1_), .Y(_200_) );
NAND2X1 NAND2X1_21 ( .A(gnd), .B(micro_ucr_hash1_a_0__1_), .Y(_201_) );
NAND3X1 NAND3X1_5 ( .A(bloque_bytes[81]), .B(_201_), .C(_200_), .Y(_202_) );
INVX1 INVX1_11 ( .A(bloque_bytes[81]), .Y(_203_) );
NOR2X1 NOR2X1_18 ( .A(gnd), .B(micro_ucr_hash1_a_0__1_), .Y(_204_) );
AND2X2 AND2X2_2 ( .A(gnd), .B(micro_ucr_hash1_a_0__1_), .Y(_205_) );
OAI21X1 OAI21X1_8 ( .A(_205_), .B(_204_), .C(_203_), .Y(_206_) );
NAND2X1 NAND2X1_22 ( .A(_206_), .B(_202_), .Y(_207_) );
XNOR2X1 XNOR2X1_6 ( .A(_207_), .B(_199_), .Y(micro_ucr_hash1_b_2__5_) );
NAND3X1 NAND3X1_6 ( .A(_202_), .B(_206_), .C(_199_), .Y(_208_) );
NOR3X1 NOR3X1_25 ( .A(_203_), .B(_204_), .C(_205_), .Y(_209_) );
INVX1 INVX1_12 ( .A(bloque_bytes[82]), .Y(_210_) );
NOR2X1 NOR2X1_19 ( .A(gnd), .B(micro_ucr_hash1_a_0__2_), .Y(_211_) );
AND2X2 AND2X2_3 ( .A(gnd), .B(micro_ucr_hash1_a_0__2_), .Y(_212_) );
NOR3X1 NOR3X1_26 ( .A(_210_), .B(_211_), .C(_212_), .Y(_213_) );
OR2X2 OR2X2_2 ( .A(gnd), .B(micro_ucr_hash1_a_0__2_), .Y(_214_) );
NAND2X1 NAND2X1_23 ( .A(gnd), .B(micro_ucr_hash1_a_0__2_), .Y(_215_) );
AOI21X1 AOI21X1_11 ( .A(_215_), .B(_214_), .C(bloque_bytes[82]), .Y(_216_) );
OAI21X1 OAI21X1_9 ( .A(_213_), .B(_216_), .C(_209_), .Y(_217_) );
NAND3X1 NAND3X1_7 ( .A(bloque_bytes[82]), .B(_215_), .C(_214_), .Y(_218_) );
OAI21X1 OAI21X1_10 ( .A(_212_), .B(_211_), .C(_210_), .Y(_219_) );
NAND3X1 NAND3X1_8 ( .A(_219_), .B(_202_), .C(_218_), .Y(_220_) );
NAND2X1 NAND2X1_24 ( .A(_220_), .B(_217_), .Y(_221_) );
XNOR2X1 XNOR2X1_7 ( .A(_221_), .B(_208_), .Y(micro_ucr_hash1_b_2__6_) );
NAND3X1 NAND3X1_9 ( .A(_218_), .B(_219_), .C(_209_), .Y(_222_) );
OAI21X1 OAI21X1_11 ( .A(_213_), .B(_216_), .C(_202_), .Y(_223_) );
NAND2X1 NAND2X1_25 ( .A(_222_), .B(_223_), .Y(_224_) );
OAI21X1 OAI21X1_12 ( .A(_224_), .B(_208_), .C(_222_), .Y(_225_) );
INVX1 INVX1_13 ( .A(bloque_bytes[83]), .Y(_226_) );
NOR2X1 NOR2X1_20 ( .A(gnd), .B(micro_ucr_hash1_a_0__3_), .Y(_227_) );
AND2X2 AND2X2_4 ( .A(gnd), .B(micro_ucr_hash1_a_0__3_), .Y(_228_) );
OAI21X1 OAI21X1_13 ( .A(_228_), .B(_227_), .C(_226_), .Y(_229_) );
OR2X2 OR2X2_3 ( .A(gnd), .B(micro_ucr_hash1_a_0__3_), .Y(_230_) );
NAND2X1 NAND2X1_26 ( .A(gnd), .B(micro_ucr_hash1_a_0__3_), .Y(_231_) );
NAND3X1 NAND3X1_10 ( .A(bloque_bytes[83]), .B(_231_), .C(_230_), .Y(_232_) );
AOI21X1 AOI21X1_12 ( .A(_229_), .B(_232_), .C(_218_), .Y(_233_) );
NAND3X1 NAND3X1_11 ( .A(_226_), .B(_231_), .C(_230_), .Y(_234_) );
OAI21X1 OAI21X1_14 ( .A(_228_), .B(_227_), .C(bloque_bytes[83]), .Y(_235_) );
AOI21X1 AOI21X1_13 ( .A(_235_), .B(_234_), .C(_213_), .Y(_236_) );
NOR2X1 NOR2X1_21 ( .A(_233_), .B(_236_), .Y(_128_) );
XOR2X1 XOR2X1_10 ( .A(_225_), .B(_128_), .Y(micro_ucr_hash1_b_2__7_) );
INVX1 INVX1_14 ( .A(bloque_bytes[84]), .Y(_129_) );
OR2X2 OR2X2_4 ( .A(gnd), .B(micro_ucr_hash1_a_0__4_), .Y(_130_) );
NAND2X1 NAND2X1_27 ( .A(gnd), .B(micro_ucr_hash1_a_0__4_), .Y(_131_) );
NAND3X1 NAND3X1_12 ( .A(_129_), .B(_131_), .C(_130_), .Y(_132_) );
NOR2X1 NOR2X1_22 ( .A(gnd), .B(micro_ucr_hash1_a_0__4_), .Y(_133_) );
AND2X2 AND2X2_5 ( .A(gnd), .B(micro_ucr_hash1_a_0__4_), .Y(_134_) );
OAI21X1 OAI21X1_15 ( .A(_134_), .B(_133_), .C(bloque_bytes[84]), .Y(_135_) );
NAND3X1 NAND3X1_13 ( .A(_229_), .B(_132_), .C(_135_), .Y(_136_) );
AOI21X1 AOI21X1_14 ( .A(_231_), .B(_230_), .C(bloque_bytes[83]), .Y(_137_) );
OAI21X1 OAI21X1_16 ( .A(_134_), .B(_133_), .C(_129_), .Y(_138_) );
NAND3X1 NAND3X1_14 ( .A(bloque_bytes[84]), .B(_131_), .C(_130_), .Y(_139_) );
NAND3X1 NAND3X1_15 ( .A(_138_), .B(_139_), .C(_137_), .Y(_140_) );
AND2X2 AND2X2_6 ( .A(_140_), .B(_136_), .Y(_141_) );
INVX2 INVX2_12 ( .A(_236_), .Y(_142_) );
NOR2X1 NOR2X1_23 ( .A(_216_), .B(_213_), .Y(_143_) );
AOI21X1 AOI21X1_15 ( .A(_209_), .B(_143_), .C(_233_), .Y(_144_) );
OAI21X1 OAI21X1_17 ( .A(_224_), .B(_208_), .C(_144_), .Y(_145_) );
NAND2X1 NAND2X1_28 ( .A(_142_), .B(_145_), .Y(_146_) );
XNOR2X1 XNOR2X1_8 ( .A(_146_), .B(_141_), .Y(micro_ucr_hash1_c_1__4_) );
NAND2X1 NAND2X1_29 ( .A(_136_), .B(_140_), .Y(_147_) );
OAI21X1 OAI21X1_18 ( .A(_146_), .B(_147_), .C(_136_), .Y(_148_) );
INVX1 INVX1_15 ( .A(bloque_bytes[85]), .Y(_149_) );
OR2X2 OR2X2_5 ( .A(vdd), .B(micro_ucr_hash1_a_0__5_), .Y(_150_) );
NAND2X1 NAND2X1_30 ( .A(vdd), .B(micro_ucr_hash1_a_0__5_), .Y(_151_) );
NAND3X1 NAND3X1_16 ( .A(_149_), .B(_151_), .C(_150_), .Y(_152_) );
NOR2X1 NOR2X1_24 ( .A(vdd), .B(micro_ucr_hash1_a_0__5_), .Y(_153_) );
AND2X2 AND2X2_7 ( .A(vdd), .B(micro_ucr_hash1_a_0__5_), .Y(_154_) );
OAI21X1 OAI21X1_19 ( .A(_154_), .B(_153_), .C(bloque_bytes[85]), .Y(_155_) );
NAND3X1 NAND3X1_17 ( .A(_138_), .B(_155_), .C(_152_), .Y(_156_) );
AOI21X1 AOI21X1_16 ( .A(_131_), .B(_130_), .C(bloque_bytes[84]), .Y(_157_) );
NAND3X1 NAND3X1_18 ( .A(bloque_bytes[85]), .B(_151_), .C(_150_), .Y(_158_) );
OAI21X1 OAI21X1_20 ( .A(_154_), .B(_153_), .C(_149_), .Y(_159_) );
NAND3X1 NAND3X1_19 ( .A(_159_), .B(_158_), .C(_157_), .Y(_160_) );
NAND2X1 NAND2X1_31 ( .A(_156_), .B(_160_), .Y(_161_) );
INVX2 INVX2_13 ( .A(_161_), .Y(_162_) );
XNOR2X1 XNOR2X1_9 ( .A(_148_), .B(_162_), .Y(micro_ucr_hash1_c_1__5_) );
AOI21X1 AOI21X1_17 ( .A(_156_), .B(_160_), .C(_147_), .Y(_163_) );
NAND3X1 NAND3X1_20 ( .A(_142_), .B(_163_), .C(_145_), .Y(_164_) );
NAND2X1 NAND2X1_32 ( .A(_159_), .B(_158_), .Y(_165_) );
OR2X2 OR2X2_6 ( .A(_165_), .B(_157_), .Y(_166_) );
INVX1 INVX1_16 ( .A(_166_), .Y(_167_) );
AOI21X1 AOI21X1_18 ( .A(_157_), .B(_165_), .C(_136_), .Y(_168_) );
NOR2X1 NOR2X1_25 ( .A(_168_), .B(_167_), .Y(_169_) );
INVX1 INVX1_17 ( .A(bloque_bytes[86]), .Y(_170_) );
XNOR2X1 XNOR2X1_10 ( .A(vdd), .B(micro_ucr_hash1_a_0__6_), .Y(_171_) );
OR2X2 OR2X2_7 ( .A(_171_), .B(_170_), .Y(_172_) );
NAND2X1 NAND2X1_33 ( .A(_170_), .B(_171_), .Y(_173_) );
NAND2X1 NAND2X1_34 ( .A(_173_), .B(_172_), .Y(_174_) );
OR2X2 OR2X2_8 ( .A(_174_), .B(_158_), .Y(_175_) );
NAND2X1 NAND2X1_35 ( .A(_158_), .B(_174_), .Y(_176_) );
NAND2X1 NAND2X1_36 ( .A(_176_), .B(_175_), .Y(_177_) );
AOI21X1 AOI21X1_19 ( .A(_169_), .B(_164_), .C(_177_), .Y(_178_) );
NAND2X1 NAND2X1_37 ( .A(_161_), .B(_141_), .Y(_179_) );
OAI21X1 OAI21X1_21 ( .A(_146_), .B(_179_), .C(_169_), .Y(_180_) );
INVX1 INVX1_18 ( .A(_177_), .Y(_181_) );
NOR2X1 NOR2X1_26 ( .A(_181_), .B(_180_), .Y(_182_) );
NOR2X1 NOR2X1_27 ( .A(_178_), .B(_182_), .Y(micro_ucr_hash1_c_1__6_) );
INVX1 INVX1_19 ( .A(_222_), .Y(_183_) );
AOI21X1 AOI21X1_20 ( .A(_142_), .B(_183_), .C(_233_), .Y(_184_) );
AOI21X1 AOI21X1_21 ( .A(_197_), .B(_198_), .C(_207_), .Y(_185_) );
NAND3X1 NAND3X1_21 ( .A(_185_), .B(_221_), .C(_128_), .Y(_186_) );
AOI21X1 AOI21X1_22 ( .A(_184_), .B(_186_), .C(_179_), .Y(_187_) );
OAI21X1 OAI21X1_22 ( .A(_162_), .B(_136_), .C(_166_), .Y(_188_) );
OAI21X1 OAI21X1_23 ( .A(_187_), .B(_188_), .C(_181_), .Y(_189_) );
XOR2X1 XOR2X1_11 ( .A(vdd), .B(bloque_bytes[87]), .Y(_190_) );
XNOR2X1 XNOR2X1_11 ( .A(_190_), .B(micro_ucr_hash1_a_0__7_), .Y(_191_) );
XNOR2X1 XNOR2X1_12 ( .A(_191_), .B(_172_), .Y(_192_) );
NAND3X1 NAND3X1_22 ( .A(_175_), .B(_192_), .C(_189_), .Y(_193_) );
INVX1 INVX1_20 ( .A(_175_), .Y(_194_) );
INVX1 INVX1_21 ( .A(_192_), .Y(_195_) );
OAI21X1 OAI21X1_24 ( .A(_178_), .B(_194_), .C(_195_), .Y(_196_) );
NAND2X1 NAND2X1_38 ( .A(_193_), .B(_196_), .Y(micro_ucr_hash1_c_1__7_) );
XOR2X1 XOR2X1_12 ( .A(micro_ucr_hash1_b_2__4_), .B(gnd), .Y(micro_ucr_hash1_a_2__0_) );
XOR2X1 XOR2X1_13 ( .A(micro_ucr_hash1_b_2__5_), .B(gnd), .Y(micro_ucr_hash1_a_2__1_) );
XOR2X1 XOR2X1_14 ( .A(micro_ucr_hash1_b_2__6_), .B(gnd), .Y(micro_ucr_hash1_a_2__2_) );
XOR2X1 XOR2X1_15 ( .A(micro_ucr_hash1_b_2__7_), .B(gnd), .Y(micro_ucr_hash1_a_2__3_) );
XOR2X1 XOR2X1_16 ( .A(micro_ucr_hash1_c_1__4_), .B(micro_ucr_hash1_b_1__4_), .Y(micro_ucr_hash1_a_2__4_) );
XOR2X1 XOR2X1_17 ( .A(micro_ucr_hash1_c_1__5_), .B(micro_ucr_hash1_b_1__5_), .Y(micro_ucr_hash1_a_2__5_) );
XOR2X1 XOR2X1_18 ( .A(micro_ucr_hash1_c_1__6_), .B(micro_ucr_hash1_b_1__6_), .Y(micro_ucr_hash1_a_2__6_) );
XOR2X1 XOR2X1_19 ( .A(micro_ucr_hash1_c_1__7_), .B(micro_ucr_hash1_b_1__7_), .Y(micro_ucr_hash1_a_2__7_) );
INVX2 INVX2_14 ( .A(bloque_bytes[72]), .Y(_306_) );
XNOR2X1 XNOR2X1_13 ( .A(gnd), .B(micro_ucr_hash1_a_1__0_), .Y(_307_) );
XNOR2X1 XNOR2X1_14 ( .A(_307_), .B(_306_), .Y(micro_ucr_hash1_b_3__4_) );
NAND2X1 NAND2X1_39 ( .A(_306_), .B(_307_), .Y(_308_) );
OR2X2 OR2X2_9 ( .A(gnd), .B(micro_ucr_hash1_a_1__1_), .Y(_309_) );
NAND2X1 NAND2X1_40 ( .A(gnd), .B(micro_ucr_hash1_a_1__1_), .Y(_310_) );
NAND3X1 NAND3X1_23 ( .A(bloque_bytes[73]), .B(_310_), .C(_309_), .Y(_311_) );
INVX1 INVX1_22 ( .A(bloque_bytes[73]), .Y(_312_) );
NOR2X1 NOR2X1_28 ( .A(gnd), .B(micro_ucr_hash1_a_1__1_), .Y(_313_) );
AND2X2 AND2X2_8 ( .A(gnd), .B(micro_ucr_hash1_a_1__1_), .Y(_314_) );
OAI21X1 OAI21X1_25 ( .A(_314_), .B(_313_), .C(_312_), .Y(_315_) );
NAND2X1 NAND2X1_41 ( .A(_315_), .B(_311_), .Y(_316_) );
XNOR2X1 XNOR2X1_15 ( .A(_316_), .B(_308_), .Y(micro_ucr_hash1_b_3__5_) );
NAND3X1 NAND3X1_24 ( .A(_311_), .B(_315_), .C(_308_), .Y(_317_) );
NOR3X1 NOR3X1_27 ( .A(_312_), .B(_313_), .C(_314_), .Y(_318_) );
INVX1 INVX1_23 ( .A(bloque_bytes[74]), .Y(_319_) );
NOR2X1 NOR2X1_29 ( .A(gnd), .B(micro_ucr_hash1_a_1__2_), .Y(_320_) );
AND2X2 AND2X2_9 ( .A(gnd), .B(micro_ucr_hash1_a_1__2_), .Y(_321_) );
NOR3X1 NOR3X1_28 ( .A(_319_), .B(_320_), .C(_321_), .Y(_322_) );
OR2X2 OR2X2_10 ( .A(gnd), .B(micro_ucr_hash1_a_1__2_), .Y(_323_) );
NAND2X1 NAND2X1_42 ( .A(gnd), .B(micro_ucr_hash1_a_1__2_), .Y(_324_) );
AOI21X1 AOI21X1_23 ( .A(_324_), .B(_323_), .C(bloque_bytes[74]), .Y(_325_) );
OAI21X1 OAI21X1_26 ( .A(_322_), .B(_325_), .C(_318_), .Y(_326_) );
NAND3X1 NAND3X1_25 ( .A(bloque_bytes[74]), .B(_324_), .C(_323_), .Y(_327_) );
OAI21X1 OAI21X1_27 ( .A(_321_), .B(_320_), .C(_319_), .Y(_328_) );
NAND3X1 NAND3X1_26 ( .A(_328_), .B(_311_), .C(_327_), .Y(_329_) );
NAND2X1 NAND2X1_43 ( .A(_329_), .B(_326_), .Y(_330_) );
XNOR2X1 XNOR2X1_16 ( .A(_330_), .B(_317_), .Y(micro_ucr_hash1_b_3__6_) );
NAND3X1 NAND3X1_27 ( .A(_327_), .B(_328_), .C(_318_), .Y(_331_) );
OAI21X1 OAI21X1_28 ( .A(_322_), .B(_325_), .C(_311_), .Y(_332_) );
NAND2X1 NAND2X1_44 ( .A(_331_), .B(_332_), .Y(_333_) );
OAI21X1 OAI21X1_29 ( .A(_333_), .B(_317_), .C(_331_), .Y(_334_) );
INVX1 INVX1_24 ( .A(bloque_bytes[75]), .Y(_335_) );
NOR2X1 NOR2X1_30 ( .A(gnd), .B(micro_ucr_hash1_a_1__3_), .Y(_336_) );
AND2X2 AND2X2_10 ( .A(gnd), .B(micro_ucr_hash1_a_1__3_), .Y(_337_) );
OAI21X1 OAI21X1_30 ( .A(_337_), .B(_336_), .C(_335_), .Y(_338_) );
OR2X2 OR2X2_11 ( .A(gnd), .B(micro_ucr_hash1_a_1__3_), .Y(_339_) );
NAND2X1 NAND2X1_45 ( .A(gnd), .B(micro_ucr_hash1_a_1__3_), .Y(_340_) );
NAND3X1 NAND3X1_28 ( .A(bloque_bytes[75]), .B(_340_), .C(_339_), .Y(_341_) );
AOI21X1 AOI21X1_24 ( .A(_338_), .B(_341_), .C(_327_), .Y(_342_) );
NAND3X1 NAND3X1_29 ( .A(_335_), .B(_340_), .C(_339_), .Y(_343_) );
OAI21X1 OAI21X1_31 ( .A(_337_), .B(_336_), .C(bloque_bytes[75]), .Y(_344_) );
AOI21X1 AOI21X1_25 ( .A(_344_), .B(_343_), .C(_322_), .Y(_345_) );
NOR2X1 NOR2X1_31 ( .A(_342_), .B(_345_), .Y(_237_) );
XOR2X1 XOR2X1_20 ( .A(_334_), .B(_237_), .Y(micro_ucr_hash1_b_3__7_) );
INVX1 INVX1_25 ( .A(bloque_bytes[76]), .Y(_238_) );
OR2X2 OR2X2_12 ( .A(micro_ucr_hash1_b_1__4_), .B(micro_ucr_hash1_a_1__4_), .Y(_239_) );
NAND2X1 NAND2X1_46 ( .A(micro_ucr_hash1_b_1__4_), .B(micro_ucr_hash1_a_1__4_), .Y(_240_) );
NAND3X1 NAND3X1_30 ( .A(_238_), .B(_240_), .C(_239_), .Y(_241_) );
NOR2X1 NOR2X1_32 ( .A(micro_ucr_hash1_b_1__4_), .B(micro_ucr_hash1_a_1__4_), .Y(_242_) );
AND2X2 AND2X2_11 ( .A(micro_ucr_hash1_b_1__4_), .B(micro_ucr_hash1_a_1__4_), .Y(_243_) );
OAI21X1 OAI21X1_32 ( .A(_243_), .B(_242_), .C(bloque_bytes[76]), .Y(_244_) );
NAND3X1 NAND3X1_31 ( .A(_338_), .B(_241_), .C(_244_), .Y(_245_) );
AOI21X1 AOI21X1_26 ( .A(_340_), .B(_339_), .C(bloque_bytes[75]), .Y(_246_) );
OAI21X1 OAI21X1_33 ( .A(_243_), .B(_242_), .C(_238_), .Y(_247_) );
NAND3X1 NAND3X1_32 ( .A(bloque_bytes[76]), .B(_240_), .C(_239_), .Y(_248_) );
NAND3X1 NAND3X1_33 ( .A(_247_), .B(_248_), .C(_246_), .Y(_249_) );
AND2X2 AND2X2_12 ( .A(_249_), .B(_245_), .Y(_250_) );
INVX2 INVX2_15 ( .A(_345_), .Y(_251_) );
NOR2X1 NOR2X1_33 ( .A(_325_), .B(_322_), .Y(_252_) );
AOI21X1 AOI21X1_27 ( .A(_318_), .B(_252_), .C(_342_), .Y(_253_) );
OAI21X1 OAI21X1_34 ( .A(_333_), .B(_317_), .C(_253_), .Y(_254_) );
NAND2X1 NAND2X1_47 ( .A(_251_), .B(_254_), .Y(_255_) );
XNOR2X1 XNOR2X1_17 ( .A(_255_), .B(_250_), .Y(micro_ucr_hash1_c_2__4_) );
NAND2X1 NAND2X1_48 ( .A(_245_), .B(_249_), .Y(_256_) );
OAI21X1 OAI21X1_35 ( .A(_255_), .B(_256_), .C(_245_), .Y(_257_) );
INVX1 INVX1_26 ( .A(bloque_bytes[77]), .Y(_258_) );
OR2X2 OR2X2_13 ( .A(micro_ucr_hash1_b_1__5_), .B(micro_ucr_hash1_a_1__5_), .Y(_259_) );
NAND2X1 NAND2X1_49 ( .A(micro_ucr_hash1_b_1__5_), .B(micro_ucr_hash1_a_1__5_), .Y(_260_) );
NAND3X1 NAND3X1_34 ( .A(_258_), .B(_260_), .C(_259_), .Y(_261_) );
NOR2X1 NOR2X1_34 ( .A(micro_ucr_hash1_b_1__5_), .B(micro_ucr_hash1_a_1__5_), .Y(_262_) );
AND2X2 AND2X2_13 ( .A(micro_ucr_hash1_b_1__5_), .B(micro_ucr_hash1_a_1__5_), .Y(_263_) );
OAI21X1 OAI21X1_36 ( .A(_263_), .B(_262_), .C(bloque_bytes[77]), .Y(_264_) );
NAND3X1 NAND3X1_35 ( .A(_247_), .B(_264_), .C(_261_), .Y(_265_) );
AOI21X1 AOI21X1_28 ( .A(_240_), .B(_239_), .C(bloque_bytes[76]), .Y(_266_) );
NAND3X1 NAND3X1_36 ( .A(bloque_bytes[77]), .B(_260_), .C(_259_), .Y(_267_) );
OAI21X1 OAI21X1_37 ( .A(_263_), .B(_262_), .C(_258_), .Y(_268_) );
NAND3X1 NAND3X1_37 ( .A(_268_), .B(_267_), .C(_266_), .Y(_269_) );
NAND2X1 NAND2X1_50 ( .A(_265_), .B(_269_), .Y(_270_) );
INVX2 INVX2_16 ( .A(_270_), .Y(_271_) );
XNOR2X1 XNOR2X1_18 ( .A(_257_), .B(_271_), .Y(micro_ucr_hash1_c_2__5_) );
AOI21X1 AOI21X1_29 ( .A(_265_), .B(_269_), .C(_256_), .Y(_272_) );
NAND3X1 NAND3X1_38 ( .A(_251_), .B(_272_), .C(_254_), .Y(_273_) );
NAND2X1 NAND2X1_51 ( .A(_268_), .B(_267_), .Y(_274_) );
OR2X2 OR2X2_14 ( .A(_274_), .B(_266_), .Y(_275_) );
INVX1 INVX1_27 ( .A(_275_), .Y(_276_) );
AOI21X1 AOI21X1_30 ( .A(_266_), .B(_274_), .C(_245_), .Y(_277_) );
NOR2X1 NOR2X1_35 ( .A(_277_), .B(_276_), .Y(_278_) );
INVX1 INVX1_28 ( .A(bloque_bytes[78]), .Y(_279_) );
XNOR2X1 XNOR2X1_19 ( .A(micro_ucr_hash1_b_1__6_), .B(micro_ucr_hash1_a_1__6_), .Y(_280_) );
OR2X2 OR2X2_15 ( .A(_280_), .B(_279_), .Y(_281_) );
NAND2X1 NAND2X1_52 ( .A(_279_), .B(_280_), .Y(_282_) );
NAND2X1 NAND2X1_53 ( .A(_282_), .B(_281_), .Y(_283_) );
OR2X2 OR2X2_16 ( .A(_283_), .B(_267_), .Y(_284_) );
NAND2X1 NAND2X1_54 ( .A(_267_), .B(_283_), .Y(_285_) );
NAND2X1 NAND2X1_55 ( .A(_285_), .B(_284_), .Y(_286_) );
AOI21X1 AOI21X1_31 ( .A(_278_), .B(_273_), .C(_286_), .Y(_287_) );
NAND2X1 NAND2X1_56 ( .A(_270_), .B(_250_), .Y(_288_) );
OAI21X1 OAI21X1_38 ( .A(_255_), .B(_288_), .C(_278_), .Y(_289_) );
INVX1 INVX1_29 ( .A(_286_), .Y(_290_) );
NOR2X1 NOR2X1_36 ( .A(_290_), .B(_289_), .Y(_291_) );
NOR2X1 NOR2X1_37 ( .A(_287_), .B(_291_), .Y(micro_ucr_hash1_c_2__6_) );
INVX1 INVX1_30 ( .A(_331_), .Y(_292_) );
AOI21X1 AOI21X1_32 ( .A(_251_), .B(_292_), .C(_342_), .Y(_293_) );
AOI21X1 AOI21X1_33 ( .A(_306_), .B(_307_), .C(_316_), .Y(_294_) );
NAND3X1 NAND3X1_39 ( .A(_294_), .B(_330_), .C(_237_), .Y(_295_) );
AOI21X1 AOI21X1_34 ( .A(_293_), .B(_295_), .C(_288_), .Y(_296_) );
OAI21X1 OAI21X1_39 ( .A(_271_), .B(_245_), .C(_275_), .Y(_297_) );
OAI21X1 OAI21X1_40 ( .A(_296_), .B(_297_), .C(_290_), .Y(_298_) );
XOR2X1 XOR2X1_21 ( .A(micro_ucr_hash1_b_1__7_), .B(bloque_bytes[79]), .Y(_299_) );
XNOR2X1 XNOR2X1_20 ( .A(_299_), .B(micro_ucr_hash1_a_1__7_), .Y(_300_) );
XNOR2X1 XNOR2X1_21 ( .A(_300_), .B(_281_), .Y(_301_) );
NAND3X1 NAND3X1_40 ( .A(_284_), .B(_301_), .C(_298_), .Y(_302_) );
INVX1 INVX1_31 ( .A(_284_), .Y(_303_) );
INVX1 INVX1_32 ( .A(_301_), .Y(_304_) );
OAI21X1 OAI21X1_41 ( .A(_287_), .B(_303_), .C(_304_), .Y(_305_) );
NAND2X1 NAND2X1_57 ( .A(_302_), .B(_305_), .Y(micro_ucr_hash1_c_2__7_) );
XOR2X1 XOR2X1_22 ( .A(micro_ucr_hash1_b_3__4_), .B(gnd), .Y(micro_ucr_hash1_a_3__0_) );
XOR2X1 XOR2X1_23 ( .A(micro_ucr_hash1_b_3__5_), .B(gnd), .Y(micro_ucr_hash1_a_3__1_) );
XOR2X1 XOR2X1_24 ( .A(micro_ucr_hash1_b_3__6_), .B(gnd), .Y(micro_ucr_hash1_a_3__2_) );
XOR2X1 XOR2X1_25 ( .A(micro_ucr_hash1_b_3__7_), .B(gnd), .Y(micro_ucr_hash1_a_3__3_) );
XOR2X1 XOR2X1_26 ( .A(micro_ucr_hash1_c_2__4_), .B(micro_ucr_hash1_b_2__4_), .Y(micro_ucr_hash1_a_3__4_) );
XOR2X1 XOR2X1_27 ( .A(micro_ucr_hash1_c_2__5_), .B(micro_ucr_hash1_b_2__5_), .Y(micro_ucr_hash1_a_3__5_) );
XOR2X1 XOR2X1_28 ( .A(micro_ucr_hash1_c_2__6_), .B(micro_ucr_hash1_b_2__6_), .Y(micro_ucr_hash1_a_3__6_) );
XOR2X1 XOR2X1_29 ( .A(micro_ucr_hash1_c_2__7_), .B(micro_ucr_hash1_b_2__7_), .Y(micro_ucr_hash1_a_3__7_) );
INVX2 INVX2_17 ( .A(bloque_bytes[64]), .Y(_415_) );
XNOR2X1 XNOR2X1_22 ( .A(gnd), .B(micro_ucr_hash1_a_2__0_), .Y(_416_) );
XNOR2X1 XNOR2X1_23 ( .A(_416_), .B(_415_), .Y(micro_ucr_hash1_b_4__4_) );
NAND2X1 NAND2X1_58 ( .A(_415_), .B(_416_), .Y(_417_) );
OR2X2 OR2X2_17 ( .A(gnd), .B(micro_ucr_hash1_a_2__1_), .Y(_418_) );
NAND2X1 NAND2X1_59 ( .A(gnd), .B(micro_ucr_hash1_a_2__1_), .Y(_419_) );
NAND3X1 NAND3X1_41 ( .A(bloque_bytes[65]), .B(_419_), .C(_418_), .Y(_420_) );
INVX1 INVX1_33 ( .A(bloque_bytes[65]), .Y(_421_) );
NOR2X1 NOR2X1_38 ( .A(gnd), .B(micro_ucr_hash1_a_2__1_), .Y(_422_) );
AND2X2 AND2X2_14 ( .A(gnd), .B(micro_ucr_hash1_a_2__1_), .Y(_423_) );
OAI21X1 OAI21X1_42 ( .A(_423_), .B(_422_), .C(_421_), .Y(_424_) );
NAND2X1 NAND2X1_60 ( .A(_424_), .B(_420_), .Y(_425_) );
XNOR2X1 XNOR2X1_24 ( .A(_425_), .B(_417_), .Y(micro_ucr_hash1_b_4__5_) );
NAND3X1 NAND3X1_42 ( .A(_420_), .B(_424_), .C(_417_), .Y(_426_) );
NOR3X1 NOR3X1_29 ( .A(_421_), .B(_422_), .C(_423_), .Y(_427_) );
INVX1 INVX1_34 ( .A(bloque_bytes[66]), .Y(_428_) );
NOR2X1 NOR2X1_39 ( .A(gnd), .B(micro_ucr_hash1_a_2__2_), .Y(_429_) );
AND2X2 AND2X2_15 ( .A(gnd), .B(micro_ucr_hash1_a_2__2_), .Y(_430_) );
NOR3X1 NOR3X1_30 ( .A(_428_), .B(_429_), .C(_430_), .Y(_431_) );
OR2X2 OR2X2_18 ( .A(gnd), .B(micro_ucr_hash1_a_2__2_), .Y(_432_) );
NAND2X1 NAND2X1_61 ( .A(gnd), .B(micro_ucr_hash1_a_2__2_), .Y(_433_) );
AOI21X1 AOI21X1_35 ( .A(_433_), .B(_432_), .C(bloque_bytes[66]), .Y(_434_) );
OAI21X1 OAI21X1_43 ( .A(_431_), .B(_434_), .C(_427_), .Y(_435_) );
NAND3X1 NAND3X1_43 ( .A(bloque_bytes[66]), .B(_433_), .C(_432_), .Y(_436_) );
OAI21X1 OAI21X1_44 ( .A(_430_), .B(_429_), .C(_428_), .Y(_437_) );
NAND3X1 NAND3X1_44 ( .A(_437_), .B(_420_), .C(_436_), .Y(_438_) );
NAND2X1 NAND2X1_62 ( .A(_438_), .B(_435_), .Y(_439_) );
XNOR2X1 XNOR2X1_25 ( .A(_439_), .B(_426_), .Y(micro_ucr_hash1_b_4__6_) );
NAND3X1 NAND3X1_45 ( .A(_436_), .B(_437_), .C(_427_), .Y(_440_) );
OAI21X1 OAI21X1_45 ( .A(_431_), .B(_434_), .C(_420_), .Y(_441_) );
NAND2X1 NAND2X1_63 ( .A(_440_), .B(_441_), .Y(_442_) );
OAI21X1 OAI21X1_46 ( .A(_442_), .B(_426_), .C(_440_), .Y(_443_) );
INVX1 INVX1_35 ( .A(bloque_bytes[67]), .Y(_444_) );
NOR2X1 NOR2X1_40 ( .A(gnd), .B(micro_ucr_hash1_a_2__3_), .Y(_445_) );
AND2X2 AND2X2_16 ( .A(gnd), .B(micro_ucr_hash1_a_2__3_), .Y(_446_) );
OAI21X1 OAI21X1_47 ( .A(_446_), .B(_445_), .C(_444_), .Y(_447_) );
OR2X2 OR2X2_19 ( .A(gnd), .B(micro_ucr_hash1_a_2__3_), .Y(_448_) );
NAND2X1 NAND2X1_64 ( .A(gnd), .B(micro_ucr_hash1_a_2__3_), .Y(_449_) );
NAND3X1 NAND3X1_46 ( .A(bloque_bytes[67]), .B(_449_), .C(_448_), .Y(_450_) );
AOI21X1 AOI21X1_36 ( .A(_447_), .B(_450_), .C(_436_), .Y(_451_) );
NAND3X1 NAND3X1_47 ( .A(_444_), .B(_449_), .C(_448_), .Y(_452_) );
OAI21X1 OAI21X1_48 ( .A(_446_), .B(_445_), .C(bloque_bytes[67]), .Y(_453_) );
AOI21X1 AOI21X1_37 ( .A(_453_), .B(_452_), .C(_431_), .Y(_454_) );
NOR2X1 NOR2X1_41 ( .A(_451_), .B(_454_), .Y(_346_) );
XOR2X1 XOR2X1_30 ( .A(_443_), .B(_346_), .Y(micro_ucr_hash1_b_4__7_) );
INVX1 INVX1_36 ( .A(bloque_bytes[68]), .Y(_347_) );
OR2X2 OR2X2_20 ( .A(micro_ucr_hash1_b_2__4_), .B(micro_ucr_hash1_a_2__4_), .Y(_348_) );
NAND2X1 NAND2X1_65 ( .A(micro_ucr_hash1_b_2__4_), .B(micro_ucr_hash1_a_2__4_), .Y(_349_) );
NAND3X1 NAND3X1_48 ( .A(_347_), .B(_349_), .C(_348_), .Y(_350_) );
NOR2X1 NOR2X1_42 ( .A(micro_ucr_hash1_b_2__4_), .B(micro_ucr_hash1_a_2__4_), .Y(_351_) );
AND2X2 AND2X2_17 ( .A(micro_ucr_hash1_b_2__4_), .B(micro_ucr_hash1_a_2__4_), .Y(_352_) );
OAI21X1 OAI21X1_49 ( .A(_352_), .B(_351_), .C(bloque_bytes[68]), .Y(_353_) );
NAND3X1 NAND3X1_49 ( .A(_447_), .B(_350_), .C(_353_), .Y(_354_) );
AOI21X1 AOI21X1_38 ( .A(_449_), .B(_448_), .C(bloque_bytes[67]), .Y(_355_) );
OAI21X1 OAI21X1_50 ( .A(_352_), .B(_351_), .C(_347_), .Y(_356_) );
NAND3X1 NAND3X1_50 ( .A(bloque_bytes[68]), .B(_349_), .C(_348_), .Y(_357_) );
NAND3X1 NAND3X1_51 ( .A(_356_), .B(_357_), .C(_355_), .Y(_358_) );
AND2X2 AND2X2_18 ( .A(_358_), .B(_354_), .Y(_359_) );
INVX2 INVX2_18 ( .A(_454_), .Y(_360_) );
NOR2X1 NOR2X1_43 ( .A(_434_), .B(_431_), .Y(_361_) );
AOI21X1 AOI21X1_39 ( .A(_427_), .B(_361_), .C(_451_), .Y(_362_) );
OAI21X1 OAI21X1_51 ( .A(_442_), .B(_426_), .C(_362_), .Y(_363_) );
NAND2X1 NAND2X1_66 ( .A(_360_), .B(_363_), .Y(_364_) );
XNOR2X1 XNOR2X1_26 ( .A(_364_), .B(_359_), .Y(micro_ucr_hash1_c_3__4_) );
NAND2X1 NAND2X1_67 ( .A(_354_), .B(_358_), .Y(_365_) );
OAI21X1 OAI21X1_52 ( .A(_364_), .B(_365_), .C(_354_), .Y(_366_) );
INVX1 INVX1_37 ( .A(bloque_bytes[69]), .Y(_367_) );
OR2X2 OR2X2_21 ( .A(micro_ucr_hash1_b_2__5_), .B(micro_ucr_hash1_a_2__5_), .Y(_368_) );
NAND2X1 NAND2X1_68 ( .A(micro_ucr_hash1_b_2__5_), .B(micro_ucr_hash1_a_2__5_), .Y(_369_) );
NAND3X1 NAND3X1_52 ( .A(_367_), .B(_369_), .C(_368_), .Y(_370_) );
NOR2X1 NOR2X1_44 ( .A(micro_ucr_hash1_b_2__5_), .B(micro_ucr_hash1_a_2__5_), .Y(_371_) );
AND2X2 AND2X2_19 ( .A(micro_ucr_hash1_b_2__5_), .B(micro_ucr_hash1_a_2__5_), .Y(_372_) );
OAI21X1 OAI21X1_53 ( .A(_372_), .B(_371_), .C(bloque_bytes[69]), .Y(_373_) );
NAND3X1 NAND3X1_53 ( .A(_356_), .B(_373_), .C(_370_), .Y(_374_) );
AOI21X1 AOI21X1_40 ( .A(_349_), .B(_348_), .C(bloque_bytes[68]), .Y(_375_) );
NAND3X1 NAND3X1_54 ( .A(bloque_bytes[69]), .B(_369_), .C(_368_), .Y(_376_) );
OAI21X1 OAI21X1_54 ( .A(_372_), .B(_371_), .C(_367_), .Y(_377_) );
NAND3X1 NAND3X1_55 ( .A(_377_), .B(_376_), .C(_375_), .Y(_378_) );
NAND2X1 NAND2X1_69 ( .A(_374_), .B(_378_), .Y(_379_) );
INVX2 INVX2_19 ( .A(_379_), .Y(_380_) );
XNOR2X1 XNOR2X1_27 ( .A(_366_), .B(_380_), .Y(micro_ucr_hash1_c_3__5_) );
AOI21X1 AOI21X1_41 ( .A(_374_), .B(_378_), .C(_365_), .Y(_381_) );
NAND3X1 NAND3X1_56 ( .A(_360_), .B(_381_), .C(_363_), .Y(_382_) );
NAND2X1 NAND2X1_70 ( .A(_377_), .B(_376_), .Y(_383_) );
OR2X2 OR2X2_22 ( .A(_383_), .B(_375_), .Y(_384_) );
INVX1 INVX1_38 ( .A(_384_), .Y(_385_) );
AOI21X1 AOI21X1_42 ( .A(_375_), .B(_383_), .C(_354_), .Y(_386_) );
NOR2X1 NOR2X1_45 ( .A(_386_), .B(_385_), .Y(_387_) );
INVX1 INVX1_39 ( .A(bloque_bytes[70]), .Y(_388_) );
XNOR2X1 XNOR2X1_28 ( .A(micro_ucr_hash1_b_2__6_), .B(micro_ucr_hash1_a_2__6_), .Y(_389_) );
OR2X2 OR2X2_23 ( .A(_389_), .B(_388_), .Y(_390_) );
NAND2X1 NAND2X1_71 ( .A(_388_), .B(_389_), .Y(_391_) );
NAND2X1 NAND2X1_72 ( .A(_391_), .B(_390_), .Y(_392_) );
OR2X2 OR2X2_24 ( .A(_392_), .B(_376_), .Y(_393_) );
NAND2X1 NAND2X1_73 ( .A(_376_), .B(_392_), .Y(_394_) );
NAND2X1 NAND2X1_74 ( .A(_394_), .B(_393_), .Y(_395_) );
AOI21X1 AOI21X1_43 ( .A(_387_), .B(_382_), .C(_395_), .Y(_396_) );
NAND2X1 NAND2X1_75 ( .A(_379_), .B(_359_), .Y(_397_) );
OAI21X1 OAI21X1_55 ( .A(_364_), .B(_397_), .C(_387_), .Y(_398_) );
INVX1 INVX1_40 ( .A(_395_), .Y(_399_) );
NOR2X1 NOR2X1_46 ( .A(_399_), .B(_398_), .Y(_400_) );
NOR2X1 NOR2X1_47 ( .A(_396_), .B(_400_), .Y(micro_ucr_hash1_c_3__6_) );
INVX1 INVX1_41 ( .A(_440_), .Y(_401_) );
AOI21X1 AOI21X1_44 ( .A(_360_), .B(_401_), .C(_451_), .Y(_402_) );
AOI21X1 AOI21X1_45 ( .A(_415_), .B(_416_), .C(_425_), .Y(_403_) );
NAND3X1 NAND3X1_57 ( .A(_403_), .B(_439_), .C(_346_), .Y(_404_) );
AOI21X1 AOI21X1_46 ( .A(_402_), .B(_404_), .C(_397_), .Y(_405_) );
OAI21X1 OAI21X1_56 ( .A(_380_), .B(_354_), .C(_384_), .Y(_406_) );
OAI21X1 OAI21X1_57 ( .A(_405_), .B(_406_), .C(_399_), .Y(_407_) );
XOR2X1 XOR2X1_31 ( .A(micro_ucr_hash1_b_2__7_), .B(bloque_bytes[71]), .Y(_408_) );
XNOR2X1 XNOR2X1_29 ( .A(_408_), .B(micro_ucr_hash1_a_2__7_), .Y(_409_) );
XNOR2X1 XNOR2X1_30 ( .A(_409_), .B(_390_), .Y(_410_) );
NAND3X1 NAND3X1_58 ( .A(_393_), .B(_410_), .C(_407_), .Y(_411_) );
INVX1 INVX1_42 ( .A(_393_), .Y(_412_) );
INVX1 INVX1_43 ( .A(_410_), .Y(_413_) );
OAI21X1 OAI21X1_58 ( .A(_396_), .B(_412_), .C(_413_), .Y(_414_) );
NAND2X1 NAND2X1_76 ( .A(_411_), .B(_414_), .Y(micro_ucr_hash1_c_3__7_) );
XOR2X1 XOR2X1_32 ( .A(micro_ucr_hash1_b_4__4_), .B(gnd), .Y(micro_ucr_hash1_a_4__0_) );
XOR2X1 XOR2X1_33 ( .A(micro_ucr_hash1_b_4__5_), .B(gnd), .Y(micro_ucr_hash1_a_4__1_) );
XOR2X1 XOR2X1_34 ( .A(micro_ucr_hash1_b_4__6_), .B(gnd), .Y(micro_ucr_hash1_a_4__2_) );
XOR2X1 XOR2X1_35 ( .A(micro_ucr_hash1_b_4__7_), .B(gnd), .Y(micro_ucr_hash1_a_4__3_) );
XOR2X1 XOR2X1_36 ( .A(micro_ucr_hash1_c_3__4_), .B(micro_ucr_hash1_b_3__4_), .Y(micro_ucr_hash1_a_4__4_) );
XOR2X1 XOR2X1_37 ( .A(micro_ucr_hash1_c_3__5_), .B(micro_ucr_hash1_b_3__5_), .Y(micro_ucr_hash1_a_4__5_) );
XOR2X1 XOR2X1_38 ( .A(micro_ucr_hash1_c_3__6_), .B(micro_ucr_hash1_b_3__6_), .Y(micro_ucr_hash1_a_4__6_) );
XOR2X1 XOR2X1_39 ( .A(micro_ucr_hash1_c_3__7_), .B(micro_ucr_hash1_b_3__7_), .Y(micro_ucr_hash1_a_4__7_) );
INVX2 INVX2_20 ( .A(bloque_bytes[56]), .Y(_524_) );
XNOR2X1 XNOR2X1_31 ( .A(gnd), .B(micro_ucr_hash1_a_3__0_), .Y(_525_) );
XNOR2X1 XNOR2X1_32 ( .A(_525_), .B(_524_), .Y(micro_ucr_hash1_b_5__4_) );
NAND2X1 NAND2X1_77 ( .A(_524_), .B(_525_), .Y(_526_) );
OR2X2 OR2X2_25 ( .A(gnd), .B(micro_ucr_hash1_a_3__1_), .Y(_527_) );
NAND2X1 NAND2X1_78 ( .A(gnd), .B(micro_ucr_hash1_a_3__1_), .Y(_528_) );
NAND3X1 NAND3X1_59 ( .A(bloque_bytes[57]), .B(_528_), .C(_527_), .Y(_529_) );
INVX1 INVX1_44 ( .A(bloque_bytes[57]), .Y(_530_) );
NOR2X1 NOR2X1_48 ( .A(gnd), .B(micro_ucr_hash1_a_3__1_), .Y(_531_) );
AND2X2 AND2X2_20 ( .A(gnd), .B(micro_ucr_hash1_a_3__1_), .Y(_532_) );
OAI21X1 OAI21X1_59 ( .A(_532_), .B(_531_), .C(_530_), .Y(_533_) );
NAND2X1 NAND2X1_79 ( .A(_533_), .B(_529_), .Y(_534_) );
XNOR2X1 XNOR2X1_33 ( .A(_534_), .B(_526_), .Y(micro_ucr_hash1_b_5__5_) );
NAND3X1 NAND3X1_60 ( .A(_529_), .B(_533_), .C(_526_), .Y(_535_) );
NOR3X1 NOR3X1_31 ( .A(_530_), .B(_531_), .C(_532_), .Y(_536_) );
INVX1 INVX1_45 ( .A(bloque_bytes[58]), .Y(_537_) );
NOR2X1 NOR2X1_49 ( .A(gnd), .B(micro_ucr_hash1_a_3__2_), .Y(_538_) );
AND2X2 AND2X2_21 ( .A(gnd), .B(micro_ucr_hash1_a_3__2_), .Y(_539_) );
NOR3X1 NOR3X1_32 ( .A(_537_), .B(_538_), .C(_539_), .Y(_540_) );
OR2X2 OR2X2_26 ( .A(gnd), .B(micro_ucr_hash1_a_3__2_), .Y(_541_) );
NAND2X1 NAND2X1_80 ( .A(gnd), .B(micro_ucr_hash1_a_3__2_), .Y(_542_) );
AOI21X1 AOI21X1_47 ( .A(_542_), .B(_541_), .C(bloque_bytes[58]), .Y(_543_) );
OAI21X1 OAI21X1_60 ( .A(_540_), .B(_543_), .C(_536_), .Y(_544_) );
NAND3X1 NAND3X1_61 ( .A(bloque_bytes[58]), .B(_542_), .C(_541_), .Y(_545_) );
OAI21X1 OAI21X1_61 ( .A(_539_), .B(_538_), .C(_537_), .Y(_546_) );
NAND3X1 NAND3X1_62 ( .A(_546_), .B(_529_), .C(_545_), .Y(_547_) );
NAND2X1 NAND2X1_81 ( .A(_547_), .B(_544_), .Y(_548_) );
XNOR2X1 XNOR2X1_34 ( .A(_548_), .B(_535_), .Y(micro_ucr_hash1_b_5__6_) );
NAND3X1 NAND3X1_63 ( .A(_545_), .B(_546_), .C(_536_), .Y(_549_) );
OAI21X1 OAI21X1_62 ( .A(_540_), .B(_543_), .C(_529_), .Y(_550_) );
NAND2X1 NAND2X1_82 ( .A(_549_), .B(_550_), .Y(_551_) );
OAI21X1 OAI21X1_63 ( .A(_551_), .B(_535_), .C(_549_), .Y(_552_) );
INVX1 INVX1_46 ( .A(bloque_bytes[59]), .Y(_553_) );
NOR2X1 NOR2X1_50 ( .A(gnd), .B(micro_ucr_hash1_a_3__3_), .Y(_554_) );
AND2X2 AND2X2_22 ( .A(gnd), .B(micro_ucr_hash1_a_3__3_), .Y(_555_) );
OAI21X1 OAI21X1_64 ( .A(_555_), .B(_554_), .C(_553_), .Y(_556_) );
OR2X2 OR2X2_27 ( .A(gnd), .B(micro_ucr_hash1_a_3__3_), .Y(_557_) );
NAND2X1 NAND2X1_83 ( .A(gnd), .B(micro_ucr_hash1_a_3__3_), .Y(_558_) );
NAND3X1 NAND3X1_64 ( .A(bloque_bytes[59]), .B(_558_), .C(_557_), .Y(_559_) );
AOI21X1 AOI21X1_48 ( .A(_556_), .B(_559_), .C(_545_), .Y(_560_) );
NAND3X1 NAND3X1_65 ( .A(_553_), .B(_558_), .C(_557_), .Y(_561_) );
OAI21X1 OAI21X1_65 ( .A(_555_), .B(_554_), .C(bloque_bytes[59]), .Y(_562_) );
AOI21X1 AOI21X1_49 ( .A(_562_), .B(_561_), .C(_540_), .Y(_563_) );
NOR2X1 NOR2X1_51 ( .A(_560_), .B(_563_), .Y(_455_) );
XOR2X1 XOR2X1_40 ( .A(_552_), .B(_455_), .Y(micro_ucr_hash1_b_5__7_) );
INVX1 INVX1_47 ( .A(bloque_bytes[60]), .Y(_456_) );
OR2X2 OR2X2_28 ( .A(micro_ucr_hash1_b_3__4_), .B(micro_ucr_hash1_a_3__4_), .Y(_457_) );
NAND2X1 NAND2X1_84 ( .A(micro_ucr_hash1_b_3__4_), .B(micro_ucr_hash1_a_3__4_), .Y(_458_) );
NAND3X1 NAND3X1_66 ( .A(_456_), .B(_458_), .C(_457_), .Y(_459_) );
NOR2X1 NOR2X1_52 ( .A(micro_ucr_hash1_b_3__4_), .B(micro_ucr_hash1_a_3__4_), .Y(_460_) );
AND2X2 AND2X2_23 ( .A(micro_ucr_hash1_b_3__4_), .B(micro_ucr_hash1_a_3__4_), .Y(_461_) );
OAI21X1 OAI21X1_66 ( .A(_461_), .B(_460_), .C(bloque_bytes[60]), .Y(_462_) );
NAND3X1 NAND3X1_67 ( .A(_556_), .B(_459_), .C(_462_), .Y(_463_) );
AOI21X1 AOI21X1_50 ( .A(_558_), .B(_557_), .C(bloque_bytes[59]), .Y(_464_) );
OAI21X1 OAI21X1_67 ( .A(_461_), .B(_460_), .C(_456_), .Y(_465_) );
NAND3X1 NAND3X1_68 ( .A(bloque_bytes[60]), .B(_458_), .C(_457_), .Y(_466_) );
NAND3X1 NAND3X1_69 ( .A(_465_), .B(_466_), .C(_464_), .Y(_467_) );
AND2X2 AND2X2_24 ( .A(_467_), .B(_463_), .Y(_468_) );
INVX2 INVX2_21 ( .A(_563_), .Y(_469_) );
NOR2X1 NOR2X1_53 ( .A(_543_), .B(_540_), .Y(_470_) );
AOI21X1 AOI21X1_51 ( .A(_536_), .B(_470_), .C(_560_), .Y(_471_) );
OAI21X1 OAI21X1_68 ( .A(_551_), .B(_535_), .C(_471_), .Y(_472_) );
NAND2X1 NAND2X1_85 ( .A(_469_), .B(_472_), .Y(_473_) );
XNOR2X1 XNOR2X1_35 ( .A(_473_), .B(_468_), .Y(micro_ucr_hash1_c_4__4_) );
NAND2X1 NAND2X1_86 ( .A(_463_), .B(_467_), .Y(_474_) );
OAI21X1 OAI21X1_69 ( .A(_473_), .B(_474_), .C(_463_), .Y(_475_) );
INVX1 INVX1_48 ( .A(bloque_bytes[61]), .Y(_476_) );
OR2X2 OR2X2_29 ( .A(micro_ucr_hash1_b_3__5_), .B(micro_ucr_hash1_a_3__5_), .Y(_477_) );
NAND2X1 NAND2X1_87 ( .A(micro_ucr_hash1_b_3__5_), .B(micro_ucr_hash1_a_3__5_), .Y(_478_) );
NAND3X1 NAND3X1_70 ( .A(_476_), .B(_478_), .C(_477_), .Y(_479_) );
NOR2X1 NOR2X1_54 ( .A(micro_ucr_hash1_b_3__5_), .B(micro_ucr_hash1_a_3__5_), .Y(_480_) );
AND2X2 AND2X2_25 ( .A(micro_ucr_hash1_b_3__5_), .B(micro_ucr_hash1_a_3__5_), .Y(_481_) );
OAI21X1 OAI21X1_70 ( .A(_481_), .B(_480_), .C(bloque_bytes[61]), .Y(_482_) );
NAND3X1 NAND3X1_71 ( .A(_465_), .B(_482_), .C(_479_), .Y(_483_) );
AOI21X1 AOI21X1_52 ( .A(_458_), .B(_457_), .C(bloque_bytes[60]), .Y(_484_) );
NAND3X1 NAND3X1_72 ( .A(bloque_bytes[61]), .B(_478_), .C(_477_), .Y(_485_) );
OAI21X1 OAI21X1_71 ( .A(_481_), .B(_480_), .C(_476_), .Y(_486_) );
NAND3X1 NAND3X1_73 ( .A(_486_), .B(_485_), .C(_484_), .Y(_487_) );
NAND2X1 NAND2X1_88 ( .A(_483_), .B(_487_), .Y(_488_) );
INVX2 INVX2_22 ( .A(_488_), .Y(_489_) );
XNOR2X1 XNOR2X1_36 ( .A(_475_), .B(_489_), .Y(micro_ucr_hash1_c_4__5_) );
AOI21X1 AOI21X1_53 ( .A(_483_), .B(_487_), .C(_474_), .Y(_490_) );
NAND3X1 NAND3X1_74 ( .A(_469_), .B(_490_), .C(_472_), .Y(_491_) );
NAND2X1 NAND2X1_89 ( .A(_486_), .B(_485_), .Y(_492_) );
OR2X2 OR2X2_30 ( .A(_492_), .B(_484_), .Y(_493_) );
INVX1 INVX1_49 ( .A(_493_), .Y(_494_) );
AOI21X1 AOI21X1_54 ( .A(_484_), .B(_492_), .C(_463_), .Y(_495_) );
NOR2X1 NOR2X1_55 ( .A(_495_), .B(_494_), .Y(_496_) );
INVX1 INVX1_50 ( .A(bloque_bytes[62]), .Y(_497_) );
XNOR2X1 XNOR2X1_37 ( .A(micro_ucr_hash1_b_3__6_), .B(micro_ucr_hash1_a_3__6_), .Y(_498_) );
OR2X2 OR2X2_31 ( .A(_498_), .B(_497_), .Y(_499_) );
NAND2X1 NAND2X1_90 ( .A(_497_), .B(_498_), .Y(_500_) );
NAND2X1 NAND2X1_91 ( .A(_500_), .B(_499_), .Y(_501_) );
OR2X2 OR2X2_32 ( .A(_501_), .B(_485_), .Y(_502_) );
NAND2X1 NAND2X1_92 ( .A(_485_), .B(_501_), .Y(_503_) );
NAND2X1 NAND2X1_93 ( .A(_503_), .B(_502_), .Y(_504_) );
AOI21X1 AOI21X1_55 ( .A(_496_), .B(_491_), .C(_504_), .Y(_505_) );
NAND2X1 NAND2X1_94 ( .A(_488_), .B(_468_), .Y(_506_) );
OAI21X1 OAI21X1_72 ( .A(_473_), .B(_506_), .C(_496_), .Y(_507_) );
INVX1 INVX1_51 ( .A(_504_), .Y(_508_) );
NOR2X1 NOR2X1_56 ( .A(_508_), .B(_507_), .Y(_509_) );
NOR2X1 NOR2X1_57 ( .A(_505_), .B(_509_), .Y(micro_ucr_hash1_c_4__6_) );
INVX1 INVX1_52 ( .A(_549_), .Y(_510_) );
AOI21X1 AOI21X1_56 ( .A(_469_), .B(_510_), .C(_560_), .Y(_511_) );
AOI21X1 AOI21X1_57 ( .A(_524_), .B(_525_), .C(_534_), .Y(_512_) );
NAND3X1 NAND3X1_75 ( .A(_512_), .B(_548_), .C(_455_), .Y(_513_) );
AOI21X1 AOI21X1_58 ( .A(_511_), .B(_513_), .C(_506_), .Y(_514_) );
OAI21X1 OAI21X1_73 ( .A(_489_), .B(_463_), .C(_493_), .Y(_515_) );
OAI21X1 OAI21X1_74 ( .A(_514_), .B(_515_), .C(_508_), .Y(_516_) );
XOR2X1 XOR2X1_41 ( .A(micro_ucr_hash1_b_3__7_), .B(bloque_bytes[63]), .Y(_517_) );
XNOR2X1 XNOR2X1_38 ( .A(_517_), .B(micro_ucr_hash1_a_3__7_), .Y(_518_) );
XNOR2X1 XNOR2X1_39 ( .A(_518_), .B(_499_), .Y(_519_) );
NAND3X1 NAND3X1_76 ( .A(_502_), .B(_519_), .C(_516_), .Y(_520_) );
INVX1 INVX1_53 ( .A(_502_), .Y(_521_) );
INVX1 INVX1_54 ( .A(_519_), .Y(_522_) );
OAI21X1 OAI21X1_75 ( .A(_505_), .B(_521_), .C(_522_), .Y(_523_) );
NAND2X1 NAND2X1_95 ( .A(_520_), .B(_523_), .Y(micro_ucr_hash1_c_4__7_) );
XOR2X1 XOR2X1_42 ( .A(micro_ucr_hash1_b_5__4_), .B(gnd), .Y(micro_ucr_hash1_a_5__0_) );
XOR2X1 XOR2X1_43 ( .A(micro_ucr_hash1_b_5__5_), .B(gnd), .Y(micro_ucr_hash1_a_5__1_) );
XOR2X1 XOR2X1_44 ( .A(micro_ucr_hash1_b_5__6_), .B(gnd), .Y(micro_ucr_hash1_a_5__2_) );
XOR2X1 XOR2X1_45 ( .A(micro_ucr_hash1_b_5__7_), .B(gnd), .Y(micro_ucr_hash1_a_5__3_) );
XOR2X1 XOR2X1_46 ( .A(micro_ucr_hash1_c_4__4_), .B(micro_ucr_hash1_b_4__4_), .Y(micro_ucr_hash1_a_5__4_) );
XOR2X1 XOR2X1_47 ( .A(micro_ucr_hash1_c_4__5_), .B(micro_ucr_hash1_b_4__5_), .Y(micro_ucr_hash1_a_5__5_) );
XOR2X1 XOR2X1_48 ( .A(micro_ucr_hash1_c_4__6_), .B(micro_ucr_hash1_b_4__6_), .Y(micro_ucr_hash1_a_5__6_) );
XOR2X1 XOR2X1_49 ( .A(micro_ucr_hash1_c_4__7_), .B(micro_ucr_hash1_b_4__7_), .Y(micro_ucr_hash1_a_5__7_) );
INVX2 INVX2_23 ( .A(bloque_bytes[48]), .Y(_633_) );
XNOR2X1 XNOR2X1_40 ( .A(gnd), .B(micro_ucr_hash1_a_4__0_), .Y(_634_) );
XNOR2X1 XNOR2X1_41 ( .A(_634_), .B(_633_), .Y(micro_ucr_hash1_b_6__4_) );
NAND2X1 NAND2X1_96 ( .A(_633_), .B(_634_), .Y(_635_) );
OR2X2 OR2X2_33 ( .A(gnd), .B(micro_ucr_hash1_a_4__1_), .Y(_636_) );
NAND2X1 NAND2X1_97 ( .A(gnd), .B(micro_ucr_hash1_a_4__1_), .Y(_637_) );
NAND3X1 NAND3X1_77 ( .A(bloque_bytes[49]), .B(_637_), .C(_636_), .Y(_638_) );
INVX1 INVX1_55 ( .A(bloque_bytes[49]), .Y(_639_) );
NOR2X1 NOR2X1_58 ( .A(gnd), .B(micro_ucr_hash1_a_4__1_), .Y(_640_) );
AND2X2 AND2X2_26 ( .A(gnd), .B(micro_ucr_hash1_a_4__1_), .Y(_641_) );
OAI21X1 OAI21X1_76 ( .A(_641_), .B(_640_), .C(_639_), .Y(_642_) );
NAND2X1 NAND2X1_98 ( .A(_642_), .B(_638_), .Y(_643_) );
XNOR2X1 XNOR2X1_42 ( .A(_643_), .B(_635_), .Y(micro_ucr_hash1_b_6__5_) );
NAND3X1 NAND3X1_78 ( .A(_638_), .B(_642_), .C(_635_), .Y(_644_) );
NOR3X1 NOR3X1_33 ( .A(_639_), .B(_640_), .C(_641_), .Y(_645_) );
INVX1 INVX1_56 ( .A(bloque_bytes[50]), .Y(_646_) );
NOR2X1 NOR2X1_59 ( .A(gnd), .B(micro_ucr_hash1_a_4__2_), .Y(_647_) );
AND2X2 AND2X2_27 ( .A(gnd), .B(micro_ucr_hash1_a_4__2_), .Y(_648_) );
NOR3X1 NOR3X1_34 ( .A(_646_), .B(_647_), .C(_648_), .Y(_649_) );
OR2X2 OR2X2_34 ( .A(gnd), .B(micro_ucr_hash1_a_4__2_), .Y(_650_) );
NAND2X1 NAND2X1_99 ( .A(gnd), .B(micro_ucr_hash1_a_4__2_), .Y(_651_) );
AOI21X1 AOI21X1_59 ( .A(_651_), .B(_650_), .C(bloque_bytes[50]), .Y(_652_) );
OAI21X1 OAI21X1_77 ( .A(_649_), .B(_652_), .C(_645_), .Y(_653_) );
NAND3X1 NAND3X1_79 ( .A(bloque_bytes[50]), .B(_651_), .C(_650_), .Y(_654_) );
OAI21X1 OAI21X1_78 ( .A(_648_), .B(_647_), .C(_646_), .Y(_655_) );
NAND3X1 NAND3X1_80 ( .A(_655_), .B(_638_), .C(_654_), .Y(_656_) );
NAND2X1 NAND2X1_100 ( .A(_656_), .B(_653_), .Y(_657_) );
XNOR2X1 XNOR2X1_43 ( .A(_657_), .B(_644_), .Y(micro_ucr_hash1_b_6__6_) );
NAND3X1 NAND3X1_81 ( .A(_654_), .B(_655_), .C(_645_), .Y(_658_) );
OAI21X1 OAI21X1_79 ( .A(_649_), .B(_652_), .C(_638_), .Y(_659_) );
NAND2X1 NAND2X1_101 ( .A(_658_), .B(_659_), .Y(_660_) );
OAI21X1 OAI21X1_80 ( .A(_660_), .B(_644_), .C(_658_), .Y(_661_) );
INVX1 INVX1_57 ( .A(bloque_bytes[51]), .Y(_662_) );
NOR2X1 NOR2X1_60 ( .A(gnd), .B(micro_ucr_hash1_a_4__3_), .Y(_663_) );
AND2X2 AND2X2_28 ( .A(gnd), .B(micro_ucr_hash1_a_4__3_), .Y(_664_) );
OAI21X1 OAI21X1_81 ( .A(_664_), .B(_663_), .C(_662_), .Y(_665_) );
OR2X2 OR2X2_35 ( .A(gnd), .B(micro_ucr_hash1_a_4__3_), .Y(_666_) );
NAND2X1 NAND2X1_102 ( .A(gnd), .B(micro_ucr_hash1_a_4__3_), .Y(_667_) );
NAND3X1 NAND3X1_82 ( .A(bloque_bytes[51]), .B(_667_), .C(_666_), .Y(_668_) );
AOI21X1 AOI21X1_60 ( .A(_665_), .B(_668_), .C(_654_), .Y(_669_) );
NAND3X1 NAND3X1_83 ( .A(_662_), .B(_667_), .C(_666_), .Y(_670_) );
OAI21X1 OAI21X1_82 ( .A(_664_), .B(_663_), .C(bloque_bytes[51]), .Y(_671_) );
AOI21X1 AOI21X1_61 ( .A(_671_), .B(_670_), .C(_649_), .Y(_672_) );
NOR2X1 NOR2X1_61 ( .A(_669_), .B(_672_), .Y(_564_) );
XOR2X1 XOR2X1_50 ( .A(_661_), .B(_564_), .Y(micro_ucr_hash1_b_6__7_) );
INVX1 INVX1_58 ( .A(bloque_bytes[52]), .Y(_565_) );
OR2X2 OR2X2_36 ( .A(micro_ucr_hash1_b_4__4_), .B(micro_ucr_hash1_a_4__4_), .Y(_566_) );
NAND2X1 NAND2X1_103 ( .A(micro_ucr_hash1_b_4__4_), .B(micro_ucr_hash1_a_4__4_), .Y(_567_) );
NAND3X1 NAND3X1_84 ( .A(_565_), .B(_567_), .C(_566_), .Y(_568_) );
NOR2X1 NOR2X1_62 ( .A(micro_ucr_hash1_b_4__4_), .B(micro_ucr_hash1_a_4__4_), .Y(_569_) );
AND2X2 AND2X2_29 ( .A(micro_ucr_hash1_b_4__4_), .B(micro_ucr_hash1_a_4__4_), .Y(_570_) );
OAI21X1 OAI21X1_83 ( .A(_570_), .B(_569_), .C(bloque_bytes[52]), .Y(_571_) );
NAND3X1 NAND3X1_85 ( .A(_665_), .B(_568_), .C(_571_), .Y(_572_) );
AOI21X1 AOI21X1_62 ( .A(_667_), .B(_666_), .C(bloque_bytes[51]), .Y(_573_) );
OAI21X1 OAI21X1_84 ( .A(_570_), .B(_569_), .C(_565_), .Y(_574_) );
NAND3X1 NAND3X1_86 ( .A(bloque_bytes[52]), .B(_567_), .C(_566_), .Y(_575_) );
NAND3X1 NAND3X1_87 ( .A(_574_), .B(_575_), .C(_573_), .Y(_576_) );
AND2X2 AND2X2_30 ( .A(_576_), .B(_572_), .Y(_577_) );
INVX2 INVX2_24 ( .A(_672_), .Y(_578_) );
NOR2X1 NOR2X1_63 ( .A(_652_), .B(_649_), .Y(_579_) );
AOI21X1 AOI21X1_63 ( .A(_645_), .B(_579_), .C(_669_), .Y(_580_) );
OAI21X1 OAI21X1_85 ( .A(_660_), .B(_644_), .C(_580_), .Y(_581_) );
NAND2X1 NAND2X1_104 ( .A(_578_), .B(_581_), .Y(_582_) );
XNOR2X1 XNOR2X1_44 ( .A(_582_), .B(_577_), .Y(micro_ucr_hash1_c_5__4_) );
NAND2X1 NAND2X1_105 ( .A(_572_), .B(_576_), .Y(_583_) );
OAI21X1 OAI21X1_86 ( .A(_582_), .B(_583_), .C(_572_), .Y(_584_) );
INVX1 INVX1_59 ( .A(bloque_bytes[53]), .Y(_585_) );
OR2X2 OR2X2_37 ( .A(micro_ucr_hash1_b_4__5_), .B(micro_ucr_hash1_a_4__5_), .Y(_586_) );
NAND2X1 NAND2X1_106 ( .A(micro_ucr_hash1_b_4__5_), .B(micro_ucr_hash1_a_4__5_), .Y(_587_) );
NAND3X1 NAND3X1_88 ( .A(_585_), .B(_587_), .C(_586_), .Y(_588_) );
NOR2X1 NOR2X1_64 ( .A(micro_ucr_hash1_b_4__5_), .B(micro_ucr_hash1_a_4__5_), .Y(_589_) );
AND2X2 AND2X2_31 ( .A(micro_ucr_hash1_b_4__5_), .B(micro_ucr_hash1_a_4__5_), .Y(_590_) );
OAI21X1 OAI21X1_87 ( .A(_590_), .B(_589_), .C(bloque_bytes[53]), .Y(_591_) );
NAND3X1 NAND3X1_89 ( .A(_574_), .B(_591_), .C(_588_), .Y(_592_) );
AOI21X1 AOI21X1_64 ( .A(_567_), .B(_566_), .C(bloque_bytes[52]), .Y(_593_) );
NAND3X1 NAND3X1_90 ( .A(bloque_bytes[53]), .B(_587_), .C(_586_), .Y(_594_) );
OAI21X1 OAI21X1_88 ( .A(_590_), .B(_589_), .C(_585_), .Y(_595_) );
NAND3X1 NAND3X1_91 ( .A(_595_), .B(_594_), .C(_593_), .Y(_596_) );
NAND2X1 NAND2X1_107 ( .A(_592_), .B(_596_), .Y(_597_) );
INVX2 INVX2_25 ( .A(_597_), .Y(_598_) );
XNOR2X1 XNOR2X1_45 ( .A(_584_), .B(_598_), .Y(micro_ucr_hash1_c_5__5_) );
AOI21X1 AOI21X1_65 ( .A(_592_), .B(_596_), .C(_583_), .Y(_599_) );
NAND3X1 NAND3X1_92 ( .A(_578_), .B(_599_), .C(_581_), .Y(_600_) );
NAND2X1 NAND2X1_108 ( .A(_595_), .B(_594_), .Y(_601_) );
OR2X2 OR2X2_38 ( .A(_601_), .B(_593_), .Y(_602_) );
INVX1 INVX1_60 ( .A(_602_), .Y(_603_) );
AOI21X1 AOI21X1_66 ( .A(_593_), .B(_601_), .C(_572_), .Y(_604_) );
NOR2X1 NOR2X1_65 ( .A(_604_), .B(_603_), .Y(_605_) );
INVX1 INVX1_61 ( .A(bloque_bytes[54]), .Y(_606_) );
XNOR2X1 XNOR2X1_46 ( .A(micro_ucr_hash1_b_4__6_), .B(micro_ucr_hash1_a_4__6_), .Y(_607_) );
OR2X2 OR2X2_39 ( .A(_607_), .B(_606_), .Y(_608_) );
NAND2X1 NAND2X1_109 ( .A(_606_), .B(_607_), .Y(_609_) );
NAND2X1 NAND2X1_110 ( .A(_609_), .B(_608_), .Y(_610_) );
OR2X2 OR2X2_40 ( .A(_610_), .B(_594_), .Y(_611_) );
NAND2X1 NAND2X1_111 ( .A(_594_), .B(_610_), .Y(_612_) );
NAND2X1 NAND2X1_112 ( .A(_612_), .B(_611_), .Y(_613_) );
AOI21X1 AOI21X1_67 ( .A(_605_), .B(_600_), .C(_613_), .Y(_614_) );
NAND2X1 NAND2X1_113 ( .A(_597_), .B(_577_), .Y(_615_) );
OAI21X1 OAI21X1_89 ( .A(_582_), .B(_615_), .C(_605_), .Y(_616_) );
INVX1 INVX1_62 ( .A(_613_), .Y(_617_) );
NOR2X1 NOR2X1_66 ( .A(_617_), .B(_616_), .Y(_618_) );
NOR2X1 NOR2X1_67 ( .A(_614_), .B(_618_), .Y(micro_ucr_hash1_c_5__6_) );
INVX1 INVX1_63 ( .A(_658_), .Y(_619_) );
AOI21X1 AOI21X1_68 ( .A(_578_), .B(_619_), .C(_669_), .Y(_620_) );
AOI21X1 AOI21X1_69 ( .A(_633_), .B(_634_), .C(_643_), .Y(_621_) );
NAND3X1 NAND3X1_93 ( .A(_621_), .B(_657_), .C(_564_), .Y(_622_) );
AOI21X1 AOI21X1_70 ( .A(_620_), .B(_622_), .C(_615_), .Y(_623_) );
OAI21X1 OAI21X1_90 ( .A(_598_), .B(_572_), .C(_602_), .Y(_624_) );
OAI21X1 OAI21X1_91 ( .A(_623_), .B(_624_), .C(_617_), .Y(_625_) );
XOR2X1 XOR2X1_51 ( .A(micro_ucr_hash1_b_4__7_), .B(bloque_bytes[55]), .Y(_626_) );
XNOR2X1 XNOR2X1_47 ( .A(_626_), .B(micro_ucr_hash1_a_4__7_), .Y(_627_) );
XNOR2X1 XNOR2X1_48 ( .A(_627_), .B(_608_), .Y(_628_) );
NAND3X1 NAND3X1_94 ( .A(_611_), .B(_628_), .C(_625_), .Y(_629_) );
INVX1 INVX1_64 ( .A(_611_), .Y(_630_) );
INVX1 INVX1_65 ( .A(_628_), .Y(_631_) );
OAI21X1 OAI21X1_92 ( .A(_614_), .B(_630_), .C(_631_), .Y(_632_) );
NAND2X1 NAND2X1_114 ( .A(_629_), .B(_632_), .Y(micro_ucr_hash1_c_5__7_) );
XOR2X1 XOR2X1_52 ( .A(micro_ucr_hash1_b_6__4_), .B(gnd), .Y(micro_ucr_hash1_a_6__0_) );
XOR2X1 XOR2X1_53 ( .A(micro_ucr_hash1_b_6__5_), .B(gnd), .Y(micro_ucr_hash1_a_6__1_) );
XOR2X1 XOR2X1_54 ( .A(micro_ucr_hash1_b_6__6_), .B(gnd), .Y(micro_ucr_hash1_a_6__2_) );
XOR2X1 XOR2X1_55 ( .A(micro_ucr_hash1_b_6__7_), .B(gnd), .Y(micro_ucr_hash1_a_6__3_) );
XOR2X1 XOR2X1_56 ( .A(micro_ucr_hash1_c_5__4_), .B(micro_ucr_hash1_b_5__4_), .Y(micro_ucr_hash1_a_6__4_) );
XOR2X1 XOR2X1_57 ( .A(micro_ucr_hash1_c_5__5_), .B(micro_ucr_hash1_b_5__5_), .Y(micro_ucr_hash1_a_6__5_) );
XOR2X1 XOR2X1_58 ( .A(micro_ucr_hash1_c_5__6_), .B(micro_ucr_hash1_b_5__6_), .Y(micro_ucr_hash1_a_6__6_) );
XOR2X1 XOR2X1_59 ( .A(micro_ucr_hash1_c_5__7_), .B(micro_ucr_hash1_b_5__7_), .Y(micro_ucr_hash1_a_6__7_) );
INVX2 INVX2_26 ( .A(bloque_bytes[40]), .Y(_742_) );
XNOR2X1 XNOR2X1_49 ( .A(gnd), .B(micro_ucr_hash1_a_5__0_), .Y(_743_) );
XNOR2X1 XNOR2X1_50 ( .A(_743_), .B(_742_), .Y(micro_ucr_hash1_b_7__4_) );
NAND2X1 NAND2X1_115 ( .A(_742_), .B(_743_), .Y(_744_) );
OR2X2 OR2X2_41 ( .A(gnd), .B(micro_ucr_hash1_a_5__1_), .Y(_745_) );
NAND2X1 NAND2X1_116 ( .A(gnd), .B(micro_ucr_hash1_a_5__1_), .Y(_746_) );
NAND3X1 NAND3X1_95 ( .A(bloque_bytes[41]), .B(_746_), .C(_745_), .Y(_747_) );
INVX1 INVX1_66 ( .A(bloque_bytes[41]), .Y(_748_) );
NOR2X1 NOR2X1_68 ( .A(gnd), .B(micro_ucr_hash1_a_5__1_), .Y(_749_) );
AND2X2 AND2X2_32 ( .A(gnd), .B(micro_ucr_hash1_a_5__1_), .Y(_750_) );
OAI21X1 OAI21X1_93 ( .A(_750_), .B(_749_), .C(_748_), .Y(_751_) );
NAND2X1 NAND2X1_117 ( .A(_751_), .B(_747_), .Y(_752_) );
XNOR2X1 XNOR2X1_51 ( .A(_752_), .B(_744_), .Y(micro_ucr_hash1_b_7__5_) );
NAND3X1 NAND3X1_96 ( .A(_747_), .B(_751_), .C(_744_), .Y(_753_) );
NOR3X1 NOR3X1_35 ( .A(_748_), .B(_749_), .C(_750_), .Y(_754_) );
INVX1 INVX1_67 ( .A(bloque_bytes[42]), .Y(_755_) );
NOR2X1 NOR2X1_69 ( .A(gnd), .B(micro_ucr_hash1_a_5__2_), .Y(_756_) );
AND2X2 AND2X2_33 ( .A(gnd), .B(micro_ucr_hash1_a_5__2_), .Y(_757_) );
NOR3X1 NOR3X1_36 ( .A(_755_), .B(_756_), .C(_757_), .Y(_758_) );
OR2X2 OR2X2_42 ( .A(gnd), .B(micro_ucr_hash1_a_5__2_), .Y(_759_) );
NAND2X1 NAND2X1_118 ( .A(gnd), .B(micro_ucr_hash1_a_5__2_), .Y(_760_) );
AOI21X1 AOI21X1_71 ( .A(_760_), .B(_759_), .C(bloque_bytes[42]), .Y(_761_) );
OAI21X1 OAI21X1_94 ( .A(_758_), .B(_761_), .C(_754_), .Y(_762_) );
NAND3X1 NAND3X1_97 ( .A(bloque_bytes[42]), .B(_760_), .C(_759_), .Y(_763_) );
OAI21X1 OAI21X1_95 ( .A(_757_), .B(_756_), .C(_755_), .Y(_764_) );
NAND3X1 NAND3X1_98 ( .A(_764_), .B(_747_), .C(_763_), .Y(_765_) );
NAND2X1 NAND2X1_119 ( .A(_765_), .B(_762_), .Y(_766_) );
XNOR2X1 XNOR2X1_52 ( .A(_766_), .B(_753_), .Y(micro_ucr_hash1_b_7__6_) );
NAND3X1 NAND3X1_99 ( .A(_763_), .B(_764_), .C(_754_), .Y(_767_) );
OAI21X1 OAI21X1_96 ( .A(_758_), .B(_761_), .C(_747_), .Y(_768_) );
NAND2X1 NAND2X1_120 ( .A(_767_), .B(_768_), .Y(_769_) );
OAI21X1 OAI21X1_97 ( .A(_769_), .B(_753_), .C(_767_), .Y(_770_) );
INVX1 INVX1_68 ( .A(bloque_bytes[43]), .Y(_771_) );
NOR2X1 NOR2X1_70 ( .A(gnd), .B(micro_ucr_hash1_a_5__3_), .Y(_772_) );
AND2X2 AND2X2_34 ( .A(gnd), .B(micro_ucr_hash1_a_5__3_), .Y(_773_) );
OAI21X1 OAI21X1_98 ( .A(_773_), .B(_772_), .C(_771_), .Y(_774_) );
OR2X2 OR2X2_43 ( .A(gnd), .B(micro_ucr_hash1_a_5__3_), .Y(_775_) );
NAND2X1 NAND2X1_121 ( .A(gnd), .B(micro_ucr_hash1_a_5__3_), .Y(_776_) );
NAND3X1 NAND3X1_100 ( .A(bloque_bytes[43]), .B(_776_), .C(_775_), .Y(_777_) );
AOI21X1 AOI21X1_72 ( .A(_774_), .B(_777_), .C(_763_), .Y(_778_) );
NAND3X1 NAND3X1_101 ( .A(_771_), .B(_776_), .C(_775_), .Y(_779_) );
OAI21X1 OAI21X1_99 ( .A(_773_), .B(_772_), .C(bloque_bytes[43]), .Y(_780_) );
AOI21X1 AOI21X1_73 ( .A(_780_), .B(_779_), .C(_758_), .Y(_781_) );
NOR2X1 NOR2X1_71 ( .A(_778_), .B(_781_), .Y(_673_) );
XOR2X1 XOR2X1_60 ( .A(_770_), .B(_673_), .Y(micro_ucr_hash1_b_7__7_) );
INVX1 INVX1_69 ( .A(bloque_bytes[44]), .Y(_674_) );
OR2X2 OR2X2_44 ( .A(micro_ucr_hash1_b_5__4_), .B(micro_ucr_hash1_a_5__4_), .Y(_675_) );
NAND2X1 NAND2X1_122 ( .A(micro_ucr_hash1_b_5__4_), .B(micro_ucr_hash1_a_5__4_), .Y(_676_) );
NAND3X1 NAND3X1_102 ( .A(_674_), .B(_676_), .C(_675_), .Y(_677_) );
NOR2X1 NOR2X1_72 ( .A(micro_ucr_hash1_b_5__4_), .B(micro_ucr_hash1_a_5__4_), .Y(_678_) );
AND2X2 AND2X2_35 ( .A(micro_ucr_hash1_b_5__4_), .B(micro_ucr_hash1_a_5__4_), .Y(_679_) );
OAI21X1 OAI21X1_100 ( .A(_679_), .B(_678_), .C(bloque_bytes[44]), .Y(_680_) );
NAND3X1 NAND3X1_103 ( .A(_774_), .B(_677_), .C(_680_), .Y(_681_) );
AOI21X1 AOI21X1_74 ( .A(_776_), .B(_775_), .C(bloque_bytes[43]), .Y(_682_) );
OAI21X1 OAI21X1_101 ( .A(_679_), .B(_678_), .C(_674_), .Y(_683_) );
NAND3X1 NAND3X1_104 ( .A(bloque_bytes[44]), .B(_676_), .C(_675_), .Y(_684_) );
NAND3X1 NAND3X1_105 ( .A(_683_), .B(_684_), .C(_682_), .Y(_685_) );
AND2X2 AND2X2_36 ( .A(_685_), .B(_681_), .Y(_686_) );
INVX2 INVX2_27 ( .A(_781_), .Y(_687_) );
NOR2X1 NOR2X1_73 ( .A(_761_), .B(_758_), .Y(_688_) );
AOI21X1 AOI21X1_75 ( .A(_754_), .B(_688_), .C(_778_), .Y(_689_) );
OAI21X1 OAI21X1_102 ( .A(_769_), .B(_753_), .C(_689_), .Y(_690_) );
NAND2X1 NAND2X1_123 ( .A(_687_), .B(_690_), .Y(_691_) );
XNOR2X1 XNOR2X1_53 ( .A(_691_), .B(_686_), .Y(micro_ucr_hash1_c_6__4_) );
NAND2X1 NAND2X1_124 ( .A(_681_), .B(_685_), .Y(_692_) );
OAI21X1 OAI21X1_103 ( .A(_691_), .B(_692_), .C(_681_), .Y(_693_) );
INVX1 INVX1_70 ( .A(bloque_bytes[45]), .Y(_694_) );
OR2X2 OR2X2_45 ( .A(micro_ucr_hash1_b_5__5_), .B(micro_ucr_hash1_a_5__5_), .Y(_695_) );
NAND2X1 NAND2X1_125 ( .A(micro_ucr_hash1_b_5__5_), .B(micro_ucr_hash1_a_5__5_), .Y(_696_) );
NAND3X1 NAND3X1_106 ( .A(_694_), .B(_696_), .C(_695_), .Y(_697_) );
NOR2X1 NOR2X1_74 ( .A(micro_ucr_hash1_b_5__5_), .B(micro_ucr_hash1_a_5__5_), .Y(_698_) );
AND2X2 AND2X2_37 ( .A(micro_ucr_hash1_b_5__5_), .B(micro_ucr_hash1_a_5__5_), .Y(_699_) );
OAI21X1 OAI21X1_104 ( .A(_699_), .B(_698_), .C(bloque_bytes[45]), .Y(_700_) );
NAND3X1 NAND3X1_107 ( .A(_683_), .B(_700_), .C(_697_), .Y(_701_) );
AOI21X1 AOI21X1_76 ( .A(_676_), .B(_675_), .C(bloque_bytes[44]), .Y(_702_) );
NAND3X1 NAND3X1_108 ( .A(bloque_bytes[45]), .B(_696_), .C(_695_), .Y(_703_) );
OAI21X1 OAI21X1_105 ( .A(_699_), .B(_698_), .C(_694_), .Y(_704_) );
NAND3X1 NAND3X1_109 ( .A(_704_), .B(_703_), .C(_702_), .Y(_705_) );
NAND2X1 NAND2X1_126 ( .A(_701_), .B(_705_), .Y(_706_) );
INVX2 INVX2_28 ( .A(_706_), .Y(_707_) );
XNOR2X1 XNOR2X1_54 ( .A(_693_), .B(_707_), .Y(micro_ucr_hash1_c_6__5_) );
AOI21X1 AOI21X1_77 ( .A(_701_), .B(_705_), .C(_692_), .Y(_708_) );
NAND3X1 NAND3X1_110 ( .A(_687_), .B(_708_), .C(_690_), .Y(_709_) );
NAND2X1 NAND2X1_127 ( .A(_704_), .B(_703_), .Y(_710_) );
OR2X2 OR2X2_46 ( .A(_710_), .B(_702_), .Y(_711_) );
INVX1 INVX1_71 ( .A(_711_), .Y(_712_) );
AOI21X1 AOI21X1_78 ( .A(_702_), .B(_710_), .C(_681_), .Y(_713_) );
NOR2X1 NOR2X1_75 ( .A(_713_), .B(_712_), .Y(_714_) );
INVX1 INVX1_72 ( .A(bloque_bytes[46]), .Y(_715_) );
XNOR2X1 XNOR2X1_55 ( .A(micro_ucr_hash1_b_5__6_), .B(micro_ucr_hash1_a_5__6_), .Y(_716_) );
OR2X2 OR2X2_47 ( .A(_716_), .B(_715_), .Y(_717_) );
NAND2X1 NAND2X1_128 ( .A(_715_), .B(_716_), .Y(_718_) );
NAND2X1 NAND2X1_129 ( .A(_718_), .B(_717_), .Y(_719_) );
OR2X2 OR2X2_48 ( .A(_719_), .B(_703_), .Y(_720_) );
NAND2X1 NAND2X1_130 ( .A(_703_), .B(_719_), .Y(_721_) );
NAND2X1 NAND2X1_131 ( .A(_721_), .B(_720_), .Y(_722_) );
AOI21X1 AOI21X1_79 ( .A(_714_), .B(_709_), .C(_722_), .Y(_723_) );
NAND2X1 NAND2X1_132 ( .A(_706_), .B(_686_), .Y(_724_) );
OAI21X1 OAI21X1_106 ( .A(_691_), .B(_724_), .C(_714_), .Y(_725_) );
INVX1 INVX1_73 ( .A(_722_), .Y(_726_) );
NOR2X1 NOR2X1_76 ( .A(_726_), .B(_725_), .Y(_727_) );
NOR2X1 NOR2X1_77 ( .A(_723_), .B(_727_), .Y(micro_ucr_hash1_c_6__6_) );
INVX1 INVX1_74 ( .A(_767_), .Y(_728_) );
AOI21X1 AOI21X1_80 ( .A(_687_), .B(_728_), .C(_778_), .Y(_729_) );
AOI21X1 AOI21X1_81 ( .A(_742_), .B(_743_), .C(_752_), .Y(_730_) );
NAND3X1 NAND3X1_111 ( .A(_730_), .B(_766_), .C(_673_), .Y(_731_) );
AOI21X1 AOI21X1_82 ( .A(_729_), .B(_731_), .C(_724_), .Y(_732_) );
OAI21X1 OAI21X1_107 ( .A(_707_), .B(_681_), .C(_711_), .Y(_733_) );
OAI21X1 OAI21X1_108 ( .A(_732_), .B(_733_), .C(_726_), .Y(_734_) );
XOR2X1 XOR2X1_61 ( .A(micro_ucr_hash1_b_5__7_), .B(bloque_bytes[47]), .Y(_735_) );
XNOR2X1 XNOR2X1_56 ( .A(_735_), .B(micro_ucr_hash1_a_5__7_), .Y(_736_) );
XNOR2X1 XNOR2X1_57 ( .A(_736_), .B(_717_), .Y(_737_) );
NAND3X1 NAND3X1_112 ( .A(_720_), .B(_737_), .C(_734_), .Y(_738_) );
INVX1 INVX1_75 ( .A(_720_), .Y(_739_) );
INVX1 INVX1_76 ( .A(_737_), .Y(_740_) );
OAI21X1 OAI21X1_109 ( .A(_723_), .B(_739_), .C(_740_), .Y(_741_) );
NAND2X1 NAND2X1_133 ( .A(_738_), .B(_741_), .Y(micro_ucr_hash1_c_6__7_) );
XOR2X1 XOR2X1_62 ( .A(micro_ucr_hash1_b_7__4_), .B(gnd), .Y(micro_ucr_hash1_a_7__0_) );
XOR2X1 XOR2X1_63 ( .A(micro_ucr_hash1_b_7__5_), .B(gnd), .Y(micro_ucr_hash1_a_7__1_) );
XOR2X1 XOR2X1_64 ( .A(micro_ucr_hash1_b_7__6_), .B(gnd), .Y(micro_ucr_hash1_a_7__2_) );
XOR2X1 XOR2X1_65 ( .A(micro_ucr_hash1_b_7__7_), .B(gnd), .Y(micro_ucr_hash1_a_7__3_) );
XOR2X1 XOR2X1_66 ( .A(micro_ucr_hash1_c_6__4_), .B(micro_ucr_hash1_b_6__4_), .Y(micro_ucr_hash1_a_7__4_) );
XOR2X1 XOR2X1_67 ( .A(micro_ucr_hash1_c_6__5_), .B(micro_ucr_hash1_b_6__5_), .Y(micro_ucr_hash1_a_7__5_) );
XOR2X1 XOR2X1_68 ( .A(micro_ucr_hash1_c_6__6_), .B(micro_ucr_hash1_b_6__6_), .Y(micro_ucr_hash1_a_7__6_) );
XOR2X1 XOR2X1_69 ( .A(micro_ucr_hash1_c_6__7_), .B(micro_ucr_hash1_b_6__7_), .Y(micro_ucr_hash1_a_7__7_) );
INVX2 INVX2_29 ( .A(bloque_bytes[32]), .Y(_851_) );
XNOR2X1 XNOR2X1_58 ( .A(gnd), .B(micro_ucr_hash1_a_6__0_), .Y(_852_) );
XNOR2X1 XNOR2X1_59 ( .A(_852_), .B(_851_), .Y(micro_ucr_hash1_b_8__4_) );
NAND2X1 NAND2X1_134 ( .A(_851_), .B(_852_), .Y(_853_) );
OR2X2 OR2X2_49 ( .A(gnd), .B(micro_ucr_hash1_a_6__1_), .Y(_854_) );
NAND2X1 NAND2X1_135 ( .A(gnd), .B(micro_ucr_hash1_a_6__1_), .Y(_855_) );
NAND3X1 NAND3X1_113 ( .A(bloque_bytes[33]), .B(_855_), .C(_854_), .Y(_856_) );
INVX1 INVX1_77 ( .A(bloque_bytes[33]), .Y(_857_) );
NOR2X1 NOR2X1_78 ( .A(gnd), .B(micro_ucr_hash1_a_6__1_), .Y(_858_) );
AND2X2 AND2X2_38 ( .A(gnd), .B(micro_ucr_hash1_a_6__1_), .Y(_859_) );
OAI21X1 OAI21X1_110 ( .A(_859_), .B(_858_), .C(_857_), .Y(_860_) );
NAND2X1 NAND2X1_136 ( .A(_860_), .B(_856_), .Y(_861_) );
XNOR2X1 XNOR2X1_60 ( .A(_861_), .B(_853_), .Y(micro_ucr_hash1_b_8__5_) );
NAND3X1 NAND3X1_114 ( .A(_856_), .B(_860_), .C(_853_), .Y(_862_) );
NOR3X1 NOR3X1_37 ( .A(_857_), .B(_858_), .C(_859_), .Y(_863_) );
INVX1 INVX1_78 ( .A(bloque_bytes[34]), .Y(_864_) );
NOR2X1 NOR2X1_79 ( .A(gnd), .B(micro_ucr_hash1_a_6__2_), .Y(_865_) );
AND2X2 AND2X2_39 ( .A(gnd), .B(micro_ucr_hash1_a_6__2_), .Y(_866_) );
NOR3X1 NOR3X1_38 ( .A(_864_), .B(_865_), .C(_866_), .Y(_867_) );
OR2X2 OR2X2_50 ( .A(gnd), .B(micro_ucr_hash1_a_6__2_), .Y(_868_) );
NAND2X1 NAND2X1_137 ( .A(gnd), .B(micro_ucr_hash1_a_6__2_), .Y(_869_) );
AOI21X1 AOI21X1_83 ( .A(_869_), .B(_868_), .C(bloque_bytes[34]), .Y(_870_) );
OAI21X1 OAI21X1_111 ( .A(_867_), .B(_870_), .C(_863_), .Y(_871_) );
NAND3X1 NAND3X1_115 ( .A(bloque_bytes[34]), .B(_869_), .C(_868_), .Y(_872_) );
OAI21X1 OAI21X1_112 ( .A(_866_), .B(_865_), .C(_864_), .Y(_873_) );
NAND3X1 NAND3X1_116 ( .A(_873_), .B(_856_), .C(_872_), .Y(_874_) );
NAND2X1 NAND2X1_138 ( .A(_874_), .B(_871_), .Y(_875_) );
XNOR2X1 XNOR2X1_61 ( .A(_875_), .B(_862_), .Y(micro_ucr_hash1_b_8__6_) );
NAND3X1 NAND3X1_117 ( .A(_872_), .B(_873_), .C(_863_), .Y(_876_) );
OAI21X1 OAI21X1_113 ( .A(_867_), .B(_870_), .C(_856_), .Y(_877_) );
NAND2X1 NAND2X1_139 ( .A(_876_), .B(_877_), .Y(_878_) );
OAI21X1 OAI21X1_114 ( .A(_878_), .B(_862_), .C(_876_), .Y(_879_) );
INVX1 INVX1_79 ( .A(bloque_bytes[35]), .Y(_880_) );
NOR2X1 NOR2X1_80 ( .A(gnd), .B(micro_ucr_hash1_a_6__3_), .Y(_881_) );
AND2X2 AND2X2_40 ( .A(gnd), .B(micro_ucr_hash1_a_6__3_), .Y(_882_) );
OAI21X1 OAI21X1_115 ( .A(_882_), .B(_881_), .C(_880_), .Y(_883_) );
OR2X2 OR2X2_51 ( .A(gnd), .B(micro_ucr_hash1_a_6__3_), .Y(_884_) );
NAND2X1 NAND2X1_140 ( .A(gnd), .B(micro_ucr_hash1_a_6__3_), .Y(_885_) );
NAND3X1 NAND3X1_118 ( .A(bloque_bytes[35]), .B(_885_), .C(_884_), .Y(_886_) );
AOI21X1 AOI21X1_84 ( .A(_883_), .B(_886_), .C(_872_), .Y(_887_) );
NAND3X1 NAND3X1_119 ( .A(_880_), .B(_885_), .C(_884_), .Y(_888_) );
OAI21X1 OAI21X1_116 ( .A(_882_), .B(_881_), .C(bloque_bytes[35]), .Y(_889_) );
AOI21X1 AOI21X1_85 ( .A(_889_), .B(_888_), .C(_867_), .Y(_890_) );
NOR2X1 NOR2X1_81 ( .A(_887_), .B(_890_), .Y(_782_) );
XOR2X1 XOR2X1_70 ( .A(_879_), .B(_782_), .Y(micro_ucr_hash1_b_8__7_) );
INVX1 INVX1_80 ( .A(bloque_bytes[36]), .Y(_783_) );
OR2X2 OR2X2_52 ( .A(micro_ucr_hash1_b_6__4_), .B(micro_ucr_hash1_a_6__4_), .Y(_784_) );
NAND2X1 NAND2X1_141 ( .A(micro_ucr_hash1_b_6__4_), .B(micro_ucr_hash1_a_6__4_), .Y(_785_) );
NAND3X1 NAND3X1_120 ( .A(_783_), .B(_785_), .C(_784_), .Y(_786_) );
NOR2X1 NOR2X1_82 ( .A(micro_ucr_hash1_b_6__4_), .B(micro_ucr_hash1_a_6__4_), .Y(_787_) );
AND2X2 AND2X2_41 ( .A(micro_ucr_hash1_b_6__4_), .B(micro_ucr_hash1_a_6__4_), .Y(_788_) );
OAI21X1 OAI21X1_117 ( .A(_788_), .B(_787_), .C(bloque_bytes[36]), .Y(_789_) );
NAND3X1 NAND3X1_121 ( .A(_883_), .B(_786_), .C(_789_), .Y(_790_) );
AOI21X1 AOI21X1_86 ( .A(_885_), .B(_884_), .C(bloque_bytes[35]), .Y(_791_) );
OAI21X1 OAI21X1_118 ( .A(_788_), .B(_787_), .C(_783_), .Y(_792_) );
NAND3X1 NAND3X1_122 ( .A(bloque_bytes[36]), .B(_785_), .C(_784_), .Y(_793_) );
NAND3X1 NAND3X1_123 ( .A(_792_), .B(_793_), .C(_791_), .Y(_794_) );
AND2X2 AND2X2_42 ( .A(_794_), .B(_790_), .Y(_795_) );
INVX2 INVX2_30 ( .A(_890_), .Y(_796_) );
NOR2X1 NOR2X1_83 ( .A(_870_), .B(_867_), .Y(_797_) );
AOI21X1 AOI21X1_87 ( .A(_863_), .B(_797_), .C(_887_), .Y(_798_) );
OAI21X1 OAI21X1_119 ( .A(_878_), .B(_862_), .C(_798_), .Y(_799_) );
NAND2X1 NAND2X1_142 ( .A(_796_), .B(_799_), .Y(_800_) );
XNOR2X1 XNOR2X1_62 ( .A(_800_), .B(_795_), .Y(micro_ucr_hash1_c_7__4_) );
NAND2X1 NAND2X1_143 ( .A(_790_), .B(_794_), .Y(_801_) );
OAI21X1 OAI21X1_120 ( .A(_800_), .B(_801_), .C(_790_), .Y(_802_) );
INVX1 INVX1_81 ( .A(bloque_bytes[37]), .Y(_803_) );
OR2X2 OR2X2_53 ( .A(micro_ucr_hash1_b_6__5_), .B(micro_ucr_hash1_a_6__5_), .Y(_804_) );
NAND2X1 NAND2X1_144 ( .A(micro_ucr_hash1_b_6__5_), .B(micro_ucr_hash1_a_6__5_), .Y(_805_) );
NAND3X1 NAND3X1_124 ( .A(_803_), .B(_805_), .C(_804_), .Y(_806_) );
NOR2X1 NOR2X1_84 ( .A(micro_ucr_hash1_b_6__5_), .B(micro_ucr_hash1_a_6__5_), .Y(_807_) );
AND2X2 AND2X2_43 ( .A(micro_ucr_hash1_b_6__5_), .B(micro_ucr_hash1_a_6__5_), .Y(_808_) );
OAI21X1 OAI21X1_121 ( .A(_808_), .B(_807_), .C(bloque_bytes[37]), .Y(_809_) );
NAND3X1 NAND3X1_125 ( .A(_792_), .B(_809_), .C(_806_), .Y(_810_) );
AOI21X1 AOI21X1_88 ( .A(_785_), .B(_784_), .C(bloque_bytes[36]), .Y(_811_) );
NAND3X1 NAND3X1_126 ( .A(bloque_bytes[37]), .B(_805_), .C(_804_), .Y(_812_) );
OAI21X1 OAI21X1_122 ( .A(_808_), .B(_807_), .C(_803_), .Y(_813_) );
NAND3X1 NAND3X1_127 ( .A(_813_), .B(_812_), .C(_811_), .Y(_814_) );
NAND2X1 NAND2X1_145 ( .A(_810_), .B(_814_), .Y(_815_) );
INVX2 INVX2_31 ( .A(_815_), .Y(_816_) );
XNOR2X1 XNOR2X1_63 ( .A(_802_), .B(_816_), .Y(micro_ucr_hash1_c_7__5_) );
AOI21X1 AOI21X1_89 ( .A(_810_), .B(_814_), .C(_801_), .Y(_817_) );
NAND3X1 NAND3X1_128 ( .A(_796_), .B(_817_), .C(_799_), .Y(_818_) );
NAND2X1 NAND2X1_146 ( .A(_813_), .B(_812_), .Y(_819_) );
OR2X2 OR2X2_54 ( .A(_819_), .B(_811_), .Y(_820_) );
INVX1 INVX1_82 ( .A(_820_), .Y(_821_) );
AOI21X1 AOI21X1_90 ( .A(_811_), .B(_819_), .C(_790_), .Y(_822_) );
NOR2X1 NOR2X1_85 ( .A(_822_), .B(_821_), .Y(_823_) );
INVX1 INVX1_83 ( .A(bloque_bytes[38]), .Y(_824_) );
XNOR2X1 XNOR2X1_64 ( .A(micro_ucr_hash1_b_6__6_), .B(micro_ucr_hash1_a_6__6_), .Y(_825_) );
OR2X2 OR2X2_55 ( .A(_825_), .B(_824_), .Y(_826_) );
NAND2X1 NAND2X1_147 ( .A(_824_), .B(_825_), .Y(_827_) );
NAND2X1 NAND2X1_148 ( .A(_827_), .B(_826_), .Y(_828_) );
OR2X2 OR2X2_56 ( .A(_828_), .B(_812_), .Y(_829_) );
NAND2X1 NAND2X1_149 ( .A(_812_), .B(_828_), .Y(_830_) );
NAND2X1 NAND2X1_150 ( .A(_830_), .B(_829_), .Y(_831_) );
AOI21X1 AOI21X1_91 ( .A(_823_), .B(_818_), .C(_831_), .Y(_832_) );
NAND2X1 NAND2X1_151 ( .A(_815_), .B(_795_), .Y(_833_) );
OAI21X1 OAI21X1_123 ( .A(_800_), .B(_833_), .C(_823_), .Y(_834_) );
INVX1 INVX1_84 ( .A(_831_), .Y(_835_) );
NOR2X1 NOR2X1_86 ( .A(_835_), .B(_834_), .Y(_836_) );
NOR2X1 NOR2X1_87 ( .A(_832_), .B(_836_), .Y(micro_ucr_hash1_c_7__6_) );
INVX1 INVX1_85 ( .A(_876_), .Y(_837_) );
AOI21X1 AOI21X1_92 ( .A(_796_), .B(_837_), .C(_887_), .Y(_838_) );
AOI21X1 AOI21X1_93 ( .A(_851_), .B(_852_), .C(_861_), .Y(_839_) );
NAND3X1 NAND3X1_129 ( .A(_839_), .B(_875_), .C(_782_), .Y(_840_) );
AOI21X1 AOI21X1_94 ( .A(_838_), .B(_840_), .C(_833_), .Y(_841_) );
OAI21X1 OAI21X1_124 ( .A(_816_), .B(_790_), .C(_820_), .Y(_842_) );
OAI21X1 OAI21X1_125 ( .A(_841_), .B(_842_), .C(_835_), .Y(_843_) );
XOR2X1 XOR2X1_71 ( .A(micro_ucr_hash1_b_6__7_), .B(bloque_bytes[39]), .Y(_844_) );
XNOR2X1 XNOR2X1_65 ( .A(_844_), .B(micro_ucr_hash1_a_6__7_), .Y(_845_) );
XNOR2X1 XNOR2X1_66 ( .A(_845_), .B(_826_), .Y(_846_) );
NAND3X1 NAND3X1_130 ( .A(_829_), .B(_846_), .C(_843_), .Y(_847_) );
INVX1 INVX1_86 ( .A(_829_), .Y(_848_) );
INVX1 INVX1_87 ( .A(_846_), .Y(_849_) );
OAI21X1 OAI21X1_126 ( .A(_832_), .B(_848_), .C(_849_), .Y(_850_) );
NAND2X1 NAND2X1_152 ( .A(_847_), .B(_850_), .Y(micro_ucr_hash1_c_7__7_) );
XOR2X1 XOR2X1_72 ( .A(micro_ucr_hash1_b_8__4_), .B(gnd), .Y(micro_ucr_hash1_a_8__0_) );
XOR2X1 XOR2X1_73 ( .A(micro_ucr_hash1_b_8__5_), .B(gnd), .Y(micro_ucr_hash1_a_8__1_) );
XOR2X1 XOR2X1_74 ( .A(micro_ucr_hash1_b_8__6_), .B(gnd), .Y(micro_ucr_hash1_a_8__2_) );
XOR2X1 XOR2X1_75 ( .A(micro_ucr_hash1_b_8__7_), .B(gnd), .Y(micro_ucr_hash1_a_8__3_) );
XOR2X1 XOR2X1_76 ( .A(micro_ucr_hash1_c_7__4_), .B(micro_ucr_hash1_b_7__4_), .Y(micro_ucr_hash1_a_8__4_) );
XOR2X1 XOR2X1_77 ( .A(micro_ucr_hash1_c_7__5_), .B(micro_ucr_hash1_b_7__5_), .Y(micro_ucr_hash1_a_8__5_) );
XOR2X1 XOR2X1_78 ( .A(micro_ucr_hash1_c_7__6_), .B(micro_ucr_hash1_b_7__6_), .Y(micro_ucr_hash1_a_8__6_) );
XOR2X1 XOR2X1_79 ( .A(micro_ucr_hash1_c_7__7_), .B(micro_ucr_hash1_b_7__7_), .Y(micro_ucr_hash1_a_8__7_) );
INVX2 INVX2_32 ( .A(bloque_bytes[24]), .Y(_960_) );
XNOR2X1 XNOR2X1_67 ( .A(gnd), .B(micro_ucr_hash1_a_7__0_), .Y(_961_) );
XNOR2X1 XNOR2X1_68 ( .A(_961_), .B(_960_), .Y(micro_ucr_hash1_b_9__4_) );
NAND2X1 NAND2X1_153 ( .A(_960_), .B(_961_), .Y(_962_) );
OR2X2 OR2X2_57 ( .A(gnd), .B(micro_ucr_hash1_a_7__1_), .Y(_963_) );
NAND2X1 NAND2X1_154 ( .A(gnd), .B(micro_ucr_hash1_a_7__1_), .Y(_964_) );
NAND3X1 NAND3X1_131 ( .A(bloque_bytes[25]), .B(_964_), .C(_963_), .Y(_965_) );
INVX1 INVX1_88 ( .A(bloque_bytes[25]), .Y(_966_) );
NOR2X1 NOR2X1_88 ( .A(gnd), .B(micro_ucr_hash1_a_7__1_), .Y(_967_) );
AND2X2 AND2X2_44 ( .A(gnd), .B(micro_ucr_hash1_a_7__1_), .Y(_968_) );
OAI21X1 OAI21X1_127 ( .A(_968_), .B(_967_), .C(_966_), .Y(_969_) );
NAND2X1 NAND2X1_155 ( .A(_969_), .B(_965_), .Y(_970_) );
XNOR2X1 XNOR2X1_69 ( .A(_970_), .B(_962_), .Y(micro_ucr_hash1_b_9__5_) );
NAND3X1 NAND3X1_132 ( .A(_965_), .B(_969_), .C(_962_), .Y(_971_) );
NOR3X1 NOR3X1_39 ( .A(_966_), .B(_967_), .C(_968_), .Y(_972_) );
INVX1 INVX1_89 ( .A(bloque_bytes[26]), .Y(_973_) );
NOR2X1 NOR2X1_89 ( .A(gnd), .B(micro_ucr_hash1_a_7__2_), .Y(_974_) );
AND2X2 AND2X2_45 ( .A(gnd), .B(micro_ucr_hash1_a_7__2_), .Y(_975_) );
NOR3X1 NOR3X1_40 ( .A(_973_), .B(_974_), .C(_975_), .Y(_976_) );
OR2X2 OR2X2_58 ( .A(gnd), .B(micro_ucr_hash1_a_7__2_), .Y(_977_) );
NAND2X1 NAND2X1_156 ( .A(gnd), .B(micro_ucr_hash1_a_7__2_), .Y(_978_) );
AOI21X1 AOI21X1_95 ( .A(_978_), .B(_977_), .C(bloque_bytes[26]), .Y(_979_) );
OAI21X1 OAI21X1_128 ( .A(_976_), .B(_979_), .C(_972_), .Y(_980_) );
NAND3X1 NAND3X1_133 ( .A(bloque_bytes[26]), .B(_978_), .C(_977_), .Y(_981_) );
OAI21X1 OAI21X1_129 ( .A(_975_), .B(_974_), .C(_973_), .Y(_982_) );
NAND3X1 NAND3X1_134 ( .A(_982_), .B(_965_), .C(_981_), .Y(_983_) );
NAND2X1 NAND2X1_157 ( .A(_983_), .B(_980_), .Y(_984_) );
XNOR2X1 XNOR2X1_70 ( .A(_984_), .B(_971_), .Y(micro_ucr_hash1_b_9__6_) );
NAND3X1 NAND3X1_135 ( .A(_981_), .B(_982_), .C(_972_), .Y(_985_) );
OAI21X1 OAI21X1_130 ( .A(_976_), .B(_979_), .C(_965_), .Y(_986_) );
NAND2X1 NAND2X1_158 ( .A(_985_), .B(_986_), .Y(_987_) );
OAI21X1 OAI21X1_131 ( .A(_987_), .B(_971_), .C(_985_), .Y(_988_) );
INVX1 INVX1_90 ( .A(bloque_bytes[27]), .Y(_989_) );
NOR2X1 NOR2X1_90 ( .A(gnd), .B(micro_ucr_hash1_a_7__3_), .Y(_990_) );
AND2X2 AND2X2_46 ( .A(gnd), .B(micro_ucr_hash1_a_7__3_), .Y(_991_) );
OAI21X1 OAI21X1_132 ( .A(_991_), .B(_990_), .C(_989_), .Y(_992_) );
OR2X2 OR2X2_59 ( .A(gnd), .B(micro_ucr_hash1_a_7__3_), .Y(_993_) );
NAND2X1 NAND2X1_159 ( .A(gnd), .B(micro_ucr_hash1_a_7__3_), .Y(_994_) );
NAND3X1 NAND3X1_136 ( .A(bloque_bytes[27]), .B(_994_), .C(_993_), .Y(_995_) );
AOI21X1 AOI21X1_96 ( .A(_992_), .B(_995_), .C(_981_), .Y(_996_) );
NAND3X1 NAND3X1_137 ( .A(_989_), .B(_994_), .C(_993_), .Y(_997_) );
OAI21X1 OAI21X1_133 ( .A(_991_), .B(_990_), .C(bloque_bytes[27]), .Y(_998_) );
AOI21X1 AOI21X1_97 ( .A(_998_), .B(_997_), .C(_976_), .Y(_999_) );
NOR2X1 NOR2X1_91 ( .A(_996_), .B(_999_), .Y(_891_) );
XOR2X1 XOR2X1_80 ( .A(_988_), .B(_891_), .Y(micro_ucr_hash1_b_9__7_) );
INVX1 INVX1_91 ( .A(bloque_bytes[28]), .Y(_892_) );
OR2X2 OR2X2_60 ( .A(micro_ucr_hash1_b_7__4_), .B(micro_ucr_hash1_a_7__4_), .Y(_893_) );
NAND2X1 NAND2X1_160 ( .A(micro_ucr_hash1_b_7__4_), .B(micro_ucr_hash1_a_7__4_), .Y(_894_) );
NAND3X1 NAND3X1_138 ( .A(_892_), .B(_894_), .C(_893_), .Y(_895_) );
NOR2X1 NOR2X1_92 ( .A(micro_ucr_hash1_b_7__4_), .B(micro_ucr_hash1_a_7__4_), .Y(_896_) );
AND2X2 AND2X2_47 ( .A(micro_ucr_hash1_b_7__4_), .B(micro_ucr_hash1_a_7__4_), .Y(_897_) );
OAI21X1 OAI21X1_134 ( .A(_897_), .B(_896_), .C(bloque_bytes[28]), .Y(_898_) );
NAND3X1 NAND3X1_139 ( .A(_992_), .B(_895_), .C(_898_), .Y(_899_) );
AOI21X1 AOI21X1_98 ( .A(_994_), .B(_993_), .C(bloque_bytes[27]), .Y(_900_) );
OAI21X1 OAI21X1_135 ( .A(_897_), .B(_896_), .C(_892_), .Y(_901_) );
NAND3X1 NAND3X1_140 ( .A(bloque_bytes[28]), .B(_894_), .C(_893_), .Y(_902_) );
NAND3X1 NAND3X1_141 ( .A(_901_), .B(_902_), .C(_900_), .Y(_903_) );
AND2X2 AND2X2_48 ( .A(_903_), .B(_899_), .Y(_904_) );
INVX2 INVX2_33 ( .A(_999_), .Y(_905_) );
NOR2X1 NOR2X1_93 ( .A(_979_), .B(_976_), .Y(_906_) );
AOI21X1 AOI21X1_99 ( .A(_972_), .B(_906_), .C(_996_), .Y(_907_) );
OAI21X1 OAI21X1_136 ( .A(_987_), .B(_971_), .C(_907_), .Y(_908_) );
NAND2X1 NAND2X1_161 ( .A(_905_), .B(_908_), .Y(_909_) );
XNOR2X1 XNOR2X1_71 ( .A(_909_), .B(_904_), .Y(micro_ucr_hash1_c_8__4_) );
NAND2X1 NAND2X1_162 ( .A(_899_), .B(_903_), .Y(_910_) );
OAI21X1 OAI21X1_137 ( .A(_909_), .B(_910_), .C(_899_), .Y(_911_) );
INVX1 INVX1_92 ( .A(bloque_bytes[29]), .Y(_912_) );
OR2X2 OR2X2_61 ( .A(micro_ucr_hash1_b_7__5_), .B(micro_ucr_hash1_a_7__5_), .Y(_913_) );
NAND2X1 NAND2X1_163 ( .A(micro_ucr_hash1_b_7__5_), .B(micro_ucr_hash1_a_7__5_), .Y(_914_) );
NAND3X1 NAND3X1_142 ( .A(_912_), .B(_914_), .C(_913_), .Y(_915_) );
NOR2X1 NOR2X1_94 ( .A(micro_ucr_hash1_b_7__5_), .B(micro_ucr_hash1_a_7__5_), .Y(_916_) );
AND2X2 AND2X2_49 ( .A(micro_ucr_hash1_b_7__5_), .B(micro_ucr_hash1_a_7__5_), .Y(_917_) );
OAI21X1 OAI21X1_138 ( .A(_917_), .B(_916_), .C(bloque_bytes[29]), .Y(_918_) );
NAND3X1 NAND3X1_143 ( .A(_901_), .B(_918_), .C(_915_), .Y(_919_) );
AOI21X1 AOI21X1_100 ( .A(_894_), .B(_893_), .C(bloque_bytes[28]), .Y(_920_) );
NAND3X1 NAND3X1_144 ( .A(bloque_bytes[29]), .B(_914_), .C(_913_), .Y(_921_) );
OAI21X1 OAI21X1_139 ( .A(_917_), .B(_916_), .C(_912_), .Y(_922_) );
NAND3X1 NAND3X1_145 ( .A(_922_), .B(_921_), .C(_920_), .Y(_923_) );
NAND2X1 NAND2X1_164 ( .A(_919_), .B(_923_), .Y(_924_) );
INVX2 INVX2_34 ( .A(_924_), .Y(_925_) );
XNOR2X1 XNOR2X1_72 ( .A(_911_), .B(_925_), .Y(micro_ucr_hash1_c_8__5_) );
AOI21X1 AOI21X1_101 ( .A(_919_), .B(_923_), .C(_910_), .Y(_926_) );
NAND3X1 NAND3X1_146 ( .A(_905_), .B(_926_), .C(_908_), .Y(_927_) );
NAND2X1 NAND2X1_165 ( .A(_922_), .B(_921_), .Y(_928_) );
OR2X2 OR2X2_62 ( .A(_928_), .B(_920_), .Y(_929_) );
INVX1 INVX1_93 ( .A(_929_), .Y(_930_) );
AOI21X1 AOI21X1_102 ( .A(_920_), .B(_928_), .C(_899_), .Y(_931_) );
NOR2X1 NOR2X1_95 ( .A(_931_), .B(_930_), .Y(_932_) );
INVX1 INVX1_94 ( .A(bloque_bytes[30]), .Y(_933_) );
XNOR2X1 XNOR2X1_73 ( .A(micro_ucr_hash1_b_7__6_), .B(micro_ucr_hash1_a_7__6_), .Y(_934_) );
OR2X2 OR2X2_63 ( .A(_934_), .B(_933_), .Y(_935_) );
NAND2X1 NAND2X1_166 ( .A(_933_), .B(_934_), .Y(_936_) );
NAND2X1 NAND2X1_167 ( .A(_936_), .B(_935_), .Y(_937_) );
OR2X2 OR2X2_64 ( .A(_937_), .B(_921_), .Y(_938_) );
NAND2X1 NAND2X1_168 ( .A(_921_), .B(_937_), .Y(_939_) );
NAND2X1 NAND2X1_169 ( .A(_939_), .B(_938_), .Y(_940_) );
AOI21X1 AOI21X1_103 ( .A(_932_), .B(_927_), .C(_940_), .Y(_941_) );
NAND2X1 NAND2X1_170 ( .A(_924_), .B(_904_), .Y(_942_) );
OAI21X1 OAI21X1_140 ( .A(_909_), .B(_942_), .C(_932_), .Y(_943_) );
INVX1 INVX1_95 ( .A(_940_), .Y(_944_) );
NOR2X1 NOR2X1_96 ( .A(_944_), .B(_943_), .Y(_945_) );
NOR2X1 NOR2X1_97 ( .A(_941_), .B(_945_), .Y(micro_ucr_hash1_c_8__6_) );
INVX1 INVX1_96 ( .A(_985_), .Y(_946_) );
AOI21X1 AOI21X1_104 ( .A(_905_), .B(_946_), .C(_996_), .Y(_947_) );
AOI21X1 AOI21X1_105 ( .A(_960_), .B(_961_), .C(_970_), .Y(_948_) );
NAND3X1 NAND3X1_147 ( .A(_948_), .B(_984_), .C(_891_), .Y(_949_) );
AOI21X1 AOI21X1_106 ( .A(_947_), .B(_949_), .C(_942_), .Y(_950_) );
OAI21X1 OAI21X1_141 ( .A(_925_), .B(_899_), .C(_929_), .Y(_951_) );
OAI21X1 OAI21X1_142 ( .A(_950_), .B(_951_), .C(_944_), .Y(_952_) );
XOR2X1 XOR2X1_81 ( .A(micro_ucr_hash1_b_7__7_), .B(bloque_bytes[31]), .Y(_953_) );
XNOR2X1 XNOR2X1_74 ( .A(_953_), .B(micro_ucr_hash1_a_7__7_), .Y(_954_) );
XNOR2X1 XNOR2X1_75 ( .A(_954_), .B(_935_), .Y(_955_) );
NAND3X1 NAND3X1_148 ( .A(_938_), .B(_955_), .C(_952_), .Y(_956_) );
INVX1 INVX1_97 ( .A(_938_), .Y(_957_) );
INVX1 INVX1_98 ( .A(_955_), .Y(_958_) );
OAI21X1 OAI21X1_143 ( .A(_941_), .B(_957_), .C(_958_), .Y(_959_) );
NAND2X1 NAND2X1_171 ( .A(_956_), .B(_959_), .Y(micro_ucr_hash1_c_8__7_) );
XOR2X1 XOR2X1_82 ( .A(micro_ucr_hash1_b_9__4_), .B(gnd), .Y(micro_ucr_hash1_a_9__0_) );
XOR2X1 XOR2X1_83 ( .A(micro_ucr_hash1_b_9__5_), .B(gnd), .Y(micro_ucr_hash1_a_9__1_) );
XOR2X1 XOR2X1_84 ( .A(micro_ucr_hash1_b_9__6_), .B(gnd), .Y(micro_ucr_hash1_a_9__2_) );
XOR2X1 XOR2X1_85 ( .A(micro_ucr_hash1_b_9__7_), .B(gnd), .Y(micro_ucr_hash1_a_9__3_) );
XOR2X1 XOR2X1_86 ( .A(micro_ucr_hash1_c_8__4_), .B(micro_ucr_hash1_b_8__4_), .Y(micro_ucr_hash1_a_9__4_) );
XOR2X1 XOR2X1_87 ( .A(micro_ucr_hash1_c_8__5_), .B(micro_ucr_hash1_b_8__5_), .Y(micro_ucr_hash1_a_9__5_) );
XOR2X1 XOR2X1_88 ( .A(micro_ucr_hash1_c_8__6_), .B(micro_ucr_hash1_b_8__6_), .Y(micro_ucr_hash1_a_9__6_) );
XOR2X1 XOR2X1_89 ( .A(micro_ucr_hash1_c_8__7_), .B(micro_ucr_hash1_b_8__7_), .Y(micro_ucr_hash1_a_9__7_) );
INVX2 INVX2_35 ( .A(bloque_bytes[16]), .Y(_1069_) );
XNOR2X1 XNOR2X1_76 ( .A(gnd), .B(micro_ucr_hash1_a_8__0_), .Y(_1070_) );
XNOR2X1 XNOR2X1_77 ( .A(_1070_), .B(_1069_), .Y(micro_ucr_hash1_b_10__4_) );
NAND2X1 NAND2X1_172 ( .A(_1069_), .B(_1070_), .Y(_1071_) );
OR2X2 OR2X2_65 ( .A(gnd), .B(micro_ucr_hash1_a_8__1_), .Y(_1072_) );
NAND2X1 NAND2X1_173 ( .A(gnd), .B(micro_ucr_hash1_a_8__1_), .Y(_1073_) );
NAND3X1 NAND3X1_149 ( .A(bloque_bytes[17]), .B(_1073_), .C(_1072_), .Y(_1074_) );
INVX1 INVX1_99 ( .A(bloque_bytes[17]), .Y(_1075_) );
NOR2X1 NOR2X1_98 ( .A(gnd), .B(micro_ucr_hash1_a_8__1_), .Y(_1076_) );
AND2X2 AND2X2_50 ( .A(gnd), .B(micro_ucr_hash1_a_8__1_), .Y(_1077_) );
OAI21X1 OAI21X1_144 ( .A(_1077_), .B(_1076_), .C(_1075_), .Y(_1078_) );
NAND2X1 NAND2X1_174 ( .A(_1078_), .B(_1074_), .Y(_1079_) );
XNOR2X1 XNOR2X1_78 ( .A(_1079_), .B(_1071_), .Y(micro_ucr_hash1_b_10__5_) );
NAND3X1 NAND3X1_150 ( .A(_1074_), .B(_1078_), .C(_1071_), .Y(_1080_) );
NOR3X1 NOR3X1_41 ( .A(_1075_), .B(_1076_), .C(_1077_), .Y(_1081_) );
INVX1 INVX1_100 ( .A(bloque_bytes[18]), .Y(_1082_) );
NOR2X1 NOR2X1_99 ( .A(gnd), .B(micro_ucr_hash1_a_8__2_), .Y(_1083_) );
AND2X2 AND2X2_51 ( .A(gnd), .B(micro_ucr_hash1_a_8__2_), .Y(_1084_) );
NOR3X1 NOR3X1_42 ( .A(_1082_), .B(_1083_), .C(_1084_), .Y(_1085_) );
OR2X2 OR2X2_66 ( .A(gnd), .B(micro_ucr_hash1_a_8__2_), .Y(_1086_) );
NAND2X1 NAND2X1_175 ( .A(gnd), .B(micro_ucr_hash1_a_8__2_), .Y(_1087_) );
AOI21X1 AOI21X1_107 ( .A(_1087_), .B(_1086_), .C(bloque_bytes[18]), .Y(_1088_) );
OAI21X1 OAI21X1_145 ( .A(_1085_), .B(_1088_), .C(_1081_), .Y(_1089_) );
NAND3X1 NAND3X1_151 ( .A(bloque_bytes[18]), .B(_1087_), .C(_1086_), .Y(_1090_) );
OAI21X1 OAI21X1_146 ( .A(_1084_), .B(_1083_), .C(_1082_), .Y(_1091_) );
NAND3X1 NAND3X1_152 ( .A(_1091_), .B(_1074_), .C(_1090_), .Y(_1092_) );
NAND2X1 NAND2X1_176 ( .A(_1092_), .B(_1089_), .Y(_1093_) );
XNOR2X1 XNOR2X1_79 ( .A(_1093_), .B(_1080_), .Y(micro_ucr_hash1_b_10__6_) );
NAND3X1 NAND3X1_153 ( .A(_1090_), .B(_1091_), .C(_1081_), .Y(_1094_) );
OAI21X1 OAI21X1_147 ( .A(_1085_), .B(_1088_), .C(_1074_), .Y(_1095_) );
NAND2X1 NAND2X1_177 ( .A(_1094_), .B(_1095_), .Y(_1096_) );
OAI21X1 OAI21X1_148 ( .A(_1096_), .B(_1080_), .C(_1094_), .Y(_1097_) );
INVX1 INVX1_101 ( .A(bloque_bytes[19]), .Y(_1098_) );
NOR2X1 NOR2X1_100 ( .A(gnd), .B(micro_ucr_hash1_a_8__3_), .Y(_1099_) );
AND2X2 AND2X2_52 ( .A(gnd), .B(micro_ucr_hash1_a_8__3_), .Y(_1100_) );
OAI21X1 OAI21X1_149 ( .A(_1100_), .B(_1099_), .C(_1098_), .Y(_1101_) );
OR2X2 OR2X2_67 ( .A(gnd), .B(micro_ucr_hash1_a_8__3_), .Y(_1102_) );
NAND2X1 NAND2X1_178 ( .A(gnd), .B(micro_ucr_hash1_a_8__3_), .Y(_1103_) );
NAND3X1 NAND3X1_154 ( .A(bloque_bytes[19]), .B(_1103_), .C(_1102_), .Y(_1104_) );
AOI21X1 AOI21X1_108 ( .A(_1101_), .B(_1104_), .C(_1090_), .Y(_1105_) );
NAND3X1 NAND3X1_155 ( .A(_1098_), .B(_1103_), .C(_1102_), .Y(_1106_) );
OAI21X1 OAI21X1_150 ( .A(_1100_), .B(_1099_), .C(bloque_bytes[19]), .Y(_1107_) );
AOI21X1 AOI21X1_109 ( .A(_1107_), .B(_1106_), .C(_1085_), .Y(_1108_) );
NOR2X1 NOR2X1_101 ( .A(_1105_), .B(_1108_), .Y(_1000_) );
XOR2X1 XOR2X1_90 ( .A(_1097_), .B(_1000_), .Y(micro_ucr_hash1_b_10__7_) );
INVX1 INVX1_102 ( .A(bloque_bytes[20]), .Y(_1001_) );
OR2X2 OR2X2_68 ( .A(micro_ucr_hash1_b_8__4_), .B(micro_ucr_hash1_a_8__4_), .Y(_1002_) );
NAND2X1 NAND2X1_179 ( .A(micro_ucr_hash1_b_8__4_), .B(micro_ucr_hash1_a_8__4_), .Y(_1003_) );
NAND3X1 NAND3X1_156 ( .A(_1001_), .B(_1003_), .C(_1002_), .Y(_1004_) );
NOR2X1 NOR2X1_102 ( .A(micro_ucr_hash1_b_8__4_), .B(micro_ucr_hash1_a_8__4_), .Y(_1005_) );
AND2X2 AND2X2_53 ( .A(micro_ucr_hash1_b_8__4_), .B(micro_ucr_hash1_a_8__4_), .Y(_1006_) );
OAI21X1 OAI21X1_151 ( .A(_1006_), .B(_1005_), .C(bloque_bytes[20]), .Y(_1007_) );
NAND3X1 NAND3X1_157 ( .A(_1101_), .B(_1004_), .C(_1007_), .Y(_1008_) );
AOI21X1 AOI21X1_110 ( .A(_1103_), .B(_1102_), .C(bloque_bytes[19]), .Y(_1009_) );
OAI21X1 OAI21X1_152 ( .A(_1006_), .B(_1005_), .C(_1001_), .Y(_1010_) );
NAND3X1 NAND3X1_158 ( .A(bloque_bytes[20]), .B(_1003_), .C(_1002_), .Y(_1011_) );
NAND3X1 NAND3X1_159 ( .A(_1010_), .B(_1011_), .C(_1009_), .Y(_1012_) );
AND2X2 AND2X2_54 ( .A(_1012_), .B(_1008_), .Y(_1013_) );
INVX2 INVX2_36 ( .A(_1108_), .Y(_1014_) );
NOR2X1 NOR2X1_103 ( .A(_1088_), .B(_1085_), .Y(_1015_) );
AOI21X1 AOI21X1_111 ( .A(_1081_), .B(_1015_), .C(_1105_), .Y(_1016_) );
OAI21X1 OAI21X1_153 ( .A(_1096_), .B(_1080_), .C(_1016_), .Y(_1017_) );
NAND2X1 NAND2X1_180 ( .A(_1014_), .B(_1017_), .Y(_1018_) );
XNOR2X1 XNOR2X1_80 ( .A(_1018_), .B(_1013_), .Y(micro_ucr_hash1_c_9__4_) );
NAND2X1 NAND2X1_181 ( .A(_1008_), .B(_1012_), .Y(_1019_) );
OAI21X1 OAI21X1_154 ( .A(_1018_), .B(_1019_), .C(_1008_), .Y(_1020_) );
INVX1 INVX1_103 ( .A(bloque_bytes[21]), .Y(_1021_) );
OR2X2 OR2X2_69 ( .A(micro_ucr_hash1_b_8__5_), .B(micro_ucr_hash1_a_8__5_), .Y(_1022_) );
NAND2X1 NAND2X1_182 ( .A(micro_ucr_hash1_b_8__5_), .B(micro_ucr_hash1_a_8__5_), .Y(_1023_) );
NAND3X1 NAND3X1_160 ( .A(_1021_), .B(_1023_), .C(_1022_), .Y(_1024_) );
NOR2X1 NOR2X1_104 ( .A(micro_ucr_hash1_b_8__5_), .B(micro_ucr_hash1_a_8__5_), .Y(_1025_) );
AND2X2 AND2X2_55 ( .A(micro_ucr_hash1_b_8__5_), .B(micro_ucr_hash1_a_8__5_), .Y(_1026_) );
OAI21X1 OAI21X1_155 ( .A(_1026_), .B(_1025_), .C(bloque_bytes[21]), .Y(_1027_) );
NAND3X1 NAND3X1_161 ( .A(_1010_), .B(_1027_), .C(_1024_), .Y(_1028_) );
AOI21X1 AOI21X1_112 ( .A(_1003_), .B(_1002_), .C(bloque_bytes[20]), .Y(_1029_) );
NAND3X1 NAND3X1_162 ( .A(bloque_bytes[21]), .B(_1023_), .C(_1022_), .Y(_1030_) );
OAI21X1 OAI21X1_156 ( .A(_1026_), .B(_1025_), .C(_1021_), .Y(_1031_) );
NAND3X1 NAND3X1_163 ( .A(_1031_), .B(_1030_), .C(_1029_), .Y(_1032_) );
NAND2X1 NAND2X1_183 ( .A(_1028_), .B(_1032_), .Y(_1033_) );
INVX2 INVX2_37 ( .A(_1033_), .Y(_1034_) );
XNOR2X1 XNOR2X1_81 ( .A(_1020_), .B(_1034_), .Y(micro_ucr_hash1_c_9__5_) );
AOI21X1 AOI21X1_113 ( .A(_1028_), .B(_1032_), .C(_1019_), .Y(_1035_) );
NAND3X1 NAND3X1_164 ( .A(_1014_), .B(_1035_), .C(_1017_), .Y(_1036_) );
NAND2X1 NAND2X1_184 ( .A(_1031_), .B(_1030_), .Y(_1037_) );
OR2X2 OR2X2_70 ( .A(_1037_), .B(_1029_), .Y(_1038_) );
INVX1 INVX1_104 ( .A(_1038_), .Y(_1039_) );
AOI21X1 AOI21X1_114 ( .A(_1029_), .B(_1037_), .C(_1008_), .Y(_1040_) );
NOR2X1 NOR2X1_105 ( .A(_1040_), .B(_1039_), .Y(_1041_) );
INVX1 INVX1_105 ( .A(bloque_bytes[22]), .Y(_1042_) );
XNOR2X1 XNOR2X1_82 ( .A(micro_ucr_hash1_b_8__6_), .B(micro_ucr_hash1_a_8__6_), .Y(_1043_) );
OR2X2 OR2X2_71 ( .A(_1043_), .B(_1042_), .Y(_1044_) );
NAND2X1 NAND2X1_185 ( .A(_1042_), .B(_1043_), .Y(_1045_) );
NAND2X1 NAND2X1_186 ( .A(_1045_), .B(_1044_), .Y(_1046_) );
OR2X2 OR2X2_72 ( .A(_1046_), .B(_1030_), .Y(_1047_) );
NAND2X1 NAND2X1_187 ( .A(_1030_), .B(_1046_), .Y(_1048_) );
NAND2X1 NAND2X1_188 ( .A(_1048_), .B(_1047_), .Y(_1049_) );
AOI21X1 AOI21X1_115 ( .A(_1041_), .B(_1036_), .C(_1049_), .Y(_1050_) );
NAND2X1 NAND2X1_189 ( .A(_1033_), .B(_1013_), .Y(_1051_) );
OAI21X1 OAI21X1_157 ( .A(_1018_), .B(_1051_), .C(_1041_), .Y(_1052_) );
INVX1 INVX1_106 ( .A(_1049_), .Y(_1053_) );
NOR2X1 NOR2X1_106 ( .A(_1053_), .B(_1052_), .Y(_1054_) );
NOR2X1 NOR2X1_107 ( .A(_1050_), .B(_1054_), .Y(micro_ucr_hash1_c_9__6_) );
INVX1 INVX1_107 ( .A(_1094_), .Y(_1055_) );
AOI21X1 AOI21X1_116 ( .A(_1014_), .B(_1055_), .C(_1105_), .Y(_1056_) );
AOI21X1 AOI21X1_117 ( .A(_1069_), .B(_1070_), .C(_1079_), .Y(_1057_) );
NAND3X1 NAND3X1_165 ( .A(_1057_), .B(_1093_), .C(_1000_), .Y(_1058_) );
AOI21X1 AOI21X1_118 ( .A(_1056_), .B(_1058_), .C(_1051_), .Y(_1059_) );
OAI21X1 OAI21X1_158 ( .A(_1034_), .B(_1008_), .C(_1038_), .Y(_1060_) );
OAI21X1 OAI21X1_159 ( .A(_1059_), .B(_1060_), .C(_1053_), .Y(_1061_) );
XOR2X1 XOR2X1_91 ( .A(micro_ucr_hash1_b_8__7_), .B(bloque_bytes[23]), .Y(_1062_) );
XNOR2X1 XNOR2X1_83 ( .A(_1062_), .B(micro_ucr_hash1_a_8__7_), .Y(_1063_) );
XNOR2X1 XNOR2X1_84 ( .A(_1063_), .B(_1044_), .Y(_1064_) );
NAND3X1 NAND3X1_166 ( .A(_1047_), .B(_1064_), .C(_1061_), .Y(_1065_) );
INVX1 INVX1_108 ( .A(_1047_), .Y(_1066_) );
INVX1 INVX1_109 ( .A(_1064_), .Y(_1067_) );
OAI21X1 OAI21X1_160 ( .A(_1050_), .B(_1066_), .C(_1067_), .Y(_1068_) );
NAND2X1 NAND2X1_190 ( .A(_1065_), .B(_1068_), .Y(micro_ucr_hash1_c_9__7_) );
XOR2X1 XOR2X1_92 ( .A(micro_ucr_hash1_b_10__4_), .B(gnd), .Y(micro_ucr_hash1_a_10__0_) );
XOR2X1 XOR2X1_93 ( .A(micro_ucr_hash1_b_10__5_), .B(gnd), .Y(micro_ucr_hash1_a_10__1_) );
XOR2X1 XOR2X1_94 ( .A(micro_ucr_hash1_b_10__6_), .B(gnd), .Y(micro_ucr_hash1_a_10__2_) );
XOR2X1 XOR2X1_95 ( .A(micro_ucr_hash1_b_10__7_), .B(gnd), .Y(micro_ucr_hash1_a_10__3_) );
XOR2X1 XOR2X1_96 ( .A(micro_ucr_hash1_c_9__4_), .B(micro_ucr_hash1_b_9__4_), .Y(micro_ucr_hash1_a_10__4_) );
XOR2X1 XOR2X1_97 ( .A(micro_ucr_hash1_c_9__5_), .B(micro_ucr_hash1_b_9__5_), .Y(micro_ucr_hash1_a_10__5_) );
XOR2X1 XOR2X1_98 ( .A(micro_ucr_hash1_c_9__6_), .B(micro_ucr_hash1_b_9__6_), .Y(micro_ucr_hash1_a_10__6_) );
XOR2X1 XOR2X1_99 ( .A(micro_ucr_hash1_c_9__7_), .B(micro_ucr_hash1_b_9__7_), .Y(micro_ucr_hash1_a_10__7_) );
INVX2 INVX2_38 ( .A(bloque_bytes[8]), .Y(_1178_) );
XNOR2X1 XNOR2X1_85 ( .A(gnd), .B(micro_ucr_hash1_a_9__0_), .Y(_1179_) );
XNOR2X1 XNOR2X1_86 ( .A(_1179_), .B(_1178_), .Y(micro_ucr_hash1_b_11__4_) );
NAND2X1 NAND2X1_191 ( .A(_1178_), .B(_1179_), .Y(_1180_) );
OR2X2 OR2X2_73 ( .A(gnd), .B(micro_ucr_hash1_a_9__1_), .Y(_1181_) );
NAND2X1 NAND2X1_192 ( .A(gnd), .B(micro_ucr_hash1_a_9__1_), .Y(_1182_) );
NAND3X1 NAND3X1_167 ( .A(bloque_bytes[9]), .B(_1182_), .C(_1181_), .Y(_1183_) );
INVX1 INVX1_110 ( .A(bloque_bytes[9]), .Y(_1184_) );
NOR2X1 NOR2X1_108 ( .A(gnd), .B(micro_ucr_hash1_a_9__1_), .Y(_1185_) );
AND2X2 AND2X2_56 ( .A(gnd), .B(micro_ucr_hash1_a_9__1_), .Y(_1186_) );
OAI21X1 OAI21X1_161 ( .A(_1186_), .B(_1185_), .C(_1184_), .Y(_1187_) );
NAND2X1 NAND2X1_193 ( .A(_1187_), .B(_1183_), .Y(_1188_) );
XNOR2X1 XNOR2X1_87 ( .A(_1188_), .B(_1180_), .Y(micro_ucr_hash1_b_11__5_) );
NAND3X1 NAND3X1_168 ( .A(_1183_), .B(_1187_), .C(_1180_), .Y(_1189_) );
NOR3X1 NOR3X1_43 ( .A(_1184_), .B(_1185_), .C(_1186_), .Y(_1190_) );
INVX1 INVX1_111 ( .A(bloque_bytes[10]), .Y(_1191_) );
NOR2X1 NOR2X1_109 ( .A(gnd), .B(micro_ucr_hash1_a_9__2_), .Y(_1192_) );
AND2X2 AND2X2_57 ( .A(gnd), .B(micro_ucr_hash1_a_9__2_), .Y(_1193_) );
NOR3X1 NOR3X1_44 ( .A(_1191_), .B(_1192_), .C(_1193_), .Y(_1194_) );
OR2X2 OR2X2_74 ( .A(gnd), .B(micro_ucr_hash1_a_9__2_), .Y(_1195_) );
NAND2X1 NAND2X1_194 ( .A(gnd), .B(micro_ucr_hash1_a_9__2_), .Y(_1196_) );
AOI21X1 AOI21X1_119 ( .A(_1196_), .B(_1195_), .C(bloque_bytes[10]), .Y(_1197_) );
OAI21X1 OAI21X1_162 ( .A(_1194_), .B(_1197_), .C(_1190_), .Y(_1198_) );
NAND3X1 NAND3X1_169 ( .A(bloque_bytes[10]), .B(_1196_), .C(_1195_), .Y(_1199_) );
OAI21X1 OAI21X1_163 ( .A(_1193_), .B(_1192_), .C(_1191_), .Y(_1200_) );
NAND3X1 NAND3X1_170 ( .A(_1200_), .B(_1183_), .C(_1199_), .Y(_1201_) );
NAND2X1 NAND2X1_195 ( .A(_1201_), .B(_1198_), .Y(_1202_) );
XNOR2X1 XNOR2X1_88 ( .A(_1202_), .B(_1189_), .Y(micro_ucr_hash1_b_11__6_) );
NAND3X1 NAND3X1_171 ( .A(_1199_), .B(_1200_), .C(_1190_), .Y(_1203_) );
OAI21X1 OAI21X1_164 ( .A(_1194_), .B(_1197_), .C(_1183_), .Y(_1204_) );
NAND2X1 NAND2X1_196 ( .A(_1203_), .B(_1204_), .Y(_1205_) );
OAI21X1 OAI21X1_165 ( .A(_1205_), .B(_1189_), .C(_1203_), .Y(_1206_) );
INVX1 INVX1_112 ( .A(bloque_bytes[11]), .Y(_1207_) );
NOR2X1 NOR2X1_110 ( .A(gnd), .B(micro_ucr_hash1_a_9__3_), .Y(_1208_) );
AND2X2 AND2X2_58 ( .A(gnd), .B(micro_ucr_hash1_a_9__3_), .Y(_1209_) );
OAI21X1 OAI21X1_166 ( .A(_1209_), .B(_1208_), .C(_1207_), .Y(_1210_) );
OR2X2 OR2X2_75 ( .A(gnd), .B(micro_ucr_hash1_a_9__3_), .Y(_1211_) );
NAND2X1 NAND2X1_197 ( .A(gnd), .B(micro_ucr_hash1_a_9__3_), .Y(_1212_) );
NAND3X1 NAND3X1_172 ( .A(bloque_bytes[11]), .B(_1212_), .C(_1211_), .Y(_1213_) );
AOI21X1 AOI21X1_120 ( .A(_1210_), .B(_1213_), .C(_1199_), .Y(_1214_) );
NAND3X1 NAND3X1_173 ( .A(_1207_), .B(_1212_), .C(_1211_), .Y(_1215_) );
OAI21X1 OAI21X1_167 ( .A(_1209_), .B(_1208_), .C(bloque_bytes[11]), .Y(_1216_) );
AOI21X1 AOI21X1_121 ( .A(_1216_), .B(_1215_), .C(_1194_), .Y(_1217_) );
NOR2X1 NOR2X1_111 ( .A(_1214_), .B(_1217_), .Y(_1109_) );
XOR2X1 XOR2X1_100 ( .A(_1206_), .B(_1109_), .Y(micro_ucr_hash1_b_11__7_) );
INVX1 INVX1_113 ( .A(bloque_bytes[12]), .Y(_1110_) );
OR2X2 OR2X2_76 ( .A(micro_ucr_hash1_b_9__4_), .B(micro_ucr_hash1_a_9__4_), .Y(_1111_) );
NAND2X1 NAND2X1_198 ( .A(micro_ucr_hash1_b_9__4_), .B(micro_ucr_hash1_a_9__4_), .Y(_1112_) );
NAND3X1 NAND3X1_174 ( .A(_1110_), .B(_1112_), .C(_1111_), .Y(_1113_) );
NOR2X1 NOR2X1_112 ( .A(micro_ucr_hash1_b_9__4_), .B(micro_ucr_hash1_a_9__4_), .Y(_1114_) );
AND2X2 AND2X2_59 ( .A(micro_ucr_hash1_b_9__4_), .B(micro_ucr_hash1_a_9__4_), .Y(_1115_) );
OAI21X1 OAI21X1_168 ( .A(_1115_), .B(_1114_), .C(bloque_bytes[12]), .Y(_1116_) );
NAND3X1 NAND3X1_175 ( .A(_1210_), .B(_1113_), .C(_1116_), .Y(_1117_) );
AOI21X1 AOI21X1_122 ( .A(_1212_), .B(_1211_), .C(bloque_bytes[11]), .Y(_1118_) );
OAI21X1 OAI21X1_169 ( .A(_1115_), .B(_1114_), .C(_1110_), .Y(_1119_) );
NAND3X1 NAND3X1_176 ( .A(bloque_bytes[12]), .B(_1112_), .C(_1111_), .Y(_1120_) );
NAND3X1 NAND3X1_177 ( .A(_1119_), .B(_1120_), .C(_1118_), .Y(_1121_) );
AND2X2 AND2X2_60 ( .A(_1121_), .B(_1117_), .Y(_1122_) );
INVX2 INVX2_39 ( .A(_1217_), .Y(_1123_) );
NOR2X1 NOR2X1_113 ( .A(_1197_), .B(_1194_), .Y(_1124_) );
AOI21X1 AOI21X1_123 ( .A(_1190_), .B(_1124_), .C(_1214_), .Y(_1125_) );
OAI21X1 OAI21X1_170 ( .A(_1205_), .B(_1189_), .C(_1125_), .Y(_1126_) );
NAND2X1 NAND2X1_199 ( .A(_1123_), .B(_1126_), .Y(_1127_) );
XNOR2X1 XNOR2X1_89 ( .A(_1127_), .B(_1122_), .Y(micro_ucr_hash1_c_10__4_) );
NAND2X1 NAND2X1_200 ( .A(_1117_), .B(_1121_), .Y(_1128_) );
OAI21X1 OAI21X1_171 ( .A(_1127_), .B(_1128_), .C(_1117_), .Y(_1129_) );
INVX1 INVX1_114 ( .A(bloque_bytes[13]), .Y(_1130_) );
OR2X2 OR2X2_77 ( .A(micro_ucr_hash1_b_9__5_), .B(micro_ucr_hash1_a_9__5_), .Y(_1131_) );
NAND2X1 NAND2X1_201 ( .A(micro_ucr_hash1_b_9__5_), .B(micro_ucr_hash1_a_9__5_), .Y(_1132_) );
NAND3X1 NAND3X1_178 ( .A(_1130_), .B(_1132_), .C(_1131_), .Y(_1133_) );
NOR2X1 NOR2X1_114 ( .A(micro_ucr_hash1_b_9__5_), .B(micro_ucr_hash1_a_9__5_), .Y(_1134_) );
AND2X2 AND2X2_61 ( .A(micro_ucr_hash1_b_9__5_), .B(micro_ucr_hash1_a_9__5_), .Y(_1135_) );
OAI21X1 OAI21X1_172 ( .A(_1135_), .B(_1134_), .C(bloque_bytes[13]), .Y(_1136_) );
NAND3X1 NAND3X1_179 ( .A(_1119_), .B(_1136_), .C(_1133_), .Y(_1137_) );
AOI21X1 AOI21X1_124 ( .A(_1112_), .B(_1111_), .C(bloque_bytes[12]), .Y(_1138_) );
NAND3X1 NAND3X1_180 ( .A(bloque_bytes[13]), .B(_1132_), .C(_1131_), .Y(_1139_) );
OAI21X1 OAI21X1_173 ( .A(_1135_), .B(_1134_), .C(_1130_), .Y(_1140_) );
NAND3X1 NAND3X1_181 ( .A(_1140_), .B(_1139_), .C(_1138_), .Y(_1141_) );
NAND2X1 NAND2X1_202 ( .A(_1137_), .B(_1141_), .Y(_1142_) );
INVX2 INVX2_40 ( .A(_1142_), .Y(_1143_) );
XNOR2X1 XNOR2X1_90 ( .A(_1129_), .B(_1143_), .Y(micro_ucr_hash1_c_10__5_) );
AOI21X1 AOI21X1_125 ( .A(_1137_), .B(_1141_), .C(_1128_), .Y(_1144_) );
NAND3X1 NAND3X1_182 ( .A(_1123_), .B(_1144_), .C(_1126_), .Y(_1145_) );
NAND2X1 NAND2X1_203 ( .A(_1140_), .B(_1139_), .Y(_1146_) );
OR2X2 OR2X2_78 ( .A(_1146_), .B(_1138_), .Y(_1147_) );
INVX1 INVX1_115 ( .A(_1147_), .Y(_1148_) );
AOI21X1 AOI21X1_126 ( .A(_1138_), .B(_1146_), .C(_1117_), .Y(_1149_) );
NOR2X1 NOR2X1_115 ( .A(_1149_), .B(_1148_), .Y(_1150_) );
INVX1 INVX1_116 ( .A(bloque_bytes[14]), .Y(_1151_) );
XNOR2X1 XNOR2X1_91 ( .A(micro_ucr_hash1_b_9__6_), .B(micro_ucr_hash1_a_9__6_), .Y(_1152_) );
OR2X2 OR2X2_79 ( .A(_1152_), .B(_1151_), .Y(_1153_) );
NAND2X1 NAND2X1_204 ( .A(_1151_), .B(_1152_), .Y(_1154_) );
NAND2X1 NAND2X1_205 ( .A(_1154_), .B(_1153_), .Y(_1155_) );
OR2X2 OR2X2_80 ( .A(_1155_), .B(_1139_), .Y(_1156_) );
NAND2X1 NAND2X1_206 ( .A(_1139_), .B(_1155_), .Y(_1157_) );
NAND2X1 NAND2X1_207 ( .A(_1157_), .B(_1156_), .Y(_1158_) );
AOI21X1 AOI21X1_127 ( .A(_1150_), .B(_1145_), .C(_1158_), .Y(_1159_) );
NAND2X1 NAND2X1_208 ( .A(_1142_), .B(_1122_), .Y(_1160_) );
OAI21X1 OAI21X1_174 ( .A(_1127_), .B(_1160_), .C(_1150_), .Y(_1161_) );
INVX1 INVX1_117 ( .A(_1158_), .Y(_1162_) );
NOR2X1 NOR2X1_116 ( .A(_1162_), .B(_1161_), .Y(_1163_) );
NOR2X1 NOR2X1_117 ( .A(_1159_), .B(_1163_), .Y(micro_ucr_hash1_c_10__6_) );
INVX1 INVX1_118 ( .A(_1203_), .Y(_1164_) );
AOI21X1 AOI21X1_128 ( .A(_1123_), .B(_1164_), .C(_1214_), .Y(_1165_) );
AOI21X1 AOI21X1_129 ( .A(_1178_), .B(_1179_), .C(_1188_), .Y(_1166_) );
NAND3X1 NAND3X1_183 ( .A(_1166_), .B(_1202_), .C(_1109_), .Y(_1167_) );
AOI21X1 AOI21X1_130 ( .A(_1165_), .B(_1167_), .C(_1160_), .Y(_1168_) );
OAI21X1 OAI21X1_175 ( .A(_1143_), .B(_1117_), .C(_1147_), .Y(_1169_) );
OAI21X1 OAI21X1_176 ( .A(_1168_), .B(_1169_), .C(_1162_), .Y(_1170_) );
XOR2X1 XOR2X1_101 ( .A(micro_ucr_hash1_b_9__7_), .B(bloque_bytes[15]), .Y(_1171_) );
XNOR2X1 XNOR2X1_92 ( .A(_1171_), .B(micro_ucr_hash1_a_9__7_), .Y(_1172_) );
XNOR2X1 XNOR2X1_93 ( .A(_1172_), .B(_1153_), .Y(_1173_) );
NAND3X1 NAND3X1_184 ( .A(_1156_), .B(_1173_), .C(_1170_), .Y(_1174_) );
INVX1 INVX1_119 ( .A(_1156_), .Y(_1175_) );
INVX1 INVX1_120 ( .A(_1173_), .Y(_1176_) );
OAI21X1 OAI21X1_177 ( .A(_1159_), .B(_1175_), .C(_1176_), .Y(_1177_) );
NAND2X1 NAND2X1_209 ( .A(_1174_), .B(_1177_), .Y(micro_ucr_hash1_c_10__7_) );
XOR2X1 XOR2X1_102 ( .A(micro_ucr_hash1_b_11__4_), .B(gnd), .Y(micro_ucr_hash1_a_11__0_) );
XOR2X1 XOR2X1_103 ( .A(micro_ucr_hash1_b_11__5_), .B(gnd), .Y(micro_ucr_hash1_a_11__1_) );
XOR2X1 XOR2X1_104 ( .A(micro_ucr_hash1_b_11__6_), .B(gnd), .Y(micro_ucr_hash1_a_11__2_) );
XOR2X1 XOR2X1_105 ( .A(micro_ucr_hash1_b_11__7_), .B(gnd), .Y(micro_ucr_hash1_a_11__3_) );
XOR2X1 XOR2X1_106 ( .A(micro_ucr_hash1_c_10__4_), .B(micro_ucr_hash1_b_10__4_), .Y(micro_ucr_hash1_a_11__4_) );
XOR2X1 XOR2X1_107 ( .A(micro_ucr_hash1_c_10__5_), .B(micro_ucr_hash1_b_10__5_), .Y(micro_ucr_hash1_a_11__5_) );
XOR2X1 XOR2X1_108 ( .A(micro_ucr_hash1_c_10__6_), .B(micro_ucr_hash1_b_10__6_), .Y(micro_ucr_hash1_a_11__6_) );
XOR2X1 XOR2X1_109 ( .A(micro_ucr_hash1_c_10__7_), .B(micro_ucr_hash1_b_10__7_), .Y(micro_ucr_hash1_a_11__7_) );
INVX2 INVX2_41 ( .A(bloque_bytes[0]), .Y(_1287_) );
XNOR2X1 XNOR2X1_94 ( .A(gnd), .B(micro_ucr_hash1_a_10__0_), .Y(_1288_) );
XNOR2X1 XNOR2X1_95 ( .A(_1288_), .B(_1287_), .Y(micro_ucr_hash1_b_12__4_) );
NAND2X1 NAND2X1_210 ( .A(_1287_), .B(_1288_), .Y(_1289_) );
OR2X2 OR2X2_81 ( .A(gnd), .B(micro_ucr_hash1_a_10__1_), .Y(_1290_) );
NAND2X1 NAND2X1_211 ( .A(gnd), .B(micro_ucr_hash1_a_10__1_), .Y(_1291_) );
NAND3X1 NAND3X1_185 ( .A(bloque_bytes[1]), .B(_1291_), .C(_1290_), .Y(_1292_) );
INVX1 INVX1_121 ( .A(bloque_bytes[1]), .Y(_1293_) );
NOR2X1 NOR2X1_118 ( .A(gnd), .B(micro_ucr_hash1_a_10__1_), .Y(_1294_) );
AND2X2 AND2X2_62 ( .A(gnd), .B(micro_ucr_hash1_a_10__1_), .Y(_1295_) );
OAI21X1 OAI21X1_178 ( .A(_1295_), .B(_1294_), .C(_1293_), .Y(_1296_) );
NAND2X1 NAND2X1_212 ( .A(_1296_), .B(_1292_), .Y(_1297_) );
XNOR2X1 XNOR2X1_96 ( .A(_1297_), .B(_1289_), .Y(micro_ucr_hash1_b_12__5_) );
NAND3X1 NAND3X1_186 ( .A(_1292_), .B(_1296_), .C(_1289_), .Y(_1298_) );
NOR3X1 NOR3X1_45 ( .A(_1293_), .B(_1294_), .C(_1295_), .Y(_1299_) );
INVX1 INVX1_122 ( .A(bloque_bytes[2]), .Y(_1300_) );
NOR2X1 NOR2X1_119 ( .A(gnd), .B(micro_ucr_hash1_a_10__2_), .Y(_1301_) );
AND2X2 AND2X2_63 ( .A(gnd), .B(micro_ucr_hash1_a_10__2_), .Y(_1302_) );
NOR3X1 NOR3X1_46 ( .A(_1300_), .B(_1301_), .C(_1302_), .Y(_1303_) );
OR2X2 OR2X2_82 ( .A(gnd), .B(micro_ucr_hash1_a_10__2_), .Y(_1304_) );
NAND2X1 NAND2X1_213 ( .A(gnd), .B(micro_ucr_hash1_a_10__2_), .Y(_1305_) );
AOI21X1 AOI21X1_131 ( .A(_1305_), .B(_1304_), .C(bloque_bytes[2]), .Y(_1306_) );
OAI21X1 OAI21X1_179 ( .A(_1303_), .B(_1306_), .C(_1299_), .Y(_1307_) );
NAND3X1 NAND3X1_187 ( .A(bloque_bytes[2]), .B(_1305_), .C(_1304_), .Y(_1308_) );
OAI21X1 OAI21X1_180 ( .A(_1302_), .B(_1301_), .C(_1300_), .Y(_1309_) );
NAND3X1 NAND3X1_188 ( .A(_1309_), .B(_1292_), .C(_1308_), .Y(_1310_) );
NAND2X1 NAND2X1_214 ( .A(_1310_), .B(_1307_), .Y(_1311_) );
XNOR2X1 XNOR2X1_97 ( .A(_1311_), .B(_1298_), .Y(micro_ucr_hash1_b_12__6_) );
NAND3X1 NAND3X1_189 ( .A(_1308_), .B(_1309_), .C(_1299_), .Y(_1312_) );
OAI21X1 OAI21X1_181 ( .A(_1303_), .B(_1306_), .C(_1292_), .Y(_1313_) );
NAND2X1 NAND2X1_215 ( .A(_1312_), .B(_1313_), .Y(_1314_) );
OAI21X1 OAI21X1_182 ( .A(_1314_), .B(_1298_), .C(_1312_), .Y(_1315_) );
INVX1 INVX1_123 ( .A(bloque_bytes[3]), .Y(_1316_) );
NOR2X1 NOR2X1_120 ( .A(gnd), .B(micro_ucr_hash1_a_10__3_), .Y(_1317_) );
AND2X2 AND2X2_64 ( .A(gnd), .B(micro_ucr_hash1_a_10__3_), .Y(_1318_) );
OAI21X1 OAI21X1_183 ( .A(_1318_), .B(_1317_), .C(_1316_), .Y(_1319_) );
OR2X2 OR2X2_83 ( .A(gnd), .B(micro_ucr_hash1_a_10__3_), .Y(_1320_) );
NAND2X1 NAND2X1_216 ( .A(gnd), .B(micro_ucr_hash1_a_10__3_), .Y(_1321_) );
NAND3X1 NAND3X1_190 ( .A(bloque_bytes[3]), .B(_1321_), .C(_1320_), .Y(_1322_) );
AOI21X1 AOI21X1_132 ( .A(_1319_), .B(_1322_), .C(_1308_), .Y(_1323_) );
NAND3X1 NAND3X1_191 ( .A(_1316_), .B(_1321_), .C(_1320_), .Y(_1324_) );
OAI21X1 OAI21X1_184 ( .A(_1318_), .B(_1317_), .C(bloque_bytes[3]), .Y(_1325_) );
AOI21X1 AOI21X1_133 ( .A(_1325_), .B(_1324_), .C(_1303_), .Y(_1326_) );
NOR2X1 NOR2X1_121 ( .A(_1323_), .B(_1326_), .Y(_1218_) );
XOR2X1 XOR2X1_110 ( .A(_1315_), .B(_1218_), .Y(micro_ucr_hash1_b_12__7_) );
INVX1 INVX1_124 ( .A(bloque_bytes[4]), .Y(_1219_) );
OR2X2 OR2X2_84 ( .A(micro_ucr_hash1_b_10__4_), .B(micro_ucr_hash1_a_10__4_), .Y(_1220_) );
NAND2X1 NAND2X1_217 ( .A(micro_ucr_hash1_b_10__4_), .B(micro_ucr_hash1_a_10__4_), .Y(_1221_) );
NAND3X1 NAND3X1_192 ( .A(_1219_), .B(_1221_), .C(_1220_), .Y(_1222_) );
NOR2X1 NOR2X1_122 ( .A(micro_ucr_hash1_b_10__4_), .B(micro_ucr_hash1_a_10__4_), .Y(_1223_) );
AND2X2 AND2X2_65 ( .A(micro_ucr_hash1_b_10__4_), .B(micro_ucr_hash1_a_10__4_), .Y(_1224_) );
OAI21X1 OAI21X1_185 ( .A(_1224_), .B(_1223_), .C(bloque_bytes[4]), .Y(_1225_) );
NAND3X1 NAND3X1_193 ( .A(_1319_), .B(_1222_), .C(_1225_), .Y(_1226_) );
AOI21X1 AOI21X1_134 ( .A(_1321_), .B(_1320_), .C(bloque_bytes[3]), .Y(_1227_) );
OAI21X1 OAI21X1_186 ( .A(_1224_), .B(_1223_), .C(_1219_), .Y(_1228_) );
NAND3X1 NAND3X1_194 ( .A(bloque_bytes[4]), .B(_1221_), .C(_1220_), .Y(_1229_) );
NAND3X1 NAND3X1_195 ( .A(_1228_), .B(_1229_), .C(_1227_), .Y(_1230_) );
AND2X2 AND2X2_66 ( .A(_1230_), .B(_1226_), .Y(_1231_) );
INVX2 INVX2_42 ( .A(_1326_), .Y(_1232_) );
NOR2X1 NOR2X1_123 ( .A(_1306_), .B(_1303_), .Y(_1233_) );
AOI21X1 AOI21X1_135 ( .A(_1299_), .B(_1233_), .C(_1323_), .Y(_1234_) );
OAI21X1 OAI21X1_187 ( .A(_1314_), .B(_1298_), .C(_1234_), .Y(_1235_) );
NAND2X1 NAND2X1_218 ( .A(_1232_), .B(_1235_), .Y(_1236_) );
XNOR2X1 XNOR2X1_98 ( .A(_1236_), .B(_1231_), .Y(micro_ucr_hash1_c_11__4_) );
NAND2X1 NAND2X1_219 ( .A(_1226_), .B(_1230_), .Y(_1237_) );
OAI21X1 OAI21X1_188 ( .A(_1236_), .B(_1237_), .C(_1226_), .Y(_1238_) );
INVX1 INVX1_125 ( .A(bloque_bytes[5]), .Y(_1239_) );
OR2X2 OR2X2_85 ( .A(micro_ucr_hash1_b_10__5_), .B(micro_ucr_hash1_a_10__5_), .Y(_1240_) );
NAND2X1 NAND2X1_220 ( .A(micro_ucr_hash1_b_10__5_), .B(micro_ucr_hash1_a_10__5_), .Y(_1241_) );
NAND3X1 NAND3X1_196 ( .A(_1239_), .B(_1241_), .C(_1240_), .Y(_1242_) );
NOR2X1 NOR2X1_124 ( .A(micro_ucr_hash1_b_10__5_), .B(micro_ucr_hash1_a_10__5_), .Y(_1243_) );
AND2X2 AND2X2_67 ( .A(micro_ucr_hash1_b_10__5_), .B(micro_ucr_hash1_a_10__5_), .Y(_1244_) );
OAI21X1 OAI21X1_189 ( .A(_1244_), .B(_1243_), .C(bloque_bytes[5]), .Y(_1245_) );
NAND3X1 NAND3X1_197 ( .A(_1228_), .B(_1245_), .C(_1242_), .Y(_1246_) );
AOI21X1 AOI21X1_136 ( .A(_1221_), .B(_1220_), .C(bloque_bytes[4]), .Y(_1247_) );
NAND3X1 NAND3X1_198 ( .A(bloque_bytes[5]), .B(_1241_), .C(_1240_), .Y(_1248_) );
OAI21X1 OAI21X1_190 ( .A(_1244_), .B(_1243_), .C(_1239_), .Y(_1249_) );
NAND3X1 NAND3X1_199 ( .A(_1249_), .B(_1248_), .C(_1247_), .Y(_1250_) );
NAND2X1 NAND2X1_221 ( .A(_1246_), .B(_1250_), .Y(_1251_) );
INVX2 INVX2_43 ( .A(_1251_), .Y(_1252_) );
XNOR2X1 XNOR2X1_99 ( .A(_1238_), .B(_1252_), .Y(micro_ucr_hash1_c_11__5_) );
AOI21X1 AOI21X1_137 ( .A(_1246_), .B(_1250_), .C(_1237_), .Y(_1253_) );
NAND3X1 NAND3X1_200 ( .A(_1232_), .B(_1253_), .C(_1235_), .Y(_1254_) );
NAND2X1 NAND2X1_222 ( .A(_1249_), .B(_1248_), .Y(_1255_) );
OR2X2 OR2X2_86 ( .A(_1255_), .B(_1247_), .Y(_1256_) );
INVX1 INVX1_126 ( .A(_1256_), .Y(_1257_) );
AOI21X1 AOI21X1_138 ( .A(_1247_), .B(_1255_), .C(_1226_), .Y(_1258_) );
NOR2X1 NOR2X1_125 ( .A(_1258_), .B(_1257_), .Y(_1259_) );
INVX1 INVX1_127 ( .A(bloque_bytes[6]), .Y(_1260_) );
XNOR2X1 XNOR2X1_100 ( .A(micro_ucr_hash1_b_10__6_), .B(micro_ucr_hash1_a_10__6_), .Y(_1261_) );
OR2X2 OR2X2_87 ( .A(_1261_), .B(_1260_), .Y(_1262_) );
NAND2X1 NAND2X1_223 ( .A(_1260_), .B(_1261_), .Y(_1263_) );
NAND2X1 NAND2X1_224 ( .A(_1263_), .B(_1262_), .Y(_1264_) );
OR2X2 OR2X2_88 ( .A(_1264_), .B(_1248_), .Y(_1265_) );
NAND2X1 NAND2X1_225 ( .A(_1248_), .B(_1264_), .Y(_1266_) );
NAND2X1 NAND2X1_226 ( .A(_1266_), .B(_1265_), .Y(_1267_) );
AOI21X1 AOI21X1_139 ( .A(_1259_), .B(_1254_), .C(_1267_), .Y(_1268_) );
NAND2X1 NAND2X1_227 ( .A(_1251_), .B(_1231_), .Y(_1269_) );
OAI21X1 OAI21X1_191 ( .A(_1236_), .B(_1269_), .C(_1259_), .Y(_1270_) );
INVX1 INVX1_128 ( .A(_1267_), .Y(_1271_) );
NOR2X1 NOR2X1_126 ( .A(_1271_), .B(_1270_), .Y(_1272_) );
NOR2X1 NOR2X1_127 ( .A(_1268_), .B(_1272_), .Y(micro_ucr_hash1_c_11__6_) );
INVX1 INVX1_129 ( .A(_1312_), .Y(_1273_) );
AOI21X1 AOI21X1_140 ( .A(_1232_), .B(_1273_), .C(_1323_), .Y(_1274_) );
AOI21X1 AOI21X1_141 ( .A(_1287_), .B(_1288_), .C(_1297_), .Y(_1275_) );
NAND3X1 NAND3X1_201 ( .A(_1275_), .B(_1311_), .C(_1218_), .Y(_1276_) );
AOI21X1 AOI21X1_142 ( .A(_1274_), .B(_1276_), .C(_1269_), .Y(_1277_) );
OAI21X1 OAI21X1_192 ( .A(_1252_), .B(_1226_), .C(_1256_), .Y(_1278_) );
OAI21X1 OAI21X1_193 ( .A(_1277_), .B(_1278_), .C(_1271_), .Y(_1279_) );
XOR2X1 XOR2X1_111 ( .A(micro_ucr_hash1_b_10__7_), .B(bloque_bytes[7]), .Y(_1280_) );
XNOR2X1 XNOR2X1_101 ( .A(_1280_), .B(micro_ucr_hash1_a_10__7_), .Y(_1281_) );
XNOR2X1 XNOR2X1_102 ( .A(_1281_), .B(_1262_), .Y(_1282_) );
NAND3X1 NAND3X1_202 ( .A(_1265_), .B(_1282_), .C(_1279_), .Y(_1283_) );
INVX1 INVX1_130 ( .A(_1265_), .Y(_1284_) );
INVX1 INVX1_131 ( .A(_1282_), .Y(_1285_) );
OAI21X1 OAI21X1_194 ( .A(_1268_), .B(_1284_), .C(_1285_), .Y(_1286_) );
NAND2X1 NAND2X1_228 ( .A(_1283_), .B(_1286_), .Y(micro_ucr_hash1_c_11__7_) );
XOR2X1 XOR2X1_112 ( .A(micro_ucr_hash1_b_12__4_), .B(gnd), .Y(micro_ucr_hash1_a_12__0_) );
XOR2X1 XOR2X1_113 ( .A(micro_ucr_hash1_b_12__5_), .B(gnd), .Y(micro_ucr_hash1_a_12__1_) );
XOR2X1 XOR2X1_114 ( .A(micro_ucr_hash1_b_12__6_), .B(gnd), .Y(micro_ucr_hash1_a_12__2_) );
XOR2X1 XOR2X1_115 ( .A(micro_ucr_hash1_b_12__7_), .B(gnd), .Y(micro_ucr_hash1_a_12__3_) );
XOR2X1 XOR2X1_116 ( .A(micro_ucr_hash1_c_11__4_), .B(micro_ucr_hash1_b_11__4_), .Y(micro_ucr_hash1_a_12__4_) );
XOR2X1 XOR2X1_117 ( .A(micro_ucr_hash1_c_11__5_), .B(micro_ucr_hash1_b_11__5_), .Y(micro_ucr_hash1_a_12__5_) );
XOR2X1 XOR2X1_118 ( .A(micro_ucr_hash1_c_11__6_), .B(micro_ucr_hash1_b_11__6_), .Y(micro_ucr_hash1_a_12__6_) );
XOR2X1 XOR2X1_119 ( .A(micro_ucr_hash1_c_11__7_), .B(micro_ucr_hash1_b_11__7_), .Y(micro_ucr_hash1_a_12__7_) );
INVX2 INVX2_44 ( .A(entrada_hash1_nonce_24_), .Y(_1396_) );
XNOR2X1 XNOR2X1_103 ( .A(gnd), .B(micro_ucr_hash1_a_11__0_), .Y(_1397_) );
XNOR2X1 XNOR2X1_104 ( .A(_1397_), .B(_1396_), .Y(micro_ucr_hash1_b_13__4_) );
NAND2X1 NAND2X1_229 ( .A(_1396_), .B(_1397_), .Y(_1398_) );
OR2X2 OR2X2_89 ( .A(gnd), .B(micro_ucr_hash1_a_11__1_), .Y(_1399_) );
NAND2X1 NAND2X1_230 ( .A(gnd), .B(micro_ucr_hash1_a_11__1_), .Y(_1400_) );
NAND3X1 NAND3X1_203 ( .A(entrada_hash1_nonce_25_), .B(_1400_), .C(_1399_), .Y(_1401_) );
INVX1 INVX1_132 ( .A(entrada_hash1_nonce_25_), .Y(_1402_) );
NOR2X1 NOR2X1_128 ( .A(gnd), .B(micro_ucr_hash1_a_11__1_), .Y(_1403_) );
AND2X2 AND2X2_68 ( .A(gnd), .B(micro_ucr_hash1_a_11__1_), .Y(_1404_) );
OAI21X1 OAI21X1_195 ( .A(_1404_), .B(_1403_), .C(_1402_), .Y(_1405_) );
NAND2X1 NAND2X1_231 ( .A(_1405_), .B(_1401_), .Y(_1406_) );
XNOR2X1 XNOR2X1_105 ( .A(_1406_), .B(_1398_), .Y(micro_ucr_hash1_b_13__5_) );
NAND3X1 NAND3X1_204 ( .A(_1401_), .B(_1405_), .C(_1398_), .Y(_1407_) );
NOR3X1 NOR3X1_47 ( .A(_1402_), .B(_1403_), .C(_1404_), .Y(_1408_) );
INVX1 INVX1_133 ( .A(entrada_hash1_nonce_26_), .Y(_1409_) );
NOR2X1 NOR2X1_129 ( .A(gnd), .B(micro_ucr_hash1_a_11__2_), .Y(_1410_) );
AND2X2 AND2X2_69 ( .A(gnd), .B(micro_ucr_hash1_a_11__2_), .Y(_1411_) );
NOR3X1 NOR3X1_48 ( .A(_1409_), .B(_1410_), .C(_1411_), .Y(_1412_) );
OR2X2 OR2X2_90 ( .A(gnd), .B(micro_ucr_hash1_a_11__2_), .Y(_1413_) );
NAND2X1 NAND2X1_232 ( .A(gnd), .B(micro_ucr_hash1_a_11__2_), .Y(_1414_) );
AOI21X1 AOI21X1_143 ( .A(_1414_), .B(_1413_), .C(entrada_hash1_nonce_26_), .Y(_1415_) );
OAI21X1 OAI21X1_196 ( .A(_1412_), .B(_1415_), .C(_1408_), .Y(_1416_) );
NAND3X1 NAND3X1_205 ( .A(entrada_hash1_nonce_26_), .B(_1414_), .C(_1413_), .Y(_1417_) );
OAI21X1 OAI21X1_197 ( .A(_1411_), .B(_1410_), .C(_1409_), .Y(_1418_) );
NAND3X1 NAND3X1_206 ( .A(_1418_), .B(_1401_), .C(_1417_), .Y(_1419_) );
NAND2X1 NAND2X1_233 ( .A(_1419_), .B(_1416_), .Y(_1420_) );
XNOR2X1 XNOR2X1_106 ( .A(_1420_), .B(_1407_), .Y(micro_ucr_hash1_b_13__6_) );
NAND3X1 NAND3X1_207 ( .A(_1417_), .B(_1418_), .C(_1408_), .Y(_1421_) );
OAI21X1 OAI21X1_198 ( .A(_1412_), .B(_1415_), .C(_1401_), .Y(_1422_) );
NAND2X1 NAND2X1_234 ( .A(_1421_), .B(_1422_), .Y(_1423_) );
OAI21X1 OAI21X1_199 ( .A(_1423_), .B(_1407_), .C(_1421_), .Y(_1424_) );
INVX1 INVX1_134 ( .A(entrada_hash1_nonce_27_), .Y(_1425_) );
NOR2X1 NOR2X1_130 ( .A(gnd), .B(micro_ucr_hash1_a_11__3_), .Y(_1426_) );
AND2X2 AND2X2_70 ( .A(gnd), .B(micro_ucr_hash1_a_11__3_), .Y(_1427_) );
OAI21X1 OAI21X1_200 ( .A(_1427_), .B(_1426_), .C(_1425_), .Y(_1428_) );
OR2X2 OR2X2_91 ( .A(gnd), .B(micro_ucr_hash1_a_11__3_), .Y(_1429_) );
NAND2X1 NAND2X1_235 ( .A(gnd), .B(micro_ucr_hash1_a_11__3_), .Y(_1430_) );
NAND3X1 NAND3X1_208 ( .A(entrada_hash1_nonce_27_), .B(_1430_), .C(_1429_), .Y(_1431_) );
AOI21X1 AOI21X1_144 ( .A(_1428_), .B(_1431_), .C(_1417_), .Y(_1432_) );
NAND3X1 NAND3X1_209 ( .A(_1425_), .B(_1430_), .C(_1429_), .Y(_1433_) );
OAI21X1 OAI21X1_201 ( .A(_1427_), .B(_1426_), .C(entrada_hash1_nonce_27_), .Y(_1434_) );
AOI21X1 AOI21X1_145 ( .A(_1434_), .B(_1433_), .C(_1412_), .Y(_1435_) );
NOR2X1 NOR2X1_131 ( .A(_1432_), .B(_1435_), .Y(_1327_) );
XOR2X1 XOR2X1_120 ( .A(_1424_), .B(_1327_), .Y(micro_ucr_hash1_b_13__7_) );
INVX1 INVX1_135 ( .A(entrada_hash1_nonce_28_), .Y(_1328_) );
OR2X2 OR2X2_92 ( .A(micro_ucr_hash1_b_11__4_), .B(micro_ucr_hash1_a_11__4_), .Y(_1329_) );
NAND2X1 NAND2X1_236 ( .A(micro_ucr_hash1_b_11__4_), .B(micro_ucr_hash1_a_11__4_), .Y(_1330_) );
NAND3X1 NAND3X1_210 ( .A(_1328_), .B(_1330_), .C(_1329_), .Y(_1331_) );
NOR2X1 NOR2X1_132 ( .A(micro_ucr_hash1_b_11__4_), .B(micro_ucr_hash1_a_11__4_), .Y(_1332_) );
AND2X2 AND2X2_71 ( .A(micro_ucr_hash1_b_11__4_), .B(micro_ucr_hash1_a_11__4_), .Y(_1333_) );
OAI21X1 OAI21X1_202 ( .A(_1333_), .B(_1332_), .C(entrada_hash1_nonce_28_), .Y(_1334_) );
NAND3X1 NAND3X1_211 ( .A(_1428_), .B(_1331_), .C(_1334_), .Y(_1335_) );
AOI21X1 AOI21X1_146 ( .A(_1430_), .B(_1429_), .C(entrada_hash1_nonce_27_), .Y(_1336_) );
OAI21X1 OAI21X1_203 ( .A(_1333_), .B(_1332_), .C(_1328_), .Y(_1337_) );
NAND3X1 NAND3X1_212 ( .A(entrada_hash1_nonce_28_), .B(_1330_), .C(_1329_), .Y(_1338_) );
NAND3X1 NAND3X1_213 ( .A(_1337_), .B(_1338_), .C(_1336_), .Y(_1339_) );
AND2X2 AND2X2_72 ( .A(_1339_), .B(_1335_), .Y(_1340_) );
INVX2 INVX2_45 ( .A(_1435_), .Y(_1341_) );
NOR2X1 NOR2X1_133 ( .A(_1415_), .B(_1412_), .Y(_1342_) );
AOI21X1 AOI21X1_147 ( .A(_1408_), .B(_1342_), .C(_1432_), .Y(_1343_) );
OAI21X1 OAI21X1_204 ( .A(_1423_), .B(_1407_), .C(_1343_), .Y(_1344_) );
NAND2X1 NAND2X1_237 ( .A(_1341_), .B(_1344_), .Y(_1345_) );
XNOR2X1 XNOR2X1_107 ( .A(_1345_), .B(_1340_), .Y(micro_ucr_hash1_c_12__4_) );
NAND2X1 NAND2X1_238 ( .A(_1335_), .B(_1339_), .Y(_1346_) );
OAI21X1 OAI21X1_205 ( .A(_1345_), .B(_1346_), .C(_1335_), .Y(_1347_) );
INVX1 INVX1_136 ( .A(entrada_hash1_nonce_29_), .Y(_1348_) );
OR2X2 OR2X2_93 ( .A(micro_ucr_hash1_b_11__5_), .B(micro_ucr_hash1_a_11__5_), .Y(_1349_) );
NAND2X1 NAND2X1_239 ( .A(micro_ucr_hash1_b_11__5_), .B(micro_ucr_hash1_a_11__5_), .Y(_1350_) );
NAND3X1 NAND3X1_214 ( .A(_1348_), .B(_1350_), .C(_1349_), .Y(_1351_) );
NOR2X1 NOR2X1_134 ( .A(micro_ucr_hash1_b_11__5_), .B(micro_ucr_hash1_a_11__5_), .Y(_1352_) );
AND2X2 AND2X2_73 ( .A(micro_ucr_hash1_b_11__5_), .B(micro_ucr_hash1_a_11__5_), .Y(_1353_) );
OAI21X1 OAI21X1_206 ( .A(_1353_), .B(_1352_), .C(entrada_hash1_nonce_29_), .Y(_1354_) );
NAND3X1 NAND3X1_215 ( .A(_1337_), .B(_1354_), .C(_1351_), .Y(_1355_) );
AOI21X1 AOI21X1_148 ( .A(_1330_), .B(_1329_), .C(entrada_hash1_nonce_28_), .Y(_1356_) );
NAND3X1 NAND3X1_216 ( .A(entrada_hash1_nonce_29_), .B(_1350_), .C(_1349_), .Y(_1357_) );
OAI21X1 OAI21X1_207 ( .A(_1353_), .B(_1352_), .C(_1348_), .Y(_1358_) );
NAND3X1 NAND3X1_217 ( .A(_1358_), .B(_1357_), .C(_1356_), .Y(_1359_) );
NAND2X1 NAND2X1_240 ( .A(_1355_), .B(_1359_), .Y(_1360_) );
INVX2 INVX2_46 ( .A(_1360_), .Y(_1361_) );
XNOR2X1 XNOR2X1_108 ( .A(_1347_), .B(_1361_), .Y(micro_ucr_hash1_c_12__5_) );
AOI21X1 AOI21X1_149 ( .A(_1355_), .B(_1359_), .C(_1346_), .Y(_1362_) );
NAND3X1 NAND3X1_218 ( .A(_1341_), .B(_1362_), .C(_1344_), .Y(_1363_) );
NAND2X1 NAND2X1_241 ( .A(_1358_), .B(_1357_), .Y(_1364_) );
OR2X2 OR2X2_94 ( .A(_1364_), .B(_1356_), .Y(_1365_) );
INVX1 INVX1_137 ( .A(_1365_), .Y(_1366_) );
AOI21X1 AOI21X1_150 ( .A(_1356_), .B(_1364_), .C(_1335_), .Y(_1367_) );
NOR2X1 NOR2X1_135 ( .A(_1367_), .B(_1366_), .Y(_1368_) );
INVX1 INVX1_138 ( .A(entrada_hash1_nonce_30_), .Y(_1369_) );
XNOR2X1 XNOR2X1_109 ( .A(micro_ucr_hash1_b_11__6_), .B(micro_ucr_hash1_a_11__6_), .Y(_1370_) );
OR2X2 OR2X2_95 ( .A(_1370_), .B(_1369_), .Y(_1371_) );
NAND2X1 NAND2X1_242 ( .A(_1369_), .B(_1370_), .Y(_1372_) );
NAND2X1 NAND2X1_243 ( .A(_1372_), .B(_1371_), .Y(_1373_) );
OR2X2 OR2X2_96 ( .A(_1373_), .B(_1357_), .Y(_1374_) );
NAND2X1 NAND2X1_244 ( .A(_1357_), .B(_1373_), .Y(_1375_) );
NAND2X1 NAND2X1_245 ( .A(_1375_), .B(_1374_), .Y(_1376_) );
AOI21X1 AOI21X1_151 ( .A(_1368_), .B(_1363_), .C(_1376_), .Y(_1377_) );
NAND2X1 NAND2X1_246 ( .A(_1360_), .B(_1340_), .Y(_1378_) );
OAI21X1 OAI21X1_208 ( .A(_1345_), .B(_1378_), .C(_1368_), .Y(_1379_) );
INVX1 INVX1_139 ( .A(_1376_), .Y(_1380_) );
NOR2X1 NOR2X1_136 ( .A(_1380_), .B(_1379_), .Y(_1381_) );
NOR2X1 NOR2X1_137 ( .A(_1377_), .B(_1381_), .Y(micro_ucr_hash1_c_12__6_) );
INVX1 INVX1_140 ( .A(_1421_), .Y(_1382_) );
AOI21X1 AOI21X1_152 ( .A(_1341_), .B(_1382_), .C(_1432_), .Y(_1383_) );
AOI21X1 AOI21X1_153 ( .A(_1396_), .B(_1397_), .C(_1406_), .Y(_1384_) );
NAND3X1 NAND3X1_219 ( .A(_1384_), .B(_1420_), .C(_1327_), .Y(_1385_) );
AOI21X1 AOI21X1_154 ( .A(_1383_), .B(_1385_), .C(_1378_), .Y(_1386_) );
OAI21X1 OAI21X1_209 ( .A(_1361_), .B(_1335_), .C(_1365_), .Y(_1387_) );
OAI21X1 OAI21X1_210 ( .A(_1386_), .B(_1387_), .C(_1380_), .Y(_1388_) );
XOR2X1 XOR2X1_121 ( .A(micro_ucr_hash1_b_11__7_), .B(entrada_hash1_nonce_31_), .Y(_1389_) );
XNOR2X1 XNOR2X1_110 ( .A(_1389_), .B(micro_ucr_hash1_a_11__7_), .Y(_1390_) );
XNOR2X1 XNOR2X1_111 ( .A(_1390_), .B(_1371_), .Y(_1391_) );
NAND3X1 NAND3X1_220 ( .A(_1374_), .B(_1391_), .C(_1388_), .Y(_1392_) );
INVX1 INVX1_141 ( .A(_1374_), .Y(_1393_) );
INVX1 INVX1_142 ( .A(_1391_), .Y(_1394_) );
OAI21X1 OAI21X1_211 ( .A(_1377_), .B(_1393_), .C(_1394_), .Y(_1395_) );
NAND2X1 NAND2X1_247 ( .A(_1392_), .B(_1395_), .Y(micro_ucr_hash1_c_12__7_) );
XOR2X1 XOR2X1_122 ( .A(micro_ucr_hash1_b_13__4_), .B(gnd), .Y(micro_ucr_hash1_a_13__0_) );
XOR2X1 XOR2X1_123 ( .A(micro_ucr_hash1_b_13__5_), .B(gnd), .Y(micro_ucr_hash1_a_13__1_) );
XOR2X1 XOR2X1_124 ( .A(micro_ucr_hash1_b_13__6_), .B(gnd), .Y(micro_ucr_hash1_a_13__2_) );
XOR2X1 XOR2X1_125 ( .A(micro_ucr_hash1_b_13__7_), .B(gnd), .Y(micro_ucr_hash1_a_13__3_) );
XOR2X1 XOR2X1_126 ( .A(micro_ucr_hash1_c_12__4_), .B(micro_ucr_hash1_b_12__4_), .Y(micro_ucr_hash1_a_13__4_) );
XOR2X1 XOR2X1_127 ( .A(micro_ucr_hash1_c_12__5_), .B(micro_ucr_hash1_b_12__5_), .Y(micro_ucr_hash1_a_13__5_) );
XOR2X1 XOR2X1_128 ( .A(micro_ucr_hash1_c_12__6_), .B(micro_ucr_hash1_b_12__6_), .Y(micro_ucr_hash1_a_13__6_) );
XOR2X1 XOR2X1_129 ( .A(micro_ucr_hash1_c_12__7_), .B(micro_ucr_hash1_b_12__7_), .Y(micro_ucr_hash1_a_13__7_) );
INVX2 INVX2_47 ( .A(entrada_hash1_nonce_16_), .Y(_1505_) );
XNOR2X1 XNOR2X1_112 ( .A(gnd), .B(micro_ucr_hash1_a_12__0_), .Y(_1506_) );
XNOR2X1 XNOR2X1_113 ( .A(_1506_), .B(_1505_), .Y(micro_ucr_hash1_b_14__4_) );
NAND2X1 NAND2X1_248 ( .A(_1505_), .B(_1506_), .Y(_1507_) );
OR2X2 OR2X2_97 ( .A(gnd), .B(micro_ucr_hash1_a_12__1_), .Y(_1508_) );
NAND2X1 NAND2X1_249 ( .A(gnd), .B(micro_ucr_hash1_a_12__1_), .Y(_1509_) );
NAND3X1 NAND3X1_221 ( .A(entrada_hash1_nonce_17_), .B(_1509_), .C(_1508_), .Y(_1510_) );
INVX1 INVX1_143 ( .A(entrada_hash1_nonce_17_), .Y(_1511_) );
NOR2X1 NOR2X1_138 ( .A(gnd), .B(micro_ucr_hash1_a_12__1_), .Y(_1512_) );
AND2X2 AND2X2_74 ( .A(gnd), .B(micro_ucr_hash1_a_12__1_), .Y(_1513_) );
OAI21X1 OAI21X1_212 ( .A(_1513_), .B(_1512_), .C(_1511_), .Y(_1514_) );
NAND2X1 NAND2X1_250 ( .A(_1514_), .B(_1510_), .Y(_1515_) );
XNOR2X1 XNOR2X1_114 ( .A(_1515_), .B(_1507_), .Y(micro_ucr_hash1_b_14__5_) );
NAND3X1 NAND3X1_222 ( .A(_1510_), .B(_1514_), .C(_1507_), .Y(_1516_) );
NOR3X1 NOR3X1_49 ( .A(_1511_), .B(_1512_), .C(_1513_), .Y(_1517_) );
INVX1 INVX1_144 ( .A(entrada_hash1_nonce_18_), .Y(_1518_) );
NOR2X1 NOR2X1_139 ( .A(gnd), .B(micro_ucr_hash1_a_12__2_), .Y(_1519_) );
AND2X2 AND2X2_75 ( .A(gnd), .B(micro_ucr_hash1_a_12__2_), .Y(_1520_) );
NOR3X1 NOR3X1_50 ( .A(_1518_), .B(_1519_), .C(_1520_), .Y(_1521_) );
OR2X2 OR2X2_98 ( .A(gnd), .B(micro_ucr_hash1_a_12__2_), .Y(_1522_) );
NAND2X1 NAND2X1_251 ( .A(gnd), .B(micro_ucr_hash1_a_12__2_), .Y(_1523_) );
AOI21X1 AOI21X1_155 ( .A(_1523_), .B(_1522_), .C(entrada_hash1_nonce_18_), .Y(_1524_) );
OAI21X1 OAI21X1_213 ( .A(_1521_), .B(_1524_), .C(_1517_), .Y(_1525_) );
NAND3X1 NAND3X1_223 ( .A(entrada_hash1_nonce_18_), .B(_1523_), .C(_1522_), .Y(_1526_) );
OAI21X1 OAI21X1_214 ( .A(_1520_), .B(_1519_), .C(_1518_), .Y(_1527_) );
NAND3X1 NAND3X1_224 ( .A(_1527_), .B(_1510_), .C(_1526_), .Y(_1528_) );
NAND2X1 NAND2X1_252 ( .A(_1528_), .B(_1525_), .Y(_1529_) );
XNOR2X1 XNOR2X1_115 ( .A(_1529_), .B(_1516_), .Y(micro_ucr_hash1_b_14__6_) );
NAND3X1 NAND3X1_225 ( .A(_1526_), .B(_1527_), .C(_1517_), .Y(_1530_) );
OAI21X1 OAI21X1_215 ( .A(_1521_), .B(_1524_), .C(_1510_), .Y(_1531_) );
NAND2X1 NAND2X1_253 ( .A(_1530_), .B(_1531_), .Y(_1532_) );
OAI21X1 OAI21X1_216 ( .A(_1532_), .B(_1516_), .C(_1530_), .Y(_1533_) );
INVX1 INVX1_145 ( .A(entrada_hash1_nonce_19_), .Y(_1534_) );
NOR2X1 NOR2X1_140 ( .A(gnd), .B(micro_ucr_hash1_a_12__3_), .Y(_1535_) );
AND2X2 AND2X2_76 ( .A(gnd), .B(micro_ucr_hash1_a_12__3_), .Y(_1536_) );
OAI21X1 OAI21X1_217 ( .A(_1536_), .B(_1535_), .C(_1534_), .Y(_1537_) );
OR2X2 OR2X2_99 ( .A(gnd), .B(micro_ucr_hash1_a_12__3_), .Y(_1538_) );
NAND2X1 NAND2X1_254 ( .A(gnd), .B(micro_ucr_hash1_a_12__3_), .Y(_1539_) );
NAND3X1 NAND3X1_226 ( .A(entrada_hash1_nonce_19_), .B(_1539_), .C(_1538_), .Y(_1540_) );
AOI21X1 AOI21X1_156 ( .A(_1537_), .B(_1540_), .C(_1526_), .Y(_1541_) );
NAND3X1 NAND3X1_227 ( .A(_1534_), .B(_1539_), .C(_1538_), .Y(_1542_) );
OAI21X1 OAI21X1_218 ( .A(_1536_), .B(_1535_), .C(entrada_hash1_nonce_19_), .Y(_1543_) );
AOI21X1 AOI21X1_157 ( .A(_1543_), .B(_1542_), .C(_1521_), .Y(_1544_) );
NOR2X1 NOR2X1_141 ( .A(_1541_), .B(_1544_), .Y(_1436_) );
XOR2X1 XOR2X1_130 ( .A(_1533_), .B(_1436_), .Y(micro_ucr_hash1_b_14__7_) );
INVX1 INVX1_146 ( .A(entrada_hash1_nonce_20_), .Y(_1437_) );
OR2X2 OR2X2_100 ( .A(micro_ucr_hash1_b_12__4_), .B(micro_ucr_hash1_a_12__4_), .Y(_1438_) );
NAND2X1 NAND2X1_255 ( .A(micro_ucr_hash1_b_12__4_), .B(micro_ucr_hash1_a_12__4_), .Y(_1439_) );
NAND3X1 NAND3X1_228 ( .A(_1437_), .B(_1439_), .C(_1438_), .Y(_1440_) );
NOR2X1 NOR2X1_142 ( .A(micro_ucr_hash1_b_12__4_), .B(micro_ucr_hash1_a_12__4_), .Y(_1441_) );
AND2X2 AND2X2_77 ( .A(micro_ucr_hash1_b_12__4_), .B(micro_ucr_hash1_a_12__4_), .Y(_1442_) );
OAI21X1 OAI21X1_219 ( .A(_1442_), .B(_1441_), .C(entrada_hash1_nonce_20_), .Y(_1443_) );
NAND3X1 NAND3X1_229 ( .A(_1537_), .B(_1440_), .C(_1443_), .Y(_1444_) );
AOI21X1 AOI21X1_158 ( .A(_1539_), .B(_1538_), .C(entrada_hash1_nonce_19_), .Y(_1445_) );
OAI21X1 OAI21X1_220 ( .A(_1442_), .B(_1441_), .C(_1437_), .Y(_1446_) );
NAND3X1 NAND3X1_230 ( .A(entrada_hash1_nonce_20_), .B(_1439_), .C(_1438_), .Y(_1447_) );
NAND3X1 NAND3X1_231 ( .A(_1446_), .B(_1447_), .C(_1445_), .Y(_1448_) );
AND2X2 AND2X2_78 ( .A(_1448_), .B(_1444_), .Y(_1449_) );
INVX2 INVX2_48 ( .A(_1544_), .Y(_1450_) );
NOR2X1 NOR2X1_143 ( .A(_1524_), .B(_1521_), .Y(_1451_) );
AOI21X1 AOI21X1_159 ( .A(_1517_), .B(_1451_), .C(_1541_), .Y(_1452_) );
OAI21X1 OAI21X1_221 ( .A(_1532_), .B(_1516_), .C(_1452_), .Y(_1453_) );
NAND2X1 NAND2X1_256 ( .A(_1450_), .B(_1453_), .Y(_1454_) );
XNOR2X1 XNOR2X1_116 ( .A(_1454_), .B(_1449_), .Y(micro_ucr_hash1_c_13__4_) );
NAND2X1 NAND2X1_257 ( .A(_1444_), .B(_1448_), .Y(_1455_) );
OAI21X1 OAI21X1_222 ( .A(_1454_), .B(_1455_), .C(_1444_), .Y(_1456_) );
INVX1 INVX1_147 ( .A(entrada_hash1_nonce_21_), .Y(_1457_) );
OR2X2 OR2X2_101 ( .A(micro_ucr_hash1_b_12__5_), .B(micro_ucr_hash1_a_12__5_), .Y(_1458_) );
NAND2X1 NAND2X1_258 ( .A(micro_ucr_hash1_b_12__5_), .B(micro_ucr_hash1_a_12__5_), .Y(_1459_) );
NAND3X1 NAND3X1_232 ( .A(_1457_), .B(_1459_), .C(_1458_), .Y(_1460_) );
NOR2X1 NOR2X1_144 ( .A(micro_ucr_hash1_b_12__5_), .B(micro_ucr_hash1_a_12__5_), .Y(_1461_) );
AND2X2 AND2X2_79 ( .A(micro_ucr_hash1_b_12__5_), .B(micro_ucr_hash1_a_12__5_), .Y(_1462_) );
OAI21X1 OAI21X1_223 ( .A(_1462_), .B(_1461_), .C(entrada_hash1_nonce_21_), .Y(_1463_) );
NAND3X1 NAND3X1_233 ( .A(_1446_), .B(_1463_), .C(_1460_), .Y(_1464_) );
AOI21X1 AOI21X1_160 ( .A(_1439_), .B(_1438_), .C(entrada_hash1_nonce_20_), .Y(_1465_) );
NAND3X1 NAND3X1_234 ( .A(entrada_hash1_nonce_21_), .B(_1459_), .C(_1458_), .Y(_1466_) );
OAI21X1 OAI21X1_224 ( .A(_1462_), .B(_1461_), .C(_1457_), .Y(_1467_) );
NAND3X1 NAND3X1_235 ( .A(_1467_), .B(_1466_), .C(_1465_), .Y(_1468_) );
NAND2X1 NAND2X1_259 ( .A(_1464_), .B(_1468_), .Y(_1469_) );
INVX2 INVX2_49 ( .A(_1469_), .Y(_1470_) );
XNOR2X1 XNOR2X1_117 ( .A(_1456_), .B(_1470_), .Y(micro_ucr_hash1_c_13__5_) );
AOI21X1 AOI21X1_161 ( .A(_1464_), .B(_1468_), .C(_1455_), .Y(_1471_) );
NAND3X1 NAND3X1_236 ( .A(_1450_), .B(_1471_), .C(_1453_), .Y(_1472_) );
NAND2X1 NAND2X1_260 ( .A(_1467_), .B(_1466_), .Y(_1473_) );
OR2X2 OR2X2_102 ( .A(_1473_), .B(_1465_), .Y(_1474_) );
INVX1 INVX1_148 ( .A(_1474_), .Y(_1475_) );
AOI21X1 AOI21X1_162 ( .A(_1465_), .B(_1473_), .C(_1444_), .Y(_1476_) );
NOR2X1 NOR2X1_145 ( .A(_1476_), .B(_1475_), .Y(_1477_) );
INVX1 INVX1_149 ( .A(entrada_hash1_nonce_22_), .Y(_1478_) );
XNOR2X1 XNOR2X1_118 ( .A(micro_ucr_hash1_b_12__6_), .B(micro_ucr_hash1_a_12__6_), .Y(_1479_) );
OR2X2 OR2X2_103 ( .A(_1479_), .B(_1478_), .Y(_1480_) );
NAND2X1 NAND2X1_261 ( .A(_1478_), .B(_1479_), .Y(_1481_) );
NAND2X1 NAND2X1_262 ( .A(_1481_), .B(_1480_), .Y(_1482_) );
OR2X2 OR2X2_104 ( .A(_1482_), .B(_1466_), .Y(_1483_) );
NAND2X1 NAND2X1_263 ( .A(_1466_), .B(_1482_), .Y(_1484_) );
NAND2X1 NAND2X1_264 ( .A(_1484_), .B(_1483_), .Y(_1485_) );
AOI21X1 AOI21X1_163 ( .A(_1477_), .B(_1472_), .C(_1485_), .Y(_1486_) );
NAND2X1 NAND2X1_265 ( .A(_1469_), .B(_1449_), .Y(_1487_) );
OAI21X1 OAI21X1_225 ( .A(_1454_), .B(_1487_), .C(_1477_), .Y(_1488_) );
INVX1 INVX1_150 ( .A(_1485_), .Y(_1489_) );
NOR2X1 NOR2X1_146 ( .A(_1489_), .B(_1488_), .Y(_1490_) );
NOR2X1 NOR2X1_147 ( .A(_1486_), .B(_1490_), .Y(micro_ucr_hash1_c_13__6_) );
INVX1 INVX1_151 ( .A(_1530_), .Y(_1491_) );
AOI21X1 AOI21X1_164 ( .A(_1450_), .B(_1491_), .C(_1541_), .Y(_1492_) );
AOI21X1 AOI21X1_165 ( .A(_1505_), .B(_1506_), .C(_1515_), .Y(_1493_) );
NAND3X1 NAND3X1_237 ( .A(_1493_), .B(_1529_), .C(_1436_), .Y(_1494_) );
AOI21X1 AOI21X1_166 ( .A(_1492_), .B(_1494_), .C(_1487_), .Y(_1495_) );
OAI21X1 OAI21X1_226 ( .A(_1470_), .B(_1444_), .C(_1474_), .Y(_1496_) );
OAI21X1 OAI21X1_227 ( .A(_1495_), .B(_1496_), .C(_1489_), .Y(_1497_) );
XOR2X1 XOR2X1_131 ( .A(micro_ucr_hash1_b_12__7_), .B(entrada_hash1_nonce_23_), .Y(_1498_) );
XNOR2X1 XNOR2X1_119 ( .A(_1498_), .B(micro_ucr_hash1_a_12__7_), .Y(_1499_) );
XNOR2X1 XNOR2X1_120 ( .A(_1499_), .B(_1480_), .Y(_1500_) );
NAND3X1 NAND3X1_238 ( .A(_1483_), .B(_1500_), .C(_1497_), .Y(_1501_) );
INVX1 INVX1_152 ( .A(_1483_), .Y(_1502_) );
INVX1 INVX1_153 ( .A(_1500_), .Y(_1503_) );
OAI21X1 OAI21X1_228 ( .A(_1486_), .B(_1502_), .C(_1503_), .Y(_1504_) );
NAND2X1 NAND2X1_266 ( .A(_1501_), .B(_1504_), .Y(micro_ucr_hash1_c_13__7_) );
XOR2X1 XOR2X1_132 ( .A(micro_ucr_hash1_b_14__4_), .B(gnd), .Y(micro_ucr_hash1_a_14__0_) );
XOR2X1 XOR2X1_133 ( .A(micro_ucr_hash1_b_14__5_), .B(gnd), .Y(micro_ucr_hash1_a_14__1_) );
XOR2X1 XOR2X1_134 ( .A(micro_ucr_hash1_b_14__6_), .B(gnd), .Y(micro_ucr_hash1_a_14__2_) );
XOR2X1 XOR2X1_135 ( .A(micro_ucr_hash1_b_14__7_), .B(gnd), .Y(micro_ucr_hash1_a_14__3_) );
XOR2X1 XOR2X1_136 ( .A(micro_ucr_hash1_c_13__4_), .B(micro_ucr_hash1_b_13__4_), .Y(micro_ucr_hash1_a_14__4_) );
XOR2X1 XOR2X1_137 ( .A(micro_ucr_hash1_c_13__5_), .B(micro_ucr_hash1_b_13__5_), .Y(micro_ucr_hash1_a_14__5_) );
XOR2X1 XOR2X1_138 ( .A(micro_ucr_hash1_c_13__6_), .B(micro_ucr_hash1_b_13__6_), .Y(micro_ucr_hash1_a_14__6_) );
XOR2X1 XOR2X1_139 ( .A(micro_ucr_hash1_c_13__7_), .B(micro_ucr_hash1_b_13__7_), .Y(micro_ucr_hash1_a_14__7_) );
INVX2 INVX2_50 ( .A(entrada_hash1_nonce_8_), .Y(_1614_) );
XNOR2X1 XNOR2X1_121 ( .A(gnd), .B(micro_ucr_hash1_a_13__0_), .Y(_1615_) );
XNOR2X1 XNOR2X1_122 ( .A(_1615_), .B(_1614_), .Y(micro_ucr_hash1_b_15__4_) );
NAND2X1 NAND2X1_267 ( .A(_1614_), .B(_1615_), .Y(_1616_) );
OR2X2 OR2X2_105 ( .A(gnd), .B(micro_ucr_hash1_a_13__1_), .Y(_1617_) );
NAND2X1 NAND2X1_268 ( .A(gnd), .B(micro_ucr_hash1_a_13__1_), .Y(_1618_) );
NAND3X1 NAND3X1_239 ( .A(entrada_hash1_nonce_9_), .B(_1618_), .C(_1617_), .Y(_1619_) );
INVX1 INVX1_154 ( .A(entrada_hash1_nonce_9_), .Y(_1620_) );
NOR2X1 NOR2X1_148 ( .A(gnd), .B(micro_ucr_hash1_a_13__1_), .Y(_1621_) );
AND2X2 AND2X2_80 ( .A(gnd), .B(micro_ucr_hash1_a_13__1_), .Y(_1622_) );
OAI21X1 OAI21X1_229 ( .A(_1622_), .B(_1621_), .C(_1620_), .Y(_1623_) );
NAND2X1 NAND2X1_269 ( .A(_1623_), .B(_1619_), .Y(_1624_) );
XNOR2X1 XNOR2X1_123 ( .A(_1624_), .B(_1616_), .Y(micro_ucr_hash1_b_15__5_) );
NAND3X1 NAND3X1_240 ( .A(_1619_), .B(_1623_), .C(_1616_), .Y(_1625_) );
NOR3X1 NOR3X1_51 ( .A(_1620_), .B(_1621_), .C(_1622_), .Y(_1626_) );
INVX1 INVX1_155 ( .A(entrada_hash1_nonce_10_), .Y(_1627_) );
NOR2X1 NOR2X1_149 ( .A(gnd), .B(micro_ucr_hash1_a_13__2_), .Y(_1628_) );
AND2X2 AND2X2_81 ( .A(gnd), .B(micro_ucr_hash1_a_13__2_), .Y(_1629_) );
NOR3X1 NOR3X1_52 ( .A(_1627_), .B(_1628_), .C(_1629_), .Y(_1630_) );
OR2X2 OR2X2_106 ( .A(gnd), .B(micro_ucr_hash1_a_13__2_), .Y(_1631_) );
NAND2X1 NAND2X1_270 ( .A(gnd), .B(micro_ucr_hash1_a_13__2_), .Y(_1632_) );
AOI21X1 AOI21X1_167 ( .A(_1632_), .B(_1631_), .C(entrada_hash1_nonce_10_), .Y(_1633_) );
OAI21X1 OAI21X1_230 ( .A(_1630_), .B(_1633_), .C(_1626_), .Y(_1634_) );
NAND3X1 NAND3X1_241 ( .A(entrada_hash1_nonce_10_), .B(_1632_), .C(_1631_), .Y(_1635_) );
OAI21X1 OAI21X1_231 ( .A(_1629_), .B(_1628_), .C(_1627_), .Y(_1636_) );
NAND3X1 NAND3X1_242 ( .A(_1636_), .B(_1619_), .C(_1635_), .Y(_1637_) );
NAND2X1 NAND2X1_271 ( .A(_1637_), .B(_1634_), .Y(_1638_) );
XNOR2X1 XNOR2X1_124 ( .A(_1638_), .B(_1625_), .Y(micro_ucr_hash1_b_15__6_) );
NAND3X1 NAND3X1_243 ( .A(_1635_), .B(_1636_), .C(_1626_), .Y(_1639_) );
OAI21X1 OAI21X1_232 ( .A(_1630_), .B(_1633_), .C(_1619_), .Y(_1640_) );
NAND2X1 NAND2X1_272 ( .A(_1639_), .B(_1640_), .Y(_1641_) );
OAI21X1 OAI21X1_233 ( .A(_1641_), .B(_1625_), .C(_1639_), .Y(_1642_) );
INVX1 INVX1_156 ( .A(entrada_hash1_nonce_11_), .Y(_1643_) );
NOR2X1 NOR2X1_150 ( .A(gnd), .B(micro_ucr_hash1_a_13__3_), .Y(_1644_) );
AND2X2 AND2X2_82 ( .A(gnd), .B(micro_ucr_hash1_a_13__3_), .Y(_1645_) );
OAI21X1 OAI21X1_234 ( .A(_1645_), .B(_1644_), .C(_1643_), .Y(_1646_) );
OR2X2 OR2X2_107 ( .A(gnd), .B(micro_ucr_hash1_a_13__3_), .Y(_1647_) );
NAND2X1 NAND2X1_273 ( .A(gnd), .B(micro_ucr_hash1_a_13__3_), .Y(_1648_) );
NAND3X1 NAND3X1_244 ( .A(entrada_hash1_nonce_11_), .B(_1648_), .C(_1647_), .Y(_1649_) );
AOI21X1 AOI21X1_168 ( .A(_1646_), .B(_1649_), .C(_1635_), .Y(_1650_) );
NAND3X1 NAND3X1_245 ( .A(_1643_), .B(_1648_), .C(_1647_), .Y(_1651_) );
OAI21X1 OAI21X1_235 ( .A(_1645_), .B(_1644_), .C(entrada_hash1_nonce_11_), .Y(_1652_) );
AOI21X1 AOI21X1_169 ( .A(_1652_), .B(_1651_), .C(_1630_), .Y(_1653_) );
NOR2X1 NOR2X1_151 ( .A(_1650_), .B(_1653_), .Y(_1545_) );
XOR2X1 XOR2X1_140 ( .A(_1642_), .B(_1545_), .Y(micro_ucr_hash1_b_15__7_) );
INVX1 INVX1_157 ( .A(entrada_hash1_nonce_12_), .Y(_1546_) );
OR2X2 OR2X2_108 ( .A(micro_ucr_hash1_b_13__4_), .B(micro_ucr_hash1_a_13__4_), .Y(_1547_) );
NAND2X1 NAND2X1_274 ( .A(micro_ucr_hash1_b_13__4_), .B(micro_ucr_hash1_a_13__4_), .Y(_1548_) );
NAND3X1 NAND3X1_246 ( .A(_1546_), .B(_1548_), .C(_1547_), .Y(_1549_) );
NOR2X1 NOR2X1_152 ( .A(micro_ucr_hash1_b_13__4_), .B(micro_ucr_hash1_a_13__4_), .Y(_1550_) );
AND2X2 AND2X2_83 ( .A(micro_ucr_hash1_b_13__4_), .B(micro_ucr_hash1_a_13__4_), .Y(_1551_) );
OAI21X1 OAI21X1_236 ( .A(_1551_), .B(_1550_), .C(entrada_hash1_nonce_12_), .Y(_1552_) );
NAND3X1 NAND3X1_247 ( .A(_1646_), .B(_1549_), .C(_1552_), .Y(_1553_) );
AOI21X1 AOI21X1_170 ( .A(_1648_), .B(_1647_), .C(entrada_hash1_nonce_11_), .Y(_1554_) );
OAI21X1 OAI21X1_237 ( .A(_1551_), .B(_1550_), .C(_1546_), .Y(_1555_) );
NAND3X1 NAND3X1_248 ( .A(entrada_hash1_nonce_12_), .B(_1548_), .C(_1547_), .Y(_1556_) );
NAND3X1 NAND3X1_249 ( .A(_1555_), .B(_1556_), .C(_1554_), .Y(_1557_) );
AND2X2 AND2X2_84 ( .A(_1557_), .B(_1553_), .Y(_1558_) );
INVX2 INVX2_51 ( .A(_1653_), .Y(_1559_) );
NOR2X1 NOR2X1_153 ( .A(_1633_), .B(_1630_), .Y(_1560_) );
AOI21X1 AOI21X1_171 ( .A(_1626_), .B(_1560_), .C(_1650_), .Y(_1561_) );
OAI21X1 OAI21X1_238 ( .A(_1641_), .B(_1625_), .C(_1561_), .Y(_1562_) );
NAND2X1 NAND2X1_275 ( .A(_1559_), .B(_1562_), .Y(_1563_) );
XNOR2X1 XNOR2X1_125 ( .A(_1563_), .B(_1558_), .Y(micro_ucr_hash1_c_14__4_) );
NAND2X1 NAND2X1_276 ( .A(_1553_), .B(_1557_), .Y(_1564_) );
OAI21X1 OAI21X1_239 ( .A(_1563_), .B(_1564_), .C(_1553_), .Y(_1565_) );
INVX1 INVX1_158 ( .A(entrada_hash1_nonce_13_), .Y(_1566_) );
OR2X2 OR2X2_109 ( .A(micro_ucr_hash1_b_13__5_), .B(micro_ucr_hash1_a_13__5_), .Y(_1567_) );
NAND2X1 NAND2X1_277 ( .A(micro_ucr_hash1_b_13__5_), .B(micro_ucr_hash1_a_13__5_), .Y(_1568_) );
NAND3X1 NAND3X1_250 ( .A(_1566_), .B(_1568_), .C(_1567_), .Y(_1569_) );
NOR2X1 NOR2X1_154 ( .A(micro_ucr_hash1_b_13__5_), .B(micro_ucr_hash1_a_13__5_), .Y(_1570_) );
AND2X2 AND2X2_85 ( .A(micro_ucr_hash1_b_13__5_), .B(micro_ucr_hash1_a_13__5_), .Y(_1571_) );
OAI21X1 OAI21X1_240 ( .A(_1571_), .B(_1570_), .C(entrada_hash1_nonce_13_), .Y(_1572_) );
NAND3X1 NAND3X1_251 ( .A(_1555_), .B(_1572_), .C(_1569_), .Y(_1573_) );
AOI21X1 AOI21X1_172 ( .A(_1548_), .B(_1547_), .C(entrada_hash1_nonce_12_), .Y(_1574_) );
NAND3X1 NAND3X1_252 ( .A(entrada_hash1_nonce_13_), .B(_1568_), .C(_1567_), .Y(_1575_) );
OAI21X1 OAI21X1_241 ( .A(_1571_), .B(_1570_), .C(_1566_), .Y(_1576_) );
NAND3X1 NAND3X1_253 ( .A(_1576_), .B(_1575_), .C(_1574_), .Y(_1577_) );
NAND2X1 NAND2X1_278 ( .A(_1573_), .B(_1577_), .Y(_1578_) );
INVX2 INVX2_52 ( .A(_1578_), .Y(_1579_) );
XNOR2X1 XNOR2X1_126 ( .A(_1565_), .B(_1579_), .Y(micro_ucr_hash1_c_14__5_) );
AOI21X1 AOI21X1_173 ( .A(_1573_), .B(_1577_), .C(_1564_), .Y(_1580_) );
NAND3X1 NAND3X1_254 ( .A(_1559_), .B(_1580_), .C(_1562_), .Y(_1581_) );
NAND2X1 NAND2X1_279 ( .A(_1576_), .B(_1575_), .Y(_1582_) );
OR2X2 OR2X2_110 ( .A(_1582_), .B(_1574_), .Y(_1583_) );
INVX1 INVX1_159 ( .A(_1583_), .Y(_1584_) );
AOI21X1 AOI21X1_174 ( .A(_1574_), .B(_1582_), .C(_1553_), .Y(_1585_) );
NOR2X1 NOR2X1_155 ( .A(_1585_), .B(_1584_), .Y(_1586_) );
INVX1 INVX1_160 ( .A(entrada_hash1_nonce_14_), .Y(_1587_) );
XNOR2X1 XNOR2X1_127 ( .A(micro_ucr_hash1_b_13__6_), .B(micro_ucr_hash1_a_13__6_), .Y(_1588_) );
OR2X2 OR2X2_111 ( .A(_1588_), .B(_1587_), .Y(_1589_) );
NAND2X1 NAND2X1_280 ( .A(_1587_), .B(_1588_), .Y(_1590_) );
NAND2X1 NAND2X1_281 ( .A(_1590_), .B(_1589_), .Y(_1591_) );
OR2X2 OR2X2_112 ( .A(_1591_), .B(_1575_), .Y(_1592_) );
NAND2X1 NAND2X1_282 ( .A(_1575_), .B(_1591_), .Y(_1593_) );
NAND2X1 NAND2X1_283 ( .A(_1593_), .B(_1592_), .Y(_1594_) );
AOI21X1 AOI21X1_175 ( .A(_1586_), .B(_1581_), .C(_1594_), .Y(_1595_) );
NAND2X1 NAND2X1_284 ( .A(_1578_), .B(_1558_), .Y(_1596_) );
OAI21X1 OAI21X1_242 ( .A(_1563_), .B(_1596_), .C(_1586_), .Y(_1597_) );
INVX1 INVX1_161 ( .A(_1594_), .Y(_1598_) );
NOR2X1 NOR2X1_156 ( .A(_1598_), .B(_1597_), .Y(_1599_) );
NOR2X1 NOR2X1_157 ( .A(_1595_), .B(_1599_), .Y(micro_ucr_hash1_c_14__6_) );
INVX1 INVX1_162 ( .A(_1639_), .Y(_1600_) );
AOI21X1 AOI21X1_176 ( .A(_1559_), .B(_1600_), .C(_1650_), .Y(_1601_) );
AOI21X1 AOI21X1_177 ( .A(_1614_), .B(_1615_), .C(_1624_), .Y(_1602_) );
NAND3X1 NAND3X1_255 ( .A(_1602_), .B(_1638_), .C(_1545_), .Y(_1603_) );
AOI21X1 AOI21X1_178 ( .A(_1601_), .B(_1603_), .C(_1596_), .Y(_1604_) );
OAI21X1 OAI21X1_243 ( .A(_1579_), .B(_1553_), .C(_1583_), .Y(_1605_) );
OAI21X1 OAI21X1_244 ( .A(_1604_), .B(_1605_), .C(_1598_), .Y(_1606_) );
XOR2X1 XOR2X1_141 ( .A(micro_ucr_hash1_b_13__7_), .B(entrada_hash1_nonce_15_), .Y(_1607_) );
XNOR2X1 XNOR2X1_128 ( .A(_1607_), .B(micro_ucr_hash1_a_13__7_), .Y(_1608_) );
XNOR2X1 XNOR2X1_129 ( .A(_1608_), .B(_1589_), .Y(_1609_) );
NAND3X1 NAND3X1_256 ( .A(_1592_), .B(_1609_), .C(_1606_), .Y(_1610_) );
INVX1 INVX1_163 ( .A(_1592_), .Y(_1611_) );
INVX1 INVX1_164 ( .A(_1609_), .Y(_1612_) );
OAI21X1 OAI21X1_245 ( .A(_1595_), .B(_1611_), .C(_1612_), .Y(_1613_) );
NAND2X1 NAND2X1_285 ( .A(_1610_), .B(_1613_), .Y(micro_ucr_hash1_c_14__7_) );
XOR2X1 XOR2X1_142 ( .A(micro_ucr_hash1_b_15__4_), .B(gnd), .Y(micro_ucr_hash1_a_15__0_) );
XOR2X1 XOR2X1_143 ( .A(micro_ucr_hash1_b_15__5_), .B(gnd), .Y(micro_ucr_hash1_a_15__1_) );
XOR2X1 XOR2X1_144 ( .A(micro_ucr_hash1_b_15__6_), .B(gnd), .Y(micro_ucr_hash1_a_15__2_) );
XOR2X1 XOR2X1_145 ( .A(micro_ucr_hash1_b_15__7_), .B(gnd), .Y(micro_ucr_hash1_a_15__3_) );
XOR2X1 XOR2X1_146 ( .A(micro_ucr_hash1_c_14__4_), .B(micro_ucr_hash1_b_14__4_), .Y(micro_ucr_hash1_a_15__4_) );
XOR2X1 XOR2X1_147 ( .A(micro_ucr_hash1_c_14__5_), .B(micro_ucr_hash1_b_14__5_), .Y(micro_ucr_hash1_a_15__5_) );
XOR2X1 XOR2X1_148 ( .A(micro_ucr_hash1_c_14__6_), .B(micro_ucr_hash1_b_14__6_), .Y(micro_ucr_hash1_a_15__6_) );
XOR2X1 XOR2X1_149 ( .A(micro_ucr_hash1_c_14__7_), .B(micro_ucr_hash1_b_14__7_), .Y(micro_ucr_hash1_a_15__7_) );
INVX2 INVX2_53 ( .A(entrada_hash1_nonce_0_), .Y(_1723_) );
XNOR2X1 XNOR2X1_130 ( .A(gnd), .B(micro_ucr_hash1_a_14__0_), .Y(_1724_) );
XNOR2X1 XNOR2X1_131 ( .A(_1724_), .B(_1723_), .Y(micro_ucr_hash1_b_16__4_) );
NAND2X1 NAND2X1_286 ( .A(_1723_), .B(_1724_), .Y(_1725_) );
OR2X2 OR2X2_113 ( .A(gnd), .B(micro_ucr_hash1_a_14__1_), .Y(_1726_) );
NAND2X1 NAND2X1_287 ( .A(gnd), .B(micro_ucr_hash1_a_14__1_), .Y(_1727_) );
NAND3X1 NAND3X1_257 ( .A(entrada_hash1_nonce_1_), .B(_1727_), .C(_1726_), .Y(_1728_) );
INVX1 INVX1_165 ( .A(entrada_hash1_nonce_1_), .Y(_1729_) );
NOR2X1 NOR2X1_158 ( .A(gnd), .B(micro_ucr_hash1_a_14__1_), .Y(_1730_) );
AND2X2 AND2X2_86 ( .A(gnd), .B(micro_ucr_hash1_a_14__1_), .Y(_1731_) );
OAI21X1 OAI21X1_246 ( .A(_1731_), .B(_1730_), .C(_1729_), .Y(_1732_) );
NAND2X1 NAND2X1_288 ( .A(_1732_), .B(_1728_), .Y(_1733_) );
XNOR2X1 XNOR2X1_132 ( .A(_1733_), .B(_1725_), .Y(micro_ucr_hash1_b_16__5_) );
NAND3X1 NAND3X1_258 ( .A(_1728_), .B(_1732_), .C(_1725_), .Y(_1734_) );
NOR3X1 NOR3X1_53 ( .A(_1729_), .B(_1730_), .C(_1731_), .Y(_1735_) );
INVX1 INVX1_166 ( .A(entrada_hash1_nonce_2_), .Y(_1736_) );
NOR2X1 NOR2X1_159 ( .A(gnd), .B(micro_ucr_hash1_a_14__2_), .Y(_1737_) );
AND2X2 AND2X2_87 ( .A(gnd), .B(micro_ucr_hash1_a_14__2_), .Y(_1738_) );
NOR3X1 NOR3X1_54 ( .A(_1736_), .B(_1737_), .C(_1738_), .Y(_1739_) );
OR2X2 OR2X2_114 ( .A(gnd), .B(micro_ucr_hash1_a_14__2_), .Y(_1740_) );
NAND2X1 NAND2X1_289 ( .A(gnd), .B(micro_ucr_hash1_a_14__2_), .Y(_1741_) );
AOI21X1 AOI21X1_179 ( .A(_1741_), .B(_1740_), .C(entrada_hash1_nonce_2_), .Y(_1742_) );
OAI21X1 OAI21X1_247 ( .A(_1739_), .B(_1742_), .C(_1735_), .Y(_1743_) );
NAND3X1 NAND3X1_259 ( .A(entrada_hash1_nonce_2_), .B(_1741_), .C(_1740_), .Y(_1744_) );
OAI21X1 OAI21X1_248 ( .A(_1738_), .B(_1737_), .C(_1736_), .Y(_1745_) );
NAND3X1 NAND3X1_260 ( .A(_1745_), .B(_1728_), .C(_1744_), .Y(_1746_) );
NAND2X1 NAND2X1_290 ( .A(_1746_), .B(_1743_), .Y(_1747_) );
XNOR2X1 XNOR2X1_133 ( .A(_1747_), .B(_1734_), .Y(micro_ucr_hash1_b_16__6_) );
NAND3X1 NAND3X1_261 ( .A(_1744_), .B(_1745_), .C(_1735_), .Y(_1748_) );
OAI21X1 OAI21X1_249 ( .A(_1739_), .B(_1742_), .C(_1728_), .Y(_1749_) );
NAND2X1 NAND2X1_291 ( .A(_1748_), .B(_1749_), .Y(_1750_) );
OAI21X1 OAI21X1_250 ( .A(_1750_), .B(_1734_), .C(_1748_), .Y(_1751_) );
INVX1 INVX1_167 ( .A(entrada_hash1_nonce_3_), .Y(_1752_) );
NOR2X1 NOR2X1_160 ( .A(gnd), .B(micro_ucr_hash1_a_14__3_), .Y(_1753_) );
AND2X2 AND2X2_88 ( .A(gnd), .B(micro_ucr_hash1_a_14__3_), .Y(_1754_) );
OAI21X1 OAI21X1_251 ( .A(_1754_), .B(_1753_), .C(_1752_), .Y(_1755_) );
OR2X2 OR2X2_115 ( .A(gnd), .B(micro_ucr_hash1_a_14__3_), .Y(_1756_) );
NAND2X1 NAND2X1_292 ( .A(gnd), .B(micro_ucr_hash1_a_14__3_), .Y(_1757_) );
NAND3X1 NAND3X1_262 ( .A(entrada_hash1_nonce_3_), .B(_1757_), .C(_1756_), .Y(_1758_) );
AOI21X1 AOI21X1_180 ( .A(_1755_), .B(_1758_), .C(_1744_), .Y(_1759_) );
NAND3X1 NAND3X1_263 ( .A(_1752_), .B(_1757_), .C(_1756_), .Y(_1760_) );
OAI21X1 OAI21X1_252 ( .A(_1754_), .B(_1753_), .C(entrada_hash1_nonce_3_), .Y(_1761_) );
AOI21X1 AOI21X1_181 ( .A(_1761_), .B(_1760_), .C(_1739_), .Y(_1762_) );
NOR2X1 NOR2X1_161 ( .A(_1759_), .B(_1762_), .Y(_1654_) );
XOR2X1 XOR2X1_150 ( .A(_1751_), .B(_1654_), .Y(micro_ucr_hash1_b_16__7_) );
INVX1 INVX1_168 ( .A(entrada_hash1_nonce_4_), .Y(_1655_) );
OR2X2 OR2X2_116 ( .A(micro_ucr_hash1_b_14__4_), .B(micro_ucr_hash1_a_14__4_), .Y(_1656_) );
NAND2X1 NAND2X1_293 ( .A(micro_ucr_hash1_b_14__4_), .B(micro_ucr_hash1_a_14__4_), .Y(_1657_) );
NAND3X1 NAND3X1_264 ( .A(_1655_), .B(_1657_), .C(_1656_), .Y(_1658_) );
NOR2X1 NOR2X1_162 ( .A(micro_ucr_hash1_b_14__4_), .B(micro_ucr_hash1_a_14__4_), .Y(_1659_) );
AND2X2 AND2X2_89 ( .A(micro_ucr_hash1_b_14__4_), .B(micro_ucr_hash1_a_14__4_), .Y(_1660_) );
OAI21X1 OAI21X1_253 ( .A(_1660_), .B(_1659_), .C(entrada_hash1_nonce_4_), .Y(_1661_) );
NAND3X1 NAND3X1_265 ( .A(_1755_), .B(_1658_), .C(_1661_), .Y(_1662_) );
AOI21X1 AOI21X1_182 ( .A(_1757_), .B(_1756_), .C(entrada_hash1_nonce_3_), .Y(_1663_) );
OAI21X1 OAI21X1_254 ( .A(_1660_), .B(_1659_), .C(_1655_), .Y(_1664_) );
NAND3X1 NAND3X1_266 ( .A(entrada_hash1_nonce_4_), .B(_1657_), .C(_1656_), .Y(_1665_) );
NAND3X1 NAND3X1_267 ( .A(_1664_), .B(_1665_), .C(_1663_), .Y(_1666_) );
AND2X2 AND2X2_90 ( .A(_1666_), .B(_1662_), .Y(_1667_) );
INVX2 INVX2_54 ( .A(_1762_), .Y(_1668_) );
NOR2X1 NOR2X1_163 ( .A(_1742_), .B(_1739_), .Y(_1669_) );
AOI21X1 AOI21X1_183 ( .A(_1735_), .B(_1669_), .C(_1759_), .Y(_1670_) );
OAI21X1 OAI21X1_255 ( .A(_1750_), .B(_1734_), .C(_1670_), .Y(_1671_) );
NAND2X1 NAND2X1_294 ( .A(_1668_), .B(_1671_), .Y(_1672_) );
XNOR2X1 XNOR2X1_134 ( .A(_1672_), .B(_1667_), .Y(micro_ucr_hash1_c_15__4_) );
NAND2X1 NAND2X1_295 ( .A(_1662_), .B(_1666_), .Y(_1673_) );
OAI21X1 OAI21X1_256 ( .A(_1672_), .B(_1673_), .C(_1662_), .Y(_1674_) );
INVX1 INVX1_169 ( .A(entrada_hash1_nonce_5_), .Y(_1675_) );
OR2X2 OR2X2_117 ( .A(micro_ucr_hash1_b_14__5_), .B(micro_ucr_hash1_a_14__5_), .Y(_1676_) );
NAND2X1 NAND2X1_296 ( .A(micro_ucr_hash1_b_14__5_), .B(micro_ucr_hash1_a_14__5_), .Y(_1677_) );
NAND3X1 NAND3X1_268 ( .A(_1675_), .B(_1677_), .C(_1676_), .Y(_1678_) );
NOR2X1 NOR2X1_164 ( .A(micro_ucr_hash1_b_14__5_), .B(micro_ucr_hash1_a_14__5_), .Y(_1679_) );
AND2X2 AND2X2_91 ( .A(micro_ucr_hash1_b_14__5_), .B(micro_ucr_hash1_a_14__5_), .Y(_1680_) );
OAI21X1 OAI21X1_257 ( .A(_1680_), .B(_1679_), .C(entrada_hash1_nonce_5_), .Y(_1681_) );
NAND3X1 NAND3X1_269 ( .A(_1664_), .B(_1681_), .C(_1678_), .Y(_1682_) );
AOI21X1 AOI21X1_184 ( .A(_1657_), .B(_1656_), .C(entrada_hash1_nonce_4_), .Y(_1683_) );
NAND3X1 NAND3X1_270 ( .A(entrada_hash1_nonce_5_), .B(_1677_), .C(_1676_), .Y(_1684_) );
OAI21X1 OAI21X1_258 ( .A(_1680_), .B(_1679_), .C(_1675_), .Y(_1685_) );
NAND3X1 NAND3X1_271 ( .A(_1685_), .B(_1684_), .C(_1683_), .Y(_1686_) );
NAND2X1 NAND2X1_297 ( .A(_1682_), .B(_1686_), .Y(_1687_) );
INVX2 INVX2_55 ( .A(_1687_), .Y(_1688_) );
XNOR2X1 XNOR2X1_135 ( .A(_1674_), .B(_1688_), .Y(micro_ucr_hash1_c_15__5_) );
AOI21X1 AOI21X1_185 ( .A(_1682_), .B(_1686_), .C(_1673_), .Y(_1689_) );
NAND3X1 NAND3X1_272 ( .A(_1668_), .B(_1689_), .C(_1671_), .Y(_1690_) );
NAND2X1 NAND2X1_298 ( .A(_1685_), .B(_1684_), .Y(_1691_) );
OR2X2 OR2X2_118 ( .A(_1691_), .B(_1683_), .Y(_1692_) );
INVX1 INVX1_170 ( .A(_1692_), .Y(_1693_) );
AOI21X1 AOI21X1_186 ( .A(_1683_), .B(_1691_), .C(_1662_), .Y(_1694_) );
NOR2X1 NOR2X1_165 ( .A(_1694_), .B(_1693_), .Y(_1695_) );
INVX1 INVX1_171 ( .A(entrada_hash1_nonce_6_), .Y(_1696_) );
XNOR2X1 XNOR2X1_136 ( .A(micro_ucr_hash1_b_14__6_), .B(micro_ucr_hash1_a_14__6_), .Y(_1697_) );
OR2X2 OR2X2_119 ( .A(_1697_), .B(_1696_), .Y(_1698_) );
NAND2X1 NAND2X1_299 ( .A(_1696_), .B(_1697_), .Y(_1699_) );
NAND2X1 NAND2X1_300 ( .A(_1699_), .B(_1698_), .Y(_1700_) );
OR2X2 OR2X2_120 ( .A(_1700_), .B(_1684_), .Y(_1701_) );
NAND2X1 NAND2X1_301 ( .A(_1684_), .B(_1700_), .Y(_1702_) );
NAND2X1 NAND2X1_302 ( .A(_1702_), .B(_1701_), .Y(_1703_) );
AOI21X1 AOI21X1_187 ( .A(_1695_), .B(_1690_), .C(_1703_), .Y(_1704_) );
NAND2X1 NAND2X1_303 ( .A(_1687_), .B(_1667_), .Y(_1705_) );
OAI21X1 OAI21X1_259 ( .A(_1672_), .B(_1705_), .C(_1695_), .Y(_1706_) );
INVX1 INVX1_172 ( .A(_1703_), .Y(_1707_) );
NOR2X1 NOR2X1_166 ( .A(_1707_), .B(_1706_), .Y(_1708_) );
NOR2X1 NOR2X1_167 ( .A(_1704_), .B(_1708_), .Y(micro_ucr_hash1_c_15__6_) );
INVX1 INVX1_173 ( .A(_1748_), .Y(_1709_) );
AOI21X1 AOI21X1_188 ( .A(_1668_), .B(_1709_), .C(_1759_), .Y(_1710_) );
AOI21X1 AOI21X1_189 ( .A(_1723_), .B(_1724_), .C(_1733_), .Y(_1711_) );
NAND3X1 NAND3X1_273 ( .A(_1711_), .B(_1747_), .C(_1654_), .Y(_1712_) );
AOI21X1 AOI21X1_190 ( .A(_1710_), .B(_1712_), .C(_1705_), .Y(_1713_) );
OAI21X1 OAI21X1_260 ( .A(_1688_), .B(_1662_), .C(_1692_), .Y(_1714_) );
OAI21X1 OAI21X1_261 ( .A(_1713_), .B(_1714_), .C(_1707_), .Y(_1715_) );
XOR2X1 XOR2X1_151 ( .A(micro_ucr_hash1_b_14__7_), .B(entrada_hash1_nonce_7_), .Y(_1716_) );
XNOR2X1 XNOR2X1_137 ( .A(_1716_), .B(micro_ucr_hash1_a_14__7_), .Y(_1717_) );
XNOR2X1 XNOR2X1_138 ( .A(_1717_), .B(_1698_), .Y(_1718_) );
NAND3X1 NAND3X1_274 ( .A(_1701_), .B(_1718_), .C(_1715_), .Y(_1719_) );
INVX1 INVX1_174 ( .A(_1701_), .Y(_1720_) );
INVX1 INVX1_175 ( .A(_1718_), .Y(_1721_) );
OAI21X1 OAI21X1_262 ( .A(_1704_), .B(_1720_), .C(_1721_), .Y(_1722_) );
NAND2X1 NAND2X1_304 ( .A(_1719_), .B(_1722_), .Y(micro_ucr_hash1_c_15__7_) );
XOR2X1 XOR2X1_152 ( .A(micro_ucr_hash1_b_16__4_), .B(gnd), .Y(micro_ucr_hash1_a_16__0_) );
XOR2X1 XOR2X1_153 ( .A(micro_ucr_hash1_b_16__5_), .B(gnd), .Y(micro_ucr_hash1_a_16__1_) );
XOR2X1 XOR2X1_154 ( .A(micro_ucr_hash1_b_16__6_), .B(gnd), .Y(micro_ucr_hash1_a_16__2_) );
XOR2X1 XOR2X1_155 ( .A(micro_ucr_hash1_b_16__7_), .B(gnd), .Y(micro_ucr_hash1_a_16__3_) );
XOR2X1 XOR2X1_156 ( .A(micro_ucr_hash1_c_15__4_), .B(micro_ucr_hash1_b_15__4_), .Y(micro_ucr_hash1_a_16__4_) );
XOR2X1 XOR2X1_157 ( .A(micro_ucr_hash1_c_15__5_), .B(micro_ucr_hash1_b_15__5_), .Y(micro_ucr_hash1_a_16__5_) );
XOR2X1 XOR2X1_158 ( .A(micro_ucr_hash1_c_15__6_), .B(micro_ucr_hash1_b_15__6_), .Y(micro_ucr_hash1_a_16__6_) );
XOR2X1 XOR2X1_159 ( .A(micro_ucr_hash1_c_15__7_), .B(micro_ucr_hash1_b_15__7_), .Y(micro_ucr_hash1_a_16__7_) );
INVX2 INVX2_56 ( .A(micro_ucr_hash1_W_16__0_), .Y(_1832_) );
XNOR2X1 XNOR2X1_139 ( .A(gnd), .B(micro_ucr_hash1_a_15__0_), .Y(_1833_) );
XNOR2X1 XNOR2X1_140 ( .A(_1833_), .B(_1832_), .Y(micro_ucr_hash1_b_17__4_) );
NAND2X1 NAND2X1_305 ( .A(_1832_), .B(_1833_), .Y(_1834_) );
OR2X2 OR2X2_121 ( .A(gnd), .B(micro_ucr_hash1_a_15__1_), .Y(_1835_) );
NAND2X1 NAND2X1_306 ( .A(gnd), .B(micro_ucr_hash1_a_15__1_), .Y(_1836_) );
NAND3X1 NAND3X1_275 ( .A(micro_ucr_hash1_W_16__1_), .B(_1836_), .C(_1835_), .Y(_1837_) );
INVX1 INVX1_176 ( .A(micro_ucr_hash1_W_16__1_), .Y(_1838_) );
NOR2X1 NOR2X1_168 ( .A(gnd), .B(micro_ucr_hash1_a_15__1_), .Y(_1839_) );
AND2X2 AND2X2_92 ( .A(gnd), .B(micro_ucr_hash1_a_15__1_), .Y(_1840_) );
OAI21X1 OAI21X1_263 ( .A(_1840_), .B(_1839_), .C(_1838_), .Y(_1841_) );
NAND2X1 NAND2X1_307 ( .A(_1841_), .B(_1837_), .Y(_1842_) );
XNOR2X1 XNOR2X1_141 ( .A(_1842_), .B(_1834_), .Y(micro_ucr_hash1_b_17__5_) );
NAND3X1 NAND3X1_276 ( .A(_1837_), .B(_1841_), .C(_1834_), .Y(_1843_) );
NOR3X1 NOR3X1_55 ( .A(_1838_), .B(_1839_), .C(_1840_), .Y(_1844_) );
INVX1 INVX1_177 ( .A(micro_ucr_hash1_W_16__2_), .Y(_1845_) );
NOR2X1 NOR2X1_169 ( .A(gnd), .B(micro_ucr_hash1_a_15__2_), .Y(_1846_) );
AND2X2 AND2X2_93 ( .A(gnd), .B(micro_ucr_hash1_a_15__2_), .Y(_1847_) );
NOR3X1 NOR3X1_56 ( .A(_1845_), .B(_1846_), .C(_1847_), .Y(_1848_) );
OR2X2 OR2X2_122 ( .A(gnd), .B(micro_ucr_hash1_a_15__2_), .Y(_1849_) );
NAND2X1 NAND2X1_308 ( .A(gnd), .B(micro_ucr_hash1_a_15__2_), .Y(_1850_) );
AOI21X1 AOI21X1_191 ( .A(_1850_), .B(_1849_), .C(micro_ucr_hash1_W_16__2_), .Y(_1851_) );
OAI21X1 OAI21X1_264 ( .A(_1848_), .B(_1851_), .C(_1844_), .Y(_1852_) );
NAND3X1 NAND3X1_277 ( .A(micro_ucr_hash1_W_16__2_), .B(_1850_), .C(_1849_), .Y(_1853_) );
OAI21X1 OAI21X1_265 ( .A(_1847_), .B(_1846_), .C(_1845_), .Y(_1854_) );
NAND3X1 NAND3X1_278 ( .A(_1854_), .B(_1837_), .C(_1853_), .Y(_1855_) );
NAND2X1 NAND2X1_309 ( .A(_1855_), .B(_1852_), .Y(_1856_) );
XNOR2X1 XNOR2X1_142 ( .A(_1856_), .B(_1843_), .Y(micro_ucr_hash1_b_17__6_) );
NAND3X1 NAND3X1_279 ( .A(_1853_), .B(_1854_), .C(_1844_), .Y(_1857_) );
OAI21X1 OAI21X1_266 ( .A(_1848_), .B(_1851_), .C(_1837_), .Y(_1858_) );
NAND2X1 NAND2X1_310 ( .A(_1857_), .B(_1858_), .Y(_1859_) );
OAI21X1 OAI21X1_267 ( .A(_1859_), .B(_1843_), .C(_1857_), .Y(_1860_) );
INVX1 INVX1_178 ( .A(micro_ucr_hash1_W_16__3_), .Y(_1861_) );
NOR2X1 NOR2X1_170 ( .A(gnd), .B(micro_ucr_hash1_a_15__3_), .Y(_1862_) );
AND2X2 AND2X2_94 ( .A(gnd), .B(micro_ucr_hash1_a_15__3_), .Y(_1863_) );
OAI21X1 OAI21X1_268 ( .A(_1863_), .B(_1862_), .C(_1861_), .Y(_1864_) );
OR2X2 OR2X2_123 ( .A(gnd), .B(micro_ucr_hash1_a_15__3_), .Y(_1865_) );
NAND2X1 NAND2X1_311 ( .A(gnd), .B(micro_ucr_hash1_a_15__3_), .Y(_1866_) );
NAND3X1 NAND3X1_280 ( .A(micro_ucr_hash1_W_16__3_), .B(_1866_), .C(_1865_), .Y(_1867_) );
AOI21X1 AOI21X1_192 ( .A(_1864_), .B(_1867_), .C(_1853_), .Y(_1868_) );
NAND3X1 NAND3X1_281 ( .A(_1861_), .B(_1866_), .C(_1865_), .Y(_1869_) );
OAI21X1 OAI21X1_269 ( .A(_1863_), .B(_1862_), .C(micro_ucr_hash1_W_16__3_), .Y(_1870_) );
AOI21X1 AOI21X1_193 ( .A(_1870_), .B(_1869_), .C(_1848_), .Y(_1871_) );
NOR2X1 NOR2X1_171 ( .A(_1868_), .B(_1871_), .Y(_1763_) );
XOR2X1 XOR2X1_160 ( .A(_1860_), .B(_1763_), .Y(micro_ucr_hash1_b_17__7_) );
INVX1 INVX1_179 ( .A(micro_ucr_hash1_W_16__4_), .Y(_1764_) );
OR2X2 OR2X2_124 ( .A(micro_ucr_hash1_b_15__4_), .B(micro_ucr_hash1_a_15__4_), .Y(_1765_) );
NAND2X1 NAND2X1_312 ( .A(micro_ucr_hash1_b_15__4_), .B(micro_ucr_hash1_a_15__4_), .Y(_1766_) );
NAND3X1 NAND3X1_282 ( .A(_1764_), .B(_1766_), .C(_1765_), .Y(_1767_) );
NOR2X1 NOR2X1_172 ( .A(micro_ucr_hash1_b_15__4_), .B(micro_ucr_hash1_a_15__4_), .Y(_1768_) );
AND2X2 AND2X2_95 ( .A(micro_ucr_hash1_b_15__4_), .B(micro_ucr_hash1_a_15__4_), .Y(_1769_) );
OAI21X1 OAI21X1_270 ( .A(_1769_), .B(_1768_), .C(micro_ucr_hash1_W_16__4_), .Y(_1770_) );
NAND3X1 NAND3X1_283 ( .A(_1864_), .B(_1767_), .C(_1770_), .Y(_1771_) );
AOI21X1 AOI21X1_194 ( .A(_1866_), .B(_1865_), .C(micro_ucr_hash1_W_16__3_), .Y(_1772_) );
OAI21X1 OAI21X1_271 ( .A(_1769_), .B(_1768_), .C(_1764_), .Y(_1773_) );
NAND3X1 NAND3X1_284 ( .A(micro_ucr_hash1_W_16__4_), .B(_1766_), .C(_1765_), .Y(_1774_) );
NAND3X1 NAND3X1_285 ( .A(_1773_), .B(_1774_), .C(_1772_), .Y(_1775_) );
AND2X2 AND2X2_96 ( .A(_1775_), .B(_1771_), .Y(_1776_) );
INVX2 INVX2_57 ( .A(_1871_), .Y(_1777_) );
NOR2X1 NOR2X1_173 ( .A(_1851_), .B(_1848_), .Y(_1778_) );
AOI21X1 AOI21X1_195 ( .A(_1844_), .B(_1778_), .C(_1868_), .Y(_1779_) );
OAI21X1 OAI21X1_272 ( .A(_1859_), .B(_1843_), .C(_1779_), .Y(_1780_) );
NAND2X1 NAND2X1_313 ( .A(_1777_), .B(_1780_), .Y(_1781_) );
XNOR2X1 XNOR2X1_143 ( .A(_1781_), .B(_1776_), .Y(micro_ucr_hash1_c_16__4_) );
NAND2X1 NAND2X1_314 ( .A(_1771_), .B(_1775_), .Y(_1782_) );
OAI21X1 OAI21X1_273 ( .A(_1781_), .B(_1782_), .C(_1771_), .Y(_1783_) );
INVX1 INVX1_180 ( .A(micro_ucr_hash1_W_16__5_), .Y(_1784_) );
OR2X2 OR2X2_125 ( .A(micro_ucr_hash1_b_15__5_), .B(micro_ucr_hash1_a_15__5_), .Y(_1785_) );
NAND2X1 NAND2X1_315 ( .A(micro_ucr_hash1_b_15__5_), .B(micro_ucr_hash1_a_15__5_), .Y(_1786_) );
NAND3X1 NAND3X1_286 ( .A(_1784_), .B(_1786_), .C(_1785_), .Y(_1787_) );
NOR2X1 NOR2X1_174 ( .A(micro_ucr_hash1_b_15__5_), .B(micro_ucr_hash1_a_15__5_), .Y(_1788_) );
AND2X2 AND2X2_97 ( .A(micro_ucr_hash1_b_15__5_), .B(micro_ucr_hash1_a_15__5_), .Y(_1789_) );
OAI21X1 OAI21X1_274 ( .A(_1789_), .B(_1788_), .C(micro_ucr_hash1_W_16__5_), .Y(_1790_) );
NAND3X1 NAND3X1_287 ( .A(_1773_), .B(_1790_), .C(_1787_), .Y(_1791_) );
AOI21X1 AOI21X1_196 ( .A(_1766_), .B(_1765_), .C(micro_ucr_hash1_W_16__4_), .Y(_1792_) );
NAND3X1 NAND3X1_288 ( .A(micro_ucr_hash1_W_16__5_), .B(_1786_), .C(_1785_), .Y(_1793_) );
OAI21X1 OAI21X1_275 ( .A(_1789_), .B(_1788_), .C(_1784_), .Y(_1794_) );
NAND3X1 NAND3X1_289 ( .A(_1794_), .B(_1793_), .C(_1792_), .Y(_1795_) );
NAND2X1 NAND2X1_316 ( .A(_1791_), .B(_1795_), .Y(_1796_) );
INVX2 INVX2_58 ( .A(_1796_), .Y(_1797_) );
XNOR2X1 XNOR2X1_144 ( .A(_1783_), .B(_1797_), .Y(micro_ucr_hash1_c_16__5_) );
AOI21X1 AOI21X1_197 ( .A(_1791_), .B(_1795_), .C(_1782_), .Y(_1798_) );
NAND3X1 NAND3X1_290 ( .A(_1777_), .B(_1798_), .C(_1780_), .Y(_1799_) );
NAND2X1 NAND2X1_317 ( .A(_1794_), .B(_1793_), .Y(_1800_) );
OR2X2 OR2X2_126 ( .A(_1800_), .B(_1792_), .Y(_1801_) );
INVX1 INVX1_181 ( .A(_1801_), .Y(_1802_) );
AOI21X1 AOI21X1_198 ( .A(_1792_), .B(_1800_), .C(_1771_), .Y(_1803_) );
NOR2X1 NOR2X1_175 ( .A(_1803_), .B(_1802_), .Y(_1804_) );
INVX1 INVX1_182 ( .A(micro_ucr_hash1_W_16__6_), .Y(_1805_) );
XNOR2X1 XNOR2X1_145 ( .A(micro_ucr_hash1_b_15__6_), .B(micro_ucr_hash1_a_15__6_), .Y(_1806_) );
OR2X2 OR2X2_127 ( .A(_1806_), .B(_1805_), .Y(_1807_) );
NAND2X1 NAND2X1_318 ( .A(_1805_), .B(_1806_), .Y(_1808_) );
NAND2X1 NAND2X1_319 ( .A(_1808_), .B(_1807_), .Y(_1809_) );
OR2X2 OR2X2_128 ( .A(_1809_), .B(_1793_), .Y(_1810_) );
NAND2X1 NAND2X1_320 ( .A(_1793_), .B(_1809_), .Y(_1811_) );
NAND2X1 NAND2X1_321 ( .A(_1811_), .B(_1810_), .Y(_1812_) );
AOI21X1 AOI21X1_199 ( .A(_1804_), .B(_1799_), .C(_1812_), .Y(_1813_) );
NAND2X1 NAND2X1_322 ( .A(_1796_), .B(_1776_), .Y(_1814_) );
OAI21X1 OAI21X1_276 ( .A(_1781_), .B(_1814_), .C(_1804_), .Y(_1815_) );
INVX1 INVX1_183 ( .A(_1812_), .Y(_1816_) );
NOR2X1 NOR2X1_176 ( .A(_1816_), .B(_1815_), .Y(_1817_) );
NOR2X1 NOR2X1_177 ( .A(_1813_), .B(_1817_), .Y(micro_ucr_hash1_c_16__6_) );
INVX1 INVX1_184 ( .A(_1857_), .Y(_1818_) );
AOI21X1 AOI21X1_200 ( .A(_1777_), .B(_1818_), .C(_1868_), .Y(_1819_) );
AOI21X1 AOI21X1_201 ( .A(_1832_), .B(_1833_), .C(_1842_), .Y(_1820_) );
NAND3X1 NAND3X1_291 ( .A(_1820_), .B(_1856_), .C(_1763_), .Y(_1821_) );
AOI21X1 AOI21X1_202 ( .A(_1819_), .B(_1821_), .C(_1814_), .Y(_1822_) );
OAI21X1 OAI21X1_277 ( .A(_1797_), .B(_1771_), .C(_1801_), .Y(_1823_) );
OAI21X1 OAI21X1_278 ( .A(_1822_), .B(_1823_), .C(_1816_), .Y(_1824_) );
XOR2X1 XOR2X1_161 ( .A(micro_ucr_hash1_b_15__7_), .B(micro_ucr_hash1_W_16__7_), .Y(_1825_) );
XNOR2X1 XNOR2X1_146 ( .A(_1825_), .B(micro_ucr_hash1_a_15__7_), .Y(_1826_) );
XNOR2X1 XNOR2X1_147 ( .A(_1826_), .B(_1807_), .Y(_1827_) );
NAND3X1 NAND3X1_292 ( .A(_1810_), .B(_1827_), .C(_1824_), .Y(_1828_) );
INVX1 INVX1_185 ( .A(_1810_), .Y(_1829_) );
INVX1 INVX1_186 ( .A(_1827_), .Y(_1830_) );
OAI21X1 OAI21X1_279 ( .A(_1813_), .B(_1829_), .C(_1830_), .Y(_1831_) );
NAND2X1 NAND2X1_323 ( .A(_1828_), .B(_1831_), .Y(micro_ucr_hash1_c_16__7_) );
XOR2X1 XOR2X1_162 ( .A(micro_ucr_hash1_b_17__4_), .B(gnd), .Y(micro_ucr_hash1_a_17__0_) );
XOR2X1 XOR2X1_163 ( .A(micro_ucr_hash1_b_17__5_), .B(gnd), .Y(micro_ucr_hash1_a_17__1_) );
XOR2X1 XOR2X1_164 ( .A(micro_ucr_hash1_b_17__6_), .B(gnd), .Y(micro_ucr_hash1_a_17__2_) );
XOR2X1 XOR2X1_165 ( .A(micro_ucr_hash1_b_17__7_), .B(gnd), .Y(micro_ucr_hash1_a_17__3_) );
XOR2X1 XOR2X1_166 ( .A(micro_ucr_hash1_c_16__4_), .B(micro_ucr_hash1_b_16__4_), .Y(micro_ucr_hash1_a_17__4_) );
XOR2X1 XOR2X1_167 ( .A(micro_ucr_hash1_c_16__5_), .B(micro_ucr_hash1_b_16__5_), .Y(micro_ucr_hash1_a_17__5_) );
XOR2X1 XOR2X1_168 ( .A(micro_ucr_hash1_c_16__6_), .B(micro_ucr_hash1_b_16__6_), .Y(micro_ucr_hash1_a_17__6_) );
XOR2X1 XOR2X1_169 ( .A(micro_ucr_hash1_c_16__7_), .B(micro_ucr_hash1_b_16__7_), .Y(micro_ucr_hash1_a_17__7_) );
INVX1 INVX1_187 ( .A(micro_ucr_hash1_W_17__0_), .Y(_1928_) );
NOR2X1 NOR2X1_178 ( .A(gnd), .B(micro_ucr_hash1_a_16__0_), .Y(_1929_) );
NAND2X1 NAND2X1_324 ( .A(_1928_), .B(_1929_), .Y(_1930_) );
OAI21X1 OAI21X1_280 ( .A(gnd), .B(micro_ucr_hash1_a_16__0_), .C(micro_ucr_hash1_W_17__0_), .Y(_1931_) );
NAND2X1 NAND2X1_325 ( .A(_1931_), .B(_1930_), .Y(micro_ucr_hash1_b_18__4_) );
OAI21X1 OAI21X1_281 ( .A(gnd), .B(micro_ucr_hash1_a_16__1_), .C(micro_ucr_hash1_W_17__1_), .Y(_1932_) );
INVX1 INVX1_188 ( .A(micro_ucr_hash1_W_17__1_), .Y(_1933_) );
NOR2X1 NOR2X1_179 ( .A(gnd), .B(micro_ucr_hash1_a_16__1_), .Y(_1934_) );
NAND2X1 NAND2X1_326 ( .A(_1933_), .B(_1934_), .Y(_1935_) );
NAND3X1 NAND3X1_293 ( .A(_1932_), .B(_1930_), .C(_1935_), .Y(_1936_) );
AND2X2 AND2X2_98 ( .A(_1929_), .B(_1928_), .Y(_1937_) );
INVX2 INVX2_59 ( .A(_1932_), .Y(_1938_) );
AND2X2 AND2X2_99 ( .A(_1934_), .B(_1933_), .Y(_1939_) );
OAI21X1 OAI21X1_282 ( .A(_1939_), .B(_1938_), .C(_1937_), .Y(_1940_) );
AND2X2 AND2X2_100 ( .A(_1940_), .B(_1936_), .Y(micro_ucr_hash1_b_18__5_) );
OAI21X1 OAI21X1_283 ( .A(gnd), .B(micro_ucr_hash1_a_16__2_), .C(micro_ucr_hash1_W_17__2_), .Y(_1941_) );
INVX1 INVX1_189 ( .A(micro_ucr_hash1_W_17__2_), .Y(_1942_) );
NOR2X1 NOR2X1_180 ( .A(gnd), .B(micro_ucr_hash1_a_16__2_), .Y(_1943_) );
NAND2X1 NAND2X1_327 ( .A(_1942_), .B(_1943_), .Y(_1944_) );
NAND2X1 NAND2X1_328 ( .A(_1941_), .B(_1944_), .Y(_1945_) );
NAND3X1 NAND3X1_294 ( .A(_1941_), .B(_1944_), .C(_1938_), .Y(_1946_) );
OAI21X1 OAI21X1_284 ( .A(_1936_), .B(_1945_), .C(_1946_), .Y(_1947_) );
INVX1 INVX1_190 ( .A(_1945_), .Y(_1948_) );
OAI21X1 OAI21X1_285 ( .A(_1937_), .B(_1939_), .C(_1932_), .Y(_1949_) );
NOR2X1 NOR2X1_181 ( .A(_1949_), .B(_1948_), .Y(_1950_) );
NOR2X1 NOR2X1_182 ( .A(_1947_), .B(_1950_), .Y(micro_ucr_hash1_b_18__6_) );
INVX1 INVX1_191 ( .A(micro_ucr_hash1_W_17__3_), .Y(_1951_) );
OAI21X1 OAI21X1_286 ( .A(gnd), .B(micro_ucr_hash1_a_16__3_), .C(_1951_), .Y(_1952_) );
NOR2X1 NOR2X1_183 ( .A(gnd), .B(micro_ucr_hash1_a_16__3_), .Y(_1953_) );
NAND2X1 NAND2X1_329 ( .A(micro_ucr_hash1_W_17__3_), .B(_1953_), .Y(_1954_) );
NAND3X1 NAND3X1_295 ( .A(_1941_), .B(_1952_), .C(_1954_), .Y(_1955_) );
INVX1 INVX1_192 ( .A(_1941_), .Y(_1956_) );
OAI21X1 OAI21X1_287 ( .A(gnd), .B(micro_ucr_hash1_a_16__3_), .C(micro_ucr_hash1_W_17__3_), .Y(_1957_) );
NAND2X1 NAND2X1_330 ( .A(_1951_), .B(_1953_), .Y(_1958_) );
NAND3X1 NAND3X1_296 ( .A(_1957_), .B(_1958_), .C(_1956_), .Y(_1959_) );
NAND2X1 NAND2X1_331 ( .A(_1955_), .B(_1959_), .Y(_1960_) );
XNOR2X1 XNOR2X1_148 ( .A(_1947_), .B(_1960_), .Y(micro_ucr_hash1_b_18__7_) );
INVX1 INVX1_193 ( .A(_1957_), .Y(_1961_) );
OAI21X1 OAI21X1_288 ( .A(micro_ucr_hash1_b_16__4_), .B(micro_ucr_hash1_a_16__4_), .C(micro_ucr_hash1_W_17__4_), .Y(_1962_) );
INVX1 INVX1_194 ( .A(micro_ucr_hash1_b_16__4_), .Y(_1963_) );
INVX1 INVX1_195 ( .A(micro_ucr_hash1_a_16__4_), .Y(_1964_) );
INVX1 INVX1_196 ( .A(micro_ucr_hash1_W_17__4_), .Y(_1965_) );
NAND3X1 NAND3X1_297 ( .A(_1963_), .B(_1964_), .C(_1965_), .Y(_1966_) );
AOI21X1 AOI21X1_203 ( .A(_1962_), .B(_1966_), .C(_1961_), .Y(_1872_) );
OAI21X1 OAI21X1_289 ( .A(micro_ucr_hash1_b_16__4_), .B(micro_ucr_hash1_a_16__4_), .C(_1965_), .Y(_1873_) );
NAND3X1 NAND3X1_298 ( .A(micro_ucr_hash1_W_17__4_), .B(_1963_), .C(_1964_), .Y(_1874_) );
AOI21X1 AOI21X1_204 ( .A(_1873_), .B(_1874_), .C(_1957_), .Y(_1875_) );
NOR2X1 NOR2X1_184 ( .A(_1875_), .B(_1872_), .Y(_1876_) );
AOI21X1 AOI21X1_205 ( .A(_1957_), .B(_1958_), .C(_1956_), .Y(_1877_) );
OAI21X1 OAI21X1_290 ( .A(_1877_), .B(_1946_), .C(_1959_), .Y(_1878_) );
NOR3X1 NOR3X1_57 ( .A(_1936_), .B(_1945_), .C(_1877_), .Y(_1879_) );
NOR2X1 NOR2X1_185 ( .A(_1878_), .B(_1879_), .Y(_1880_) );
XNOR2X1 XNOR2X1_149 ( .A(_1880_), .B(_1876_), .Y(micro_ucr_hash1_c_17__4_) );
NAND3X1 NAND3X1_299 ( .A(_1962_), .B(_1966_), .C(_1961_), .Y(_1881_) );
OAI21X1 OAI21X1_291 ( .A(_1880_), .B(_1872_), .C(_1881_), .Y(_1882_) );
INVX1 INVX1_197 ( .A(micro_ucr_hash1_W_17__5_), .Y(_1883_) );
OAI21X1 OAI21X1_292 ( .A(micro_ucr_hash1_b_16__5_), .B(micro_ucr_hash1_a_16__5_), .C(_1883_), .Y(_1884_) );
NOR2X1 NOR2X1_186 ( .A(micro_ucr_hash1_b_16__5_), .B(micro_ucr_hash1_a_16__5_), .Y(_1885_) );
NAND2X1 NAND2X1_332 ( .A(micro_ucr_hash1_W_17__5_), .B(_1885_), .Y(_1886_) );
NAND3X1 NAND3X1_300 ( .A(_1962_), .B(_1884_), .C(_1886_), .Y(_1887_) );
INVX1 INVX1_198 ( .A(_1962_), .Y(_1888_) );
NAND2X1 NAND2X1_333 ( .A(_1883_), .B(_1885_), .Y(_1889_) );
OAI21X1 OAI21X1_293 ( .A(micro_ucr_hash1_b_16__5_), .B(micro_ucr_hash1_a_16__5_), .C(micro_ucr_hash1_W_17__5_), .Y(_1890_) );
NAND3X1 NAND3X1_301 ( .A(_1890_), .B(_1889_), .C(_1888_), .Y(_1891_) );
NAND2X1 NAND2X1_334 ( .A(_1887_), .B(_1891_), .Y(_1892_) );
XOR2X1 XOR2X1_170 ( .A(_1882_), .B(_1892_), .Y(micro_ucr_hash1_c_17__5_) );
OAI21X1 OAI21X1_294 ( .A(gnd), .B(micro_ucr_hash1_a_16__2_), .C(_1942_), .Y(_1893_) );
NAND2X1 NAND2X1_335 ( .A(micro_ucr_hash1_W_17__2_), .B(_1943_), .Y(_1894_) );
AOI21X1 AOI21X1_206 ( .A(_1893_), .B(_1894_), .C(_1932_), .Y(_1895_) );
INVX1 INVX1_199 ( .A(_1959_), .Y(_1896_) );
AOI21X1 AOI21X1_207 ( .A(_1955_), .B(_1895_), .C(_1896_), .Y(_1897_) );
NOR3X1 NOR3X1_58 ( .A(_1937_), .B(_1938_), .C(_1939_), .Y(_1898_) );
NAND3X1 NAND3X1_302 ( .A(_1948_), .B(_1955_), .C(_1898_), .Y(_1899_) );
NAND2X1 NAND2X1_336 ( .A(_1892_), .B(_1876_), .Y(_1900_) );
AOI21X1 AOI21X1_208 ( .A(_1897_), .B(_1899_), .C(_1900_), .Y(_1901_) );
AOI22X1 AOI22X1_8 ( .A(_1889_), .B(_1890_), .C(_1881_), .D(_1962_), .Y(_1902_) );
INVX1 INVX1_200 ( .A(_1889_), .Y(_1903_) );
OAI21X1 OAI21X1_295 ( .A(micro_ucr_hash1_b_16__6_), .B(micro_ucr_hash1_a_16__6_), .C(micro_ucr_hash1_W_17__6_), .Y(_1904_) );
INVX1 INVX1_201 ( .A(micro_ucr_hash1_W_17__6_), .Y(_1905_) );
NOR2X1 NOR2X1_187 ( .A(micro_ucr_hash1_b_16__6_), .B(micro_ucr_hash1_a_16__6_), .Y(_1906_) );
NAND2X1 NAND2X1_337 ( .A(_1905_), .B(_1906_), .Y(_1907_) );
NAND2X1 NAND2X1_338 ( .A(_1904_), .B(_1907_), .Y(_1908_) );
NOR2X1 NOR2X1_188 ( .A(_1903_), .B(_1908_), .Y(_1909_) );
INVX1 INVX1_202 ( .A(_1909_), .Y(_1910_) );
NAND2X1 NAND2X1_339 ( .A(_1903_), .B(_1908_), .Y(_1911_) );
NAND2X1 NAND2X1_340 ( .A(_1911_), .B(_1910_), .Y(_1912_) );
INVX1 INVX1_203 ( .A(_1912_), .Y(_1913_) );
OAI21X1 OAI21X1_296 ( .A(_1901_), .B(_1902_), .C(_1913_), .Y(_1914_) );
NAND3X1 NAND3X1_303 ( .A(_1957_), .B(_1873_), .C(_1874_), .Y(_1915_) );
NAND2X1 NAND2X1_341 ( .A(_1915_), .B(_1881_), .Y(_1916_) );
AOI21X1 AOI21X1_209 ( .A(_1887_), .B(_1891_), .C(_1916_), .Y(_1917_) );
OAI21X1 OAI21X1_297 ( .A(_1878_), .B(_1879_), .C(_1917_), .Y(_1918_) );
INVX1 INVX1_204 ( .A(_1902_), .Y(_1919_) );
NAND3X1 NAND3X1_304 ( .A(_1919_), .B(_1912_), .C(_1918_), .Y(_1920_) );
AND2X2 AND2X2_101 ( .A(_1914_), .B(_1920_), .Y(micro_ucr_hash1_c_17__6_) );
AOI21X1 AOI21X1_210 ( .A(_1919_), .B(_1918_), .C(_1912_), .Y(_1921_) );
NOR2X1 NOR2X1_189 ( .A(micro_ucr_hash1_b_16__7_), .B(micro_ucr_hash1_a_16__7_), .Y(_1922_) );
XNOR2X1 XNOR2X1_150 ( .A(_1922_), .B(micro_ucr_hash1_W_17__7_), .Y(_1923_) );
XNOR2X1 XNOR2X1_151 ( .A(_1923_), .B(_1904_), .Y(_1924_) );
OAI21X1 OAI21X1_298 ( .A(_1921_), .B(_1909_), .C(_1924_), .Y(_1925_) );
INVX1 INVX1_205 ( .A(_1924_), .Y(_1926_) );
NAND3X1 NAND3X1_305 ( .A(_1910_), .B(_1926_), .C(_1914_), .Y(_1927_) );
NAND2X1 NAND2X1_342 ( .A(_1925_), .B(_1927_), .Y(micro_ucr_hash1_c_17__7_) );
XOR2X1 XOR2X1_171 ( .A(micro_ucr_hash1_b_18__4_), .B(gnd), .Y(micro_ucr_hash1_a_18__0_) );
XOR2X1 XOR2X1_172 ( .A(micro_ucr_hash1_b_18__5_), .B(gnd), .Y(micro_ucr_hash1_a_18__1_) );
XOR2X1 XOR2X1_173 ( .A(micro_ucr_hash1_b_18__6_), .B(gnd), .Y(micro_ucr_hash1_a_18__2_) );
XOR2X1 XOR2X1_174 ( .A(micro_ucr_hash1_b_18__7_), .B(gnd), .Y(micro_ucr_hash1_a_18__3_) );
XOR2X1 XOR2X1_175 ( .A(micro_ucr_hash1_c_17__4_), .B(micro_ucr_hash1_b_17__4_), .Y(micro_ucr_hash1_a_18__4_) );
XOR2X1 XOR2X1_176 ( .A(micro_ucr_hash1_c_17__5_), .B(micro_ucr_hash1_b_17__5_), .Y(micro_ucr_hash1_a_18__5_) );
XOR2X1 XOR2X1_177 ( .A(micro_ucr_hash1_c_17__6_), .B(micro_ucr_hash1_b_17__6_), .Y(micro_ucr_hash1_a_18__6_) );
XOR2X1 XOR2X1_178 ( .A(micro_ucr_hash1_c_17__7_), .B(micro_ucr_hash1_b_17__7_), .Y(micro_ucr_hash1_a_18__7_) );
INVX1 INVX1_206 ( .A(micro_ucr_hash1_W_18__0_), .Y(_2023_) );
NOR2X1 NOR2X1_190 ( .A(gnd), .B(micro_ucr_hash1_a_17__0_), .Y(_2024_) );
NAND2X1 NAND2X1_343 ( .A(_2023_), .B(_2024_), .Y(_2025_) );
OAI21X1 OAI21X1_299 ( .A(gnd), .B(micro_ucr_hash1_a_17__0_), .C(micro_ucr_hash1_W_18__0_), .Y(_2026_) );
NAND2X1 NAND2X1_344 ( .A(_2026_), .B(_2025_), .Y(micro_ucr_hash1_b_19__4_) );
OAI21X1 OAI21X1_300 ( .A(gnd), .B(micro_ucr_hash1_a_17__1_), .C(micro_ucr_hash1_W_18__1_), .Y(_2027_) );
INVX1 INVX1_207 ( .A(micro_ucr_hash1_W_18__1_), .Y(_2028_) );
NOR2X1 NOR2X1_191 ( .A(gnd), .B(micro_ucr_hash1_a_17__1_), .Y(_2029_) );
NAND2X1 NAND2X1_345 ( .A(_2028_), .B(_2029_), .Y(_2030_) );
NAND3X1 NAND3X1_306 ( .A(_2027_), .B(_2025_), .C(_2030_), .Y(_2031_) );
AND2X2 AND2X2_102 ( .A(_2024_), .B(_2023_), .Y(_2032_) );
INVX2 INVX2_60 ( .A(_2027_), .Y(_2033_) );
AND2X2 AND2X2_103 ( .A(_2029_), .B(_2028_), .Y(_2034_) );
OAI21X1 OAI21X1_301 ( .A(_2034_), .B(_2033_), .C(_2032_), .Y(_2035_) );
AND2X2 AND2X2_104 ( .A(_2035_), .B(_2031_), .Y(micro_ucr_hash1_b_19__5_) );
OAI21X1 OAI21X1_302 ( .A(gnd), .B(micro_ucr_hash1_a_17__2_), .C(micro_ucr_hash1_W_18__2_), .Y(_2036_) );
INVX1 INVX1_208 ( .A(micro_ucr_hash1_W_18__2_), .Y(_2037_) );
NOR2X1 NOR2X1_192 ( .A(gnd), .B(micro_ucr_hash1_a_17__2_), .Y(_2038_) );
NAND2X1 NAND2X1_346 ( .A(_2037_), .B(_2038_), .Y(_2039_) );
NAND2X1 NAND2X1_347 ( .A(_2036_), .B(_2039_), .Y(_2040_) );
NAND3X1 NAND3X1_307 ( .A(_2036_), .B(_2039_), .C(_2033_), .Y(_2041_) );
OAI21X1 OAI21X1_303 ( .A(_2031_), .B(_2040_), .C(_2041_), .Y(_2042_) );
INVX1 INVX1_209 ( .A(_2040_), .Y(_2043_) );
OAI21X1 OAI21X1_304 ( .A(_2032_), .B(_2034_), .C(_2027_), .Y(_2044_) );
NOR2X1 NOR2X1_193 ( .A(_2044_), .B(_2043_), .Y(_2045_) );
NOR2X1 NOR2X1_194 ( .A(_2042_), .B(_2045_), .Y(micro_ucr_hash1_b_19__6_) );
INVX1 INVX1_210 ( .A(micro_ucr_hash1_W_18__3_), .Y(_2046_) );
OAI21X1 OAI21X1_305 ( .A(gnd), .B(micro_ucr_hash1_a_17__3_), .C(_2046_), .Y(_2047_) );
NOR2X1 NOR2X1_195 ( .A(gnd), .B(micro_ucr_hash1_a_17__3_), .Y(_2048_) );
NAND2X1 NAND2X1_348 ( .A(micro_ucr_hash1_W_18__3_), .B(_2048_), .Y(_2049_) );
NAND3X1 NAND3X1_308 ( .A(_2036_), .B(_2047_), .C(_2049_), .Y(_2050_) );
INVX1 INVX1_211 ( .A(_2036_), .Y(_2051_) );
OAI21X1 OAI21X1_306 ( .A(gnd), .B(micro_ucr_hash1_a_17__3_), .C(micro_ucr_hash1_W_18__3_), .Y(_2052_) );
NAND2X1 NAND2X1_349 ( .A(_2046_), .B(_2048_), .Y(_2053_) );
NAND3X1 NAND3X1_309 ( .A(_2052_), .B(_2053_), .C(_2051_), .Y(_2054_) );
NAND2X1 NAND2X1_350 ( .A(_2050_), .B(_2054_), .Y(_2055_) );
XNOR2X1 XNOR2X1_152 ( .A(_2042_), .B(_2055_), .Y(micro_ucr_hash1_b_19__7_) );
INVX1 INVX1_212 ( .A(_2052_), .Y(_2056_) );
OAI21X1 OAI21X1_307 ( .A(micro_ucr_hash1_b_17__4_), .B(micro_ucr_hash1_a_17__4_), .C(micro_ucr_hash1_W_18__4_), .Y(_2057_) );
INVX1 INVX1_213 ( .A(micro_ucr_hash1_b_17__4_), .Y(_2058_) );
INVX1 INVX1_214 ( .A(micro_ucr_hash1_a_17__4_), .Y(_2059_) );
INVX1 INVX1_215 ( .A(micro_ucr_hash1_W_18__4_), .Y(_2060_) );
NAND3X1 NAND3X1_310 ( .A(_2058_), .B(_2059_), .C(_2060_), .Y(_2061_) );
AOI21X1 AOI21X1_211 ( .A(_2057_), .B(_2061_), .C(_2056_), .Y(_1967_) );
OAI21X1 OAI21X1_308 ( .A(micro_ucr_hash1_b_17__4_), .B(micro_ucr_hash1_a_17__4_), .C(_2060_), .Y(_1968_) );
NAND3X1 NAND3X1_311 ( .A(micro_ucr_hash1_W_18__4_), .B(_2058_), .C(_2059_), .Y(_1969_) );
AOI21X1 AOI21X1_212 ( .A(_1968_), .B(_1969_), .C(_2052_), .Y(_1970_) );
NOR2X1 NOR2X1_196 ( .A(_1970_), .B(_1967_), .Y(_1971_) );
AOI21X1 AOI21X1_213 ( .A(_2052_), .B(_2053_), .C(_2051_), .Y(_1972_) );
OAI21X1 OAI21X1_309 ( .A(_1972_), .B(_2041_), .C(_2054_), .Y(_1973_) );
NOR3X1 NOR3X1_59 ( .A(_2031_), .B(_2040_), .C(_1972_), .Y(_1974_) );
NOR2X1 NOR2X1_197 ( .A(_1973_), .B(_1974_), .Y(_1975_) );
XNOR2X1 XNOR2X1_153 ( .A(_1975_), .B(_1971_), .Y(micro_ucr_hash1_c_18__4_) );
NAND3X1 NAND3X1_312 ( .A(_2057_), .B(_2061_), .C(_2056_), .Y(_1976_) );
OAI21X1 OAI21X1_310 ( .A(_1975_), .B(_1967_), .C(_1976_), .Y(_1977_) );
INVX1 INVX1_216 ( .A(micro_ucr_hash1_W_18__5_), .Y(_1978_) );
OAI21X1 OAI21X1_311 ( .A(micro_ucr_hash1_b_17__5_), .B(micro_ucr_hash1_a_17__5_), .C(_1978_), .Y(_1979_) );
NOR2X1 NOR2X1_198 ( .A(micro_ucr_hash1_b_17__5_), .B(micro_ucr_hash1_a_17__5_), .Y(_1980_) );
NAND2X1 NAND2X1_351 ( .A(micro_ucr_hash1_W_18__5_), .B(_1980_), .Y(_1981_) );
NAND3X1 NAND3X1_313 ( .A(_2057_), .B(_1979_), .C(_1981_), .Y(_1982_) );
INVX1 INVX1_217 ( .A(_2057_), .Y(_1983_) );
NAND2X1 NAND2X1_352 ( .A(_1978_), .B(_1980_), .Y(_1984_) );
OAI21X1 OAI21X1_312 ( .A(micro_ucr_hash1_b_17__5_), .B(micro_ucr_hash1_a_17__5_), .C(micro_ucr_hash1_W_18__5_), .Y(_1985_) );
NAND3X1 NAND3X1_314 ( .A(_1985_), .B(_1984_), .C(_1983_), .Y(_1986_) );
NAND2X1 NAND2X1_353 ( .A(_1982_), .B(_1986_), .Y(_1987_) );
XOR2X1 XOR2X1_179 ( .A(_1977_), .B(_1987_), .Y(micro_ucr_hash1_c_18__5_) );
OAI21X1 OAI21X1_313 ( .A(gnd), .B(micro_ucr_hash1_a_17__2_), .C(_2037_), .Y(_1988_) );
NAND2X1 NAND2X1_354 ( .A(micro_ucr_hash1_W_18__2_), .B(_2038_), .Y(_1989_) );
AOI21X1 AOI21X1_214 ( .A(_1988_), .B(_1989_), .C(_2027_), .Y(_1990_) );
INVX1 INVX1_218 ( .A(_2054_), .Y(_1991_) );
AOI21X1 AOI21X1_215 ( .A(_2050_), .B(_1990_), .C(_1991_), .Y(_1992_) );
NOR3X1 NOR3X1_60 ( .A(_2032_), .B(_2033_), .C(_2034_), .Y(_1993_) );
NAND3X1 NAND3X1_315 ( .A(_2043_), .B(_2050_), .C(_1993_), .Y(_1994_) );
NAND2X1 NAND2X1_355 ( .A(_1987_), .B(_1971_), .Y(_1995_) );
AOI21X1 AOI21X1_216 ( .A(_1992_), .B(_1994_), .C(_1995_), .Y(_1996_) );
AOI22X1 AOI22X1_9 ( .A(_1984_), .B(_1985_), .C(_1976_), .D(_2057_), .Y(_1997_) );
INVX1 INVX1_219 ( .A(_1984_), .Y(_1998_) );
OAI21X1 OAI21X1_314 ( .A(micro_ucr_hash1_b_17__6_), .B(micro_ucr_hash1_a_17__6_), .C(micro_ucr_hash1_W_18__6_), .Y(_1999_) );
INVX1 INVX1_220 ( .A(micro_ucr_hash1_W_18__6_), .Y(_2000_) );
NOR2X1 NOR2X1_199 ( .A(micro_ucr_hash1_b_17__6_), .B(micro_ucr_hash1_a_17__6_), .Y(_2001_) );
NAND2X1 NAND2X1_356 ( .A(_2000_), .B(_2001_), .Y(_2002_) );
NAND2X1 NAND2X1_357 ( .A(_1999_), .B(_2002_), .Y(_2003_) );
NOR2X1 NOR2X1_200 ( .A(_1998_), .B(_2003_), .Y(_2004_) );
INVX1 INVX1_221 ( .A(_2004_), .Y(_2005_) );
NAND2X1 NAND2X1_358 ( .A(_1998_), .B(_2003_), .Y(_2006_) );
NAND2X1 NAND2X1_359 ( .A(_2006_), .B(_2005_), .Y(_2007_) );
INVX1 INVX1_222 ( .A(_2007_), .Y(_2008_) );
OAI21X1 OAI21X1_315 ( .A(_1996_), .B(_1997_), .C(_2008_), .Y(_2009_) );
NAND3X1 NAND3X1_316 ( .A(_2052_), .B(_1968_), .C(_1969_), .Y(_2010_) );
NAND2X1 NAND2X1_360 ( .A(_2010_), .B(_1976_), .Y(_2011_) );
AOI21X1 AOI21X1_217 ( .A(_1982_), .B(_1986_), .C(_2011_), .Y(_2012_) );
OAI21X1 OAI21X1_316 ( .A(_1973_), .B(_1974_), .C(_2012_), .Y(_2013_) );
INVX1 INVX1_223 ( .A(_1997_), .Y(_2014_) );
NAND3X1 NAND3X1_317 ( .A(_2014_), .B(_2007_), .C(_2013_), .Y(_2015_) );
AND2X2 AND2X2_105 ( .A(_2009_), .B(_2015_), .Y(micro_ucr_hash1_c_18__6_) );
AOI21X1 AOI21X1_218 ( .A(_2014_), .B(_2013_), .C(_2007_), .Y(_2016_) );
NOR2X1 NOR2X1_201 ( .A(micro_ucr_hash1_b_17__7_), .B(micro_ucr_hash1_a_17__7_), .Y(_2017_) );
XNOR2X1 XNOR2X1_154 ( .A(_2017_), .B(micro_ucr_hash1_W_18__7_), .Y(_2018_) );
XNOR2X1 XNOR2X1_155 ( .A(_2018_), .B(_1999_), .Y(_2019_) );
OAI21X1 OAI21X1_317 ( .A(_2016_), .B(_2004_), .C(_2019_), .Y(_2020_) );
INVX1 INVX1_224 ( .A(_2019_), .Y(_2021_) );
NAND3X1 NAND3X1_318 ( .A(_2005_), .B(_2021_), .C(_2009_), .Y(_2022_) );
NAND2X1 NAND2X1_361 ( .A(_2020_), .B(_2022_), .Y(micro_ucr_hash1_c_18__7_) );
XOR2X1 XOR2X1_180 ( .A(micro_ucr_hash1_b_19__4_), .B(gnd), .Y(micro_ucr_hash1_a_19__0_) );
XOR2X1 XOR2X1_181 ( .A(micro_ucr_hash1_b_19__5_), .B(gnd), .Y(micro_ucr_hash1_a_19__1_) );
XOR2X1 XOR2X1_182 ( .A(micro_ucr_hash1_b_19__6_), .B(gnd), .Y(micro_ucr_hash1_a_19__2_) );
XOR2X1 XOR2X1_183 ( .A(micro_ucr_hash1_b_19__7_), .B(gnd), .Y(micro_ucr_hash1_a_19__3_) );
XOR2X1 XOR2X1_184 ( .A(micro_ucr_hash1_c_18__4_), .B(micro_ucr_hash1_b_18__4_), .Y(micro_ucr_hash1_a_19__4_) );
XOR2X1 XOR2X1_185 ( .A(micro_ucr_hash1_c_18__5_), .B(micro_ucr_hash1_b_18__5_), .Y(micro_ucr_hash1_a_19__5_) );
XOR2X1 XOR2X1_186 ( .A(micro_ucr_hash1_c_18__6_), .B(micro_ucr_hash1_b_18__6_), .Y(micro_ucr_hash1_a_19__6_) );
XOR2X1 XOR2X1_187 ( .A(micro_ucr_hash1_c_18__7_), .B(micro_ucr_hash1_b_18__7_), .Y(micro_ucr_hash1_a_19__7_) );
INVX1 INVX1_225 ( .A(micro_ucr_hash1_W_19__0_), .Y(_2118_) );
NOR2X1 NOR2X1_202 ( .A(gnd), .B(micro_ucr_hash1_a_18__0_), .Y(_2119_) );
NAND2X1 NAND2X1_362 ( .A(_2118_), .B(_2119_), .Y(_2120_) );
OAI21X1 OAI21X1_318 ( .A(gnd), .B(micro_ucr_hash1_a_18__0_), .C(micro_ucr_hash1_W_19__0_), .Y(_2121_) );
NAND2X1 NAND2X1_363 ( .A(_2121_), .B(_2120_), .Y(micro_ucr_hash1_b_20__4_) );
OAI21X1 OAI21X1_319 ( .A(gnd), .B(micro_ucr_hash1_a_18__1_), .C(micro_ucr_hash1_W_19__1_), .Y(_2122_) );
INVX1 INVX1_226 ( .A(micro_ucr_hash1_W_19__1_), .Y(_2123_) );
NOR2X1 NOR2X1_203 ( .A(gnd), .B(micro_ucr_hash1_a_18__1_), .Y(_2124_) );
NAND2X1 NAND2X1_364 ( .A(_2123_), .B(_2124_), .Y(_2125_) );
NAND3X1 NAND3X1_319 ( .A(_2122_), .B(_2120_), .C(_2125_), .Y(_2126_) );
AND2X2 AND2X2_106 ( .A(_2119_), .B(_2118_), .Y(_2127_) );
INVX2 INVX2_61 ( .A(_2122_), .Y(_2128_) );
AND2X2 AND2X2_107 ( .A(_2124_), .B(_2123_), .Y(_2129_) );
OAI21X1 OAI21X1_320 ( .A(_2129_), .B(_2128_), .C(_2127_), .Y(_2130_) );
AND2X2 AND2X2_108 ( .A(_2130_), .B(_2126_), .Y(micro_ucr_hash1_b_20__5_) );
OAI21X1 OAI21X1_321 ( .A(gnd), .B(micro_ucr_hash1_a_18__2_), .C(micro_ucr_hash1_W_19__2_), .Y(_2131_) );
INVX1 INVX1_227 ( .A(micro_ucr_hash1_W_19__2_), .Y(_2132_) );
NOR2X1 NOR2X1_204 ( .A(gnd), .B(micro_ucr_hash1_a_18__2_), .Y(_2133_) );
NAND2X1 NAND2X1_365 ( .A(_2132_), .B(_2133_), .Y(_2134_) );
NAND2X1 NAND2X1_366 ( .A(_2131_), .B(_2134_), .Y(_2135_) );
NAND3X1 NAND3X1_320 ( .A(_2131_), .B(_2134_), .C(_2128_), .Y(_2136_) );
OAI21X1 OAI21X1_322 ( .A(_2126_), .B(_2135_), .C(_2136_), .Y(_2137_) );
INVX1 INVX1_228 ( .A(_2135_), .Y(_2138_) );
OAI21X1 OAI21X1_323 ( .A(_2127_), .B(_2129_), .C(_2122_), .Y(_2139_) );
NOR2X1 NOR2X1_205 ( .A(_2139_), .B(_2138_), .Y(_2140_) );
NOR2X1 NOR2X1_206 ( .A(_2137_), .B(_2140_), .Y(micro_ucr_hash1_b_20__6_) );
INVX1 INVX1_229 ( .A(micro_ucr_hash1_W_19__3_), .Y(_2141_) );
OAI21X1 OAI21X1_324 ( .A(gnd), .B(micro_ucr_hash1_a_18__3_), .C(_2141_), .Y(_2142_) );
NOR2X1 NOR2X1_207 ( .A(gnd), .B(micro_ucr_hash1_a_18__3_), .Y(_2143_) );
NAND2X1 NAND2X1_367 ( .A(micro_ucr_hash1_W_19__3_), .B(_2143_), .Y(_2144_) );
NAND3X1 NAND3X1_321 ( .A(_2131_), .B(_2142_), .C(_2144_), .Y(_2145_) );
INVX1 INVX1_230 ( .A(_2131_), .Y(_2146_) );
OAI21X1 OAI21X1_325 ( .A(gnd), .B(micro_ucr_hash1_a_18__3_), .C(micro_ucr_hash1_W_19__3_), .Y(_2147_) );
NAND2X1 NAND2X1_368 ( .A(_2141_), .B(_2143_), .Y(_2148_) );
NAND3X1 NAND3X1_322 ( .A(_2147_), .B(_2148_), .C(_2146_), .Y(_2149_) );
NAND2X1 NAND2X1_369 ( .A(_2145_), .B(_2149_), .Y(_2150_) );
XNOR2X1 XNOR2X1_156 ( .A(_2137_), .B(_2150_), .Y(micro_ucr_hash1_b_20__7_) );
INVX1 INVX1_231 ( .A(_2147_), .Y(_2151_) );
OAI21X1 OAI21X1_326 ( .A(micro_ucr_hash1_b_18__4_), .B(micro_ucr_hash1_a_18__4_), .C(micro_ucr_hash1_W_19__4_), .Y(_2152_) );
INVX1 INVX1_232 ( .A(micro_ucr_hash1_b_18__4_), .Y(_2153_) );
INVX1 INVX1_233 ( .A(micro_ucr_hash1_a_18__4_), .Y(_2154_) );
INVX1 INVX1_234 ( .A(micro_ucr_hash1_W_19__4_), .Y(_2155_) );
NAND3X1 NAND3X1_323 ( .A(_2153_), .B(_2154_), .C(_2155_), .Y(_2156_) );
AOI21X1 AOI21X1_219 ( .A(_2152_), .B(_2156_), .C(_2151_), .Y(_2062_) );
OAI21X1 OAI21X1_327 ( .A(micro_ucr_hash1_b_18__4_), .B(micro_ucr_hash1_a_18__4_), .C(_2155_), .Y(_2063_) );
NAND3X1 NAND3X1_324 ( .A(micro_ucr_hash1_W_19__4_), .B(_2153_), .C(_2154_), .Y(_2064_) );
AOI21X1 AOI21X1_220 ( .A(_2063_), .B(_2064_), .C(_2147_), .Y(_2065_) );
NOR2X1 NOR2X1_208 ( .A(_2065_), .B(_2062_), .Y(_2066_) );
AOI21X1 AOI21X1_221 ( .A(_2147_), .B(_2148_), .C(_2146_), .Y(_2067_) );
OAI21X1 OAI21X1_328 ( .A(_2067_), .B(_2136_), .C(_2149_), .Y(_2068_) );
NOR3X1 NOR3X1_61 ( .A(_2126_), .B(_2135_), .C(_2067_), .Y(_2069_) );
NOR2X1 NOR2X1_209 ( .A(_2068_), .B(_2069_), .Y(_2070_) );
XNOR2X1 XNOR2X1_157 ( .A(_2070_), .B(_2066_), .Y(micro_ucr_hash1_c_19__4_) );
NAND3X1 NAND3X1_325 ( .A(_2152_), .B(_2156_), .C(_2151_), .Y(_2071_) );
OAI21X1 OAI21X1_329 ( .A(_2070_), .B(_2062_), .C(_2071_), .Y(_2072_) );
INVX1 INVX1_235 ( .A(micro_ucr_hash1_W_19__5_), .Y(_2073_) );
OAI21X1 OAI21X1_330 ( .A(micro_ucr_hash1_b_18__5_), .B(micro_ucr_hash1_a_18__5_), .C(_2073_), .Y(_2074_) );
NOR2X1 NOR2X1_210 ( .A(micro_ucr_hash1_b_18__5_), .B(micro_ucr_hash1_a_18__5_), .Y(_2075_) );
NAND2X1 NAND2X1_370 ( .A(micro_ucr_hash1_W_19__5_), .B(_2075_), .Y(_2076_) );
NAND3X1 NAND3X1_326 ( .A(_2152_), .B(_2074_), .C(_2076_), .Y(_2077_) );
INVX1 INVX1_236 ( .A(_2152_), .Y(_2078_) );
NAND2X1 NAND2X1_371 ( .A(_2073_), .B(_2075_), .Y(_2079_) );
OAI21X1 OAI21X1_331 ( .A(micro_ucr_hash1_b_18__5_), .B(micro_ucr_hash1_a_18__5_), .C(micro_ucr_hash1_W_19__5_), .Y(_2080_) );
NAND3X1 NAND3X1_327 ( .A(_2080_), .B(_2079_), .C(_2078_), .Y(_2081_) );
NAND2X1 NAND2X1_372 ( .A(_2077_), .B(_2081_), .Y(_2082_) );
XOR2X1 XOR2X1_188 ( .A(_2072_), .B(_2082_), .Y(micro_ucr_hash1_c_19__5_) );
OAI21X1 OAI21X1_332 ( .A(gnd), .B(micro_ucr_hash1_a_18__2_), .C(_2132_), .Y(_2083_) );
NAND2X1 NAND2X1_373 ( .A(micro_ucr_hash1_W_19__2_), .B(_2133_), .Y(_2084_) );
AOI21X1 AOI21X1_222 ( .A(_2083_), .B(_2084_), .C(_2122_), .Y(_2085_) );
INVX1 INVX1_237 ( .A(_2149_), .Y(_2086_) );
AOI21X1 AOI21X1_223 ( .A(_2145_), .B(_2085_), .C(_2086_), .Y(_2087_) );
NOR3X1 NOR3X1_62 ( .A(_2127_), .B(_2128_), .C(_2129_), .Y(_2088_) );
NAND3X1 NAND3X1_328 ( .A(_2138_), .B(_2145_), .C(_2088_), .Y(_2089_) );
NAND2X1 NAND2X1_374 ( .A(_2082_), .B(_2066_), .Y(_2090_) );
AOI21X1 AOI21X1_224 ( .A(_2087_), .B(_2089_), .C(_2090_), .Y(_2091_) );
AOI22X1 AOI22X1_10 ( .A(_2079_), .B(_2080_), .C(_2071_), .D(_2152_), .Y(_2092_) );
INVX1 INVX1_238 ( .A(_2079_), .Y(_2093_) );
OAI21X1 OAI21X1_333 ( .A(micro_ucr_hash1_b_18__6_), .B(micro_ucr_hash1_a_18__6_), .C(micro_ucr_hash1_W_19__6_), .Y(_2094_) );
INVX1 INVX1_239 ( .A(micro_ucr_hash1_W_19__6_), .Y(_2095_) );
NOR2X1 NOR2X1_211 ( .A(micro_ucr_hash1_b_18__6_), .B(micro_ucr_hash1_a_18__6_), .Y(_2096_) );
NAND2X1 NAND2X1_375 ( .A(_2095_), .B(_2096_), .Y(_2097_) );
NAND2X1 NAND2X1_376 ( .A(_2094_), .B(_2097_), .Y(_2098_) );
NOR2X1 NOR2X1_212 ( .A(_2093_), .B(_2098_), .Y(_2099_) );
INVX1 INVX1_240 ( .A(_2099_), .Y(_2100_) );
NAND2X1 NAND2X1_377 ( .A(_2093_), .B(_2098_), .Y(_2101_) );
NAND2X1 NAND2X1_378 ( .A(_2101_), .B(_2100_), .Y(_2102_) );
INVX1 INVX1_241 ( .A(_2102_), .Y(_2103_) );
OAI21X1 OAI21X1_334 ( .A(_2091_), .B(_2092_), .C(_2103_), .Y(_2104_) );
NAND3X1 NAND3X1_329 ( .A(_2147_), .B(_2063_), .C(_2064_), .Y(_2105_) );
NAND2X1 NAND2X1_379 ( .A(_2105_), .B(_2071_), .Y(_2106_) );
AOI21X1 AOI21X1_225 ( .A(_2077_), .B(_2081_), .C(_2106_), .Y(_2107_) );
OAI21X1 OAI21X1_335 ( .A(_2068_), .B(_2069_), .C(_2107_), .Y(_2108_) );
INVX1 INVX1_242 ( .A(_2092_), .Y(_2109_) );
NAND3X1 NAND3X1_330 ( .A(_2109_), .B(_2102_), .C(_2108_), .Y(_2110_) );
AND2X2 AND2X2_109 ( .A(_2104_), .B(_2110_), .Y(micro_ucr_hash1_c_19__6_) );
AOI21X1 AOI21X1_226 ( .A(_2109_), .B(_2108_), .C(_2102_), .Y(_2111_) );
NOR2X1 NOR2X1_213 ( .A(micro_ucr_hash1_b_18__7_), .B(micro_ucr_hash1_a_18__7_), .Y(_2112_) );
XNOR2X1 XNOR2X1_158 ( .A(_2112_), .B(micro_ucr_hash1_W_19__7_), .Y(_2113_) );
XNOR2X1 XNOR2X1_159 ( .A(_2113_), .B(_2094_), .Y(_2114_) );
OAI21X1 OAI21X1_336 ( .A(_2111_), .B(_2099_), .C(_2114_), .Y(_2115_) );
INVX1 INVX1_243 ( .A(_2114_), .Y(_2116_) );
NAND3X1 NAND3X1_331 ( .A(_2100_), .B(_2116_), .C(_2104_), .Y(_2117_) );
NAND2X1 NAND2X1_380 ( .A(_2115_), .B(_2117_), .Y(micro_ucr_hash1_c_19__7_) );
XOR2X1 XOR2X1_189 ( .A(micro_ucr_hash1_b_20__4_), .B(gnd), .Y(micro_ucr_hash1_a_20__0_) );
XOR2X1 XOR2X1_190 ( .A(micro_ucr_hash1_b_20__5_), .B(gnd), .Y(micro_ucr_hash1_a_20__1_) );
XOR2X1 XOR2X1_191 ( .A(micro_ucr_hash1_b_20__6_), .B(gnd), .Y(micro_ucr_hash1_a_20__2_) );
XOR2X1 XOR2X1_192 ( .A(micro_ucr_hash1_b_20__7_), .B(gnd), .Y(micro_ucr_hash1_a_20__3_) );
XOR2X1 XOR2X1_193 ( .A(micro_ucr_hash1_c_19__4_), .B(micro_ucr_hash1_b_19__4_), .Y(micro_ucr_hash1_a_20__4_) );
XOR2X1 XOR2X1_194 ( .A(micro_ucr_hash1_c_19__5_), .B(micro_ucr_hash1_b_19__5_), .Y(micro_ucr_hash1_a_20__5_) );
XOR2X1 XOR2X1_195 ( .A(micro_ucr_hash1_c_19__6_), .B(micro_ucr_hash1_b_19__6_), .Y(micro_ucr_hash1_a_20__6_) );
XOR2X1 XOR2X1_196 ( .A(micro_ucr_hash1_c_19__7_), .B(micro_ucr_hash1_b_19__7_), .Y(micro_ucr_hash1_a_20__7_) );
INVX1 INVX1_244 ( .A(micro_ucr_hash1_W_20__0_), .Y(_2213_) );
NOR2X1 NOR2X1_214 ( .A(gnd), .B(micro_ucr_hash1_a_19__0_), .Y(_2214_) );
NAND2X1 NAND2X1_381 ( .A(_2213_), .B(_2214_), .Y(_2215_) );
OAI21X1 OAI21X1_337 ( .A(gnd), .B(micro_ucr_hash1_a_19__0_), .C(micro_ucr_hash1_W_20__0_), .Y(_2216_) );
NAND2X1 NAND2X1_382 ( .A(_2216_), .B(_2215_), .Y(micro_ucr_hash1_b_21__4_) );
OAI21X1 OAI21X1_338 ( .A(gnd), .B(micro_ucr_hash1_a_19__1_), .C(micro_ucr_hash1_W_20__1_), .Y(_2217_) );
INVX1 INVX1_245 ( .A(micro_ucr_hash1_W_20__1_), .Y(_2218_) );
NOR2X1 NOR2X1_215 ( .A(gnd), .B(micro_ucr_hash1_a_19__1_), .Y(_2219_) );
NAND2X1 NAND2X1_383 ( .A(_2218_), .B(_2219_), .Y(_2220_) );
NAND3X1 NAND3X1_332 ( .A(_2217_), .B(_2215_), .C(_2220_), .Y(_2221_) );
AND2X2 AND2X2_110 ( .A(_2214_), .B(_2213_), .Y(_2222_) );
INVX2 INVX2_62 ( .A(_2217_), .Y(_2223_) );
AND2X2 AND2X2_111 ( .A(_2219_), .B(_2218_), .Y(_2224_) );
OAI21X1 OAI21X1_339 ( .A(_2224_), .B(_2223_), .C(_2222_), .Y(_2225_) );
AND2X2 AND2X2_112 ( .A(_2225_), .B(_2221_), .Y(micro_ucr_hash1_b_21__5_) );
OAI21X1 OAI21X1_340 ( .A(gnd), .B(micro_ucr_hash1_a_19__2_), .C(micro_ucr_hash1_W_20__2_), .Y(_2226_) );
INVX1 INVX1_246 ( .A(micro_ucr_hash1_W_20__2_), .Y(_2227_) );
NOR2X1 NOR2X1_216 ( .A(gnd), .B(micro_ucr_hash1_a_19__2_), .Y(_2228_) );
NAND2X1 NAND2X1_384 ( .A(_2227_), .B(_2228_), .Y(_2229_) );
NAND2X1 NAND2X1_385 ( .A(_2226_), .B(_2229_), .Y(_2230_) );
NAND3X1 NAND3X1_333 ( .A(_2226_), .B(_2229_), .C(_2223_), .Y(_2231_) );
OAI21X1 OAI21X1_341 ( .A(_2221_), .B(_2230_), .C(_2231_), .Y(_2232_) );
INVX1 INVX1_247 ( .A(_2230_), .Y(_2233_) );
OAI21X1 OAI21X1_342 ( .A(_2222_), .B(_2224_), .C(_2217_), .Y(_2234_) );
NOR2X1 NOR2X1_217 ( .A(_2234_), .B(_2233_), .Y(_2235_) );
NOR2X1 NOR2X1_218 ( .A(_2232_), .B(_2235_), .Y(micro_ucr_hash1_b_21__6_) );
INVX1 INVX1_248 ( .A(micro_ucr_hash1_W_20__3_), .Y(_2236_) );
OAI21X1 OAI21X1_343 ( .A(gnd), .B(micro_ucr_hash1_a_19__3_), .C(_2236_), .Y(_2237_) );
NOR2X1 NOR2X1_219 ( .A(gnd), .B(micro_ucr_hash1_a_19__3_), .Y(_2238_) );
NAND2X1 NAND2X1_386 ( .A(micro_ucr_hash1_W_20__3_), .B(_2238_), .Y(_2239_) );
NAND3X1 NAND3X1_334 ( .A(_2226_), .B(_2237_), .C(_2239_), .Y(_2240_) );
INVX1 INVX1_249 ( .A(_2226_), .Y(_2241_) );
OAI21X1 OAI21X1_344 ( .A(gnd), .B(micro_ucr_hash1_a_19__3_), .C(micro_ucr_hash1_W_20__3_), .Y(_2242_) );
NAND2X1 NAND2X1_387 ( .A(_2236_), .B(_2238_), .Y(_2243_) );
NAND3X1 NAND3X1_335 ( .A(_2242_), .B(_2243_), .C(_2241_), .Y(_2244_) );
NAND2X1 NAND2X1_388 ( .A(_2240_), .B(_2244_), .Y(_2245_) );
XNOR2X1 XNOR2X1_160 ( .A(_2232_), .B(_2245_), .Y(micro_ucr_hash1_b_21__7_) );
INVX1 INVX1_250 ( .A(_2242_), .Y(_2246_) );
OAI21X1 OAI21X1_345 ( .A(micro_ucr_hash1_b_19__4_), .B(micro_ucr_hash1_a_19__4_), .C(micro_ucr_hash1_W_20__4_), .Y(_2247_) );
INVX1 INVX1_251 ( .A(micro_ucr_hash1_b_19__4_), .Y(_2248_) );
INVX1 INVX1_252 ( .A(micro_ucr_hash1_a_19__4_), .Y(_2249_) );
INVX1 INVX1_253 ( .A(micro_ucr_hash1_W_20__4_), .Y(_2250_) );
NAND3X1 NAND3X1_336 ( .A(_2248_), .B(_2249_), .C(_2250_), .Y(_2251_) );
AOI21X1 AOI21X1_227 ( .A(_2247_), .B(_2251_), .C(_2246_), .Y(_2157_) );
OAI21X1 OAI21X1_346 ( .A(micro_ucr_hash1_b_19__4_), .B(micro_ucr_hash1_a_19__4_), .C(_2250_), .Y(_2158_) );
NAND3X1 NAND3X1_337 ( .A(micro_ucr_hash1_W_20__4_), .B(_2248_), .C(_2249_), .Y(_2159_) );
AOI21X1 AOI21X1_228 ( .A(_2158_), .B(_2159_), .C(_2242_), .Y(_2160_) );
NOR2X1 NOR2X1_220 ( .A(_2160_), .B(_2157_), .Y(_2161_) );
AOI21X1 AOI21X1_229 ( .A(_2242_), .B(_2243_), .C(_2241_), .Y(_2162_) );
OAI21X1 OAI21X1_347 ( .A(_2162_), .B(_2231_), .C(_2244_), .Y(_2163_) );
NOR3X1 NOR3X1_63 ( .A(_2221_), .B(_2230_), .C(_2162_), .Y(_2164_) );
NOR2X1 NOR2X1_221 ( .A(_2163_), .B(_2164_), .Y(_2165_) );
XNOR2X1 XNOR2X1_161 ( .A(_2165_), .B(_2161_), .Y(micro_ucr_hash1_c_20__4_) );
NAND3X1 NAND3X1_338 ( .A(_2247_), .B(_2251_), .C(_2246_), .Y(_2166_) );
OAI21X1 OAI21X1_348 ( .A(_2165_), .B(_2157_), .C(_2166_), .Y(_2167_) );
INVX1 INVX1_254 ( .A(micro_ucr_hash1_W_20__5_), .Y(_2168_) );
OAI21X1 OAI21X1_349 ( .A(micro_ucr_hash1_b_19__5_), .B(micro_ucr_hash1_a_19__5_), .C(_2168_), .Y(_2169_) );
NOR2X1 NOR2X1_222 ( .A(micro_ucr_hash1_b_19__5_), .B(micro_ucr_hash1_a_19__5_), .Y(_2170_) );
NAND2X1 NAND2X1_389 ( .A(micro_ucr_hash1_W_20__5_), .B(_2170_), .Y(_2171_) );
NAND3X1 NAND3X1_339 ( .A(_2247_), .B(_2169_), .C(_2171_), .Y(_2172_) );
INVX1 INVX1_255 ( .A(_2247_), .Y(_2173_) );
NAND2X1 NAND2X1_390 ( .A(_2168_), .B(_2170_), .Y(_2174_) );
OAI21X1 OAI21X1_350 ( .A(micro_ucr_hash1_b_19__5_), .B(micro_ucr_hash1_a_19__5_), .C(micro_ucr_hash1_W_20__5_), .Y(_2175_) );
NAND3X1 NAND3X1_340 ( .A(_2175_), .B(_2174_), .C(_2173_), .Y(_2176_) );
NAND2X1 NAND2X1_391 ( .A(_2172_), .B(_2176_), .Y(_2177_) );
XOR2X1 XOR2X1_197 ( .A(_2167_), .B(_2177_), .Y(micro_ucr_hash1_c_20__5_) );
OAI21X1 OAI21X1_351 ( .A(gnd), .B(micro_ucr_hash1_a_19__2_), .C(_2227_), .Y(_2178_) );
NAND2X1 NAND2X1_392 ( .A(micro_ucr_hash1_W_20__2_), .B(_2228_), .Y(_2179_) );
AOI21X1 AOI21X1_230 ( .A(_2178_), .B(_2179_), .C(_2217_), .Y(_2180_) );
INVX1 INVX1_256 ( .A(_2244_), .Y(_2181_) );
AOI21X1 AOI21X1_231 ( .A(_2240_), .B(_2180_), .C(_2181_), .Y(_2182_) );
NOR3X1 NOR3X1_64 ( .A(_2222_), .B(_2223_), .C(_2224_), .Y(_2183_) );
NAND3X1 NAND3X1_341 ( .A(_2233_), .B(_2240_), .C(_2183_), .Y(_2184_) );
NAND2X1 NAND2X1_393 ( .A(_2177_), .B(_2161_), .Y(_2185_) );
AOI21X1 AOI21X1_232 ( .A(_2182_), .B(_2184_), .C(_2185_), .Y(_2186_) );
AOI22X1 AOI22X1_11 ( .A(_2174_), .B(_2175_), .C(_2166_), .D(_2247_), .Y(_2187_) );
INVX1 INVX1_257 ( .A(_2174_), .Y(_2188_) );
OAI21X1 OAI21X1_352 ( .A(micro_ucr_hash1_b_19__6_), .B(micro_ucr_hash1_a_19__6_), .C(micro_ucr_hash1_W_20__6_), .Y(_2189_) );
INVX1 INVX1_258 ( .A(micro_ucr_hash1_W_20__6_), .Y(_2190_) );
NOR2X1 NOR2X1_223 ( .A(micro_ucr_hash1_b_19__6_), .B(micro_ucr_hash1_a_19__6_), .Y(_2191_) );
NAND2X1 NAND2X1_394 ( .A(_2190_), .B(_2191_), .Y(_2192_) );
NAND2X1 NAND2X1_395 ( .A(_2189_), .B(_2192_), .Y(_2193_) );
NOR2X1 NOR2X1_224 ( .A(_2188_), .B(_2193_), .Y(_2194_) );
INVX1 INVX1_259 ( .A(_2194_), .Y(_2195_) );
NAND2X1 NAND2X1_396 ( .A(_2188_), .B(_2193_), .Y(_2196_) );
NAND2X1 NAND2X1_397 ( .A(_2196_), .B(_2195_), .Y(_2197_) );
INVX1 INVX1_260 ( .A(_2197_), .Y(_2198_) );
OAI21X1 OAI21X1_353 ( .A(_2186_), .B(_2187_), .C(_2198_), .Y(_2199_) );
NAND3X1 NAND3X1_342 ( .A(_2242_), .B(_2158_), .C(_2159_), .Y(_2200_) );
NAND2X1 NAND2X1_398 ( .A(_2200_), .B(_2166_), .Y(_2201_) );
AOI21X1 AOI21X1_233 ( .A(_2172_), .B(_2176_), .C(_2201_), .Y(_2202_) );
OAI21X1 OAI21X1_354 ( .A(_2163_), .B(_2164_), .C(_2202_), .Y(_2203_) );
INVX1 INVX1_261 ( .A(_2187_), .Y(_2204_) );
NAND3X1 NAND3X1_343 ( .A(_2204_), .B(_2197_), .C(_2203_), .Y(_2205_) );
AND2X2 AND2X2_113 ( .A(_2199_), .B(_2205_), .Y(micro_ucr_hash1_c_20__6_) );
AOI21X1 AOI21X1_234 ( .A(_2204_), .B(_2203_), .C(_2197_), .Y(_2206_) );
NOR2X1 NOR2X1_225 ( .A(micro_ucr_hash1_b_19__7_), .B(micro_ucr_hash1_a_19__7_), .Y(_2207_) );
XNOR2X1 XNOR2X1_162 ( .A(_2207_), .B(micro_ucr_hash1_W_20__7_), .Y(_2208_) );
XNOR2X1 XNOR2X1_163 ( .A(_2208_), .B(_2189_), .Y(_2209_) );
OAI21X1 OAI21X1_355 ( .A(_2206_), .B(_2194_), .C(_2209_), .Y(_2210_) );
INVX1 INVX1_262 ( .A(_2209_), .Y(_2211_) );
NAND3X1 NAND3X1_344 ( .A(_2195_), .B(_2211_), .C(_2199_), .Y(_2212_) );
NAND2X1 NAND2X1_399 ( .A(_2210_), .B(_2212_), .Y(micro_ucr_hash1_c_20__7_) );
XOR2X1 XOR2X1_198 ( .A(micro_ucr_hash1_b_21__4_), .B(gnd), .Y(micro_ucr_hash1_a_21__0_) );
XOR2X1 XOR2X1_199 ( .A(micro_ucr_hash1_b_21__5_), .B(gnd), .Y(micro_ucr_hash1_a_21__1_) );
XOR2X1 XOR2X1_200 ( .A(micro_ucr_hash1_b_21__6_), .B(gnd), .Y(micro_ucr_hash1_a_21__2_) );
XOR2X1 XOR2X1_201 ( .A(micro_ucr_hash1_b_21__7_), .B(gnd), .Y(micro_ucr_hash1_a_21__3_) );
XOR2X1 XOR2X1_202 ( .A(micro_ucr_hash1_c_20__4_), .B(micro_ucr_hash1_b_20__4_), .Y(micro_ucr_hash1_a_21__4_) );
XOR2X1 XOR2X1_203 ( .A(micro_ucr_hash1_c_20__5_), .B(micro_ucr_hash1_b_20__5_), .Y(micro_ucr_hash1_a_21__5_) );
XOR2X1 XOR2X1_204 ( .A(micro_ucr_hash1_c_20__6_), .B(micro_ucr_hash1_b_20__6_), .Y(micro_ucr_hash1_a_21__6_) );
XOR2X1 XOR2X1_205 ( .A(micro_ucr_hash1_c_20__7_), .B(micro_ucr_hash1_b_20__7_), .Y(micro_ucr_hash1_a_21__7_) );
INVX1 INVX1_263 ( .A(micro_ucr_hash1_W_21__0_), .Y(_2308_) );
NOR2X1 NOR2X1_226 ( .A(gnd), .B(micro_ucr_hash1_a_20__0_), .Y(_2309_) );
NAND2X1 NAND2X1_400 ( .A(_2308_), .B(_2309_), .Y(_2310_) );
OAI21X1 OAI21X1_356 ( .A(gnd), .B(micro_ucr_hash1_a_20__0_), .C(micro_ucr_hash1_W_21__0_), .Y(_2311_) );
NAND2X1 NAND2X1_401 ( .A(_2311_), .B(_2310_), .Y(micro_ucr_hash1_b_22__4_) );
OAI21X1 OAI21X1_357 ( .A(gnd), .B(micro_ucr_hash1_a_20__1_), .C(micro_ucr_hash1_W_21__1_), .Y(_2312_) );
INVX1 INVX1_264 ( .A(micro_ucr_hash1_W_21__1_), .Y(_2313_) );
NOR2X1 NOR2X1_227 ( .A(gnd), .B(micro_ucr_hash1_a_20__1_), .Y(_2314_) );
NAND2X1 NAND2X1_402 ( .A(_2313_), .B(_2314_), .Y(_2315_) );
NAND3X1 NAND3X1_345 ( .A(_2312_), .B(_2310_), .C(_2315_), .Y(_2316_) );
AND2X2 AND2X2_114 ( .A(_2309_), .B(_2308_), .Y(_2317_) );
INVX2 INVX2_63 ( .A(_2312_), .Y(_2318_) );
AND2X2 AND2X2_115 ( .A(_2314_), .B(_2313_), .Y(_2319_) );
OAI21X1 OAI21X1_358 ( .A(_2319_), .B(_2318_), .C(_2317_), .Y(_2320_) );
AND2X2 AND2X2_116 ( .A(_2320_), .B(_2316_), .Y(micro_ucr_hash1_b_22__5_) );
OAI21X1 OAI21X1_359 ( .A(gnd), .B(micro_ucr_hash1_a_20__2_), .C(micro_ucr_hash1_W_21__2_), .Y(_2321_) );
INVX1 INVX1_265 ( .A(micro_ucr_hash1_W_21__2_), .Y(_2322_) );
NOR2X1 NOR2X1_228 ( .A(gnd), .B(micro_ucr_hash1_a_20__2_), .Y(_2323_) );
NAND2X1 NAND2X1_403 ( .A(_2322_), .B(_2323_), .Y(_2324_) );
NAND2X1 NAND2X1_404 ( .A(_2321_), .B(_2324_), .Y(_2325_) );
NAND3X1 NAND3X1_346 ( .A(_2321_), .B(_2324_), .C(_2318_), .Y(_2326_) );
OAI21X1 OAI21X1_360 ( .A(_2316_), .B(_2325_), .C(_2326_), .Y(_2327_) );
INVX1 INVX1_266 ( .A(_2325_), .Y(_2328_) );
OAI21X1 OAI21X1_361 ( .A(_2317_), .B(_2319_), .C(_2312_), .Y(_2329_) );
NOR2X1 NOR2X1_229 ( .A(_2329_), .B(_2328_), .Y(_2330_) );
NOR2X1 NOR2X1_230 ( .A(_2327_), .B(_2330_), .Y(micro_ucr_hash1_b_22__6_) );
INVX1 INVX1_267 ( .A(micro_ucr_hash1_W_21__3_), .Y(_2331_) );
OAI21X1 OAI21X1_362 ( .A(gnd), .B(micro_ucr_hash1_a_20__3_), .C(_2331_), .Y(_2332_) );
NOR2X1 NOR2X1_231 ( .A(gnd), .B(micro_ucr_hash1_a_20__3_), .Y(_2333_) );
NAND2X1 NAND2X1_405 ( .A(micro_ucr_hash1_W_21__3_), .B(_2333_), .Y(_2334_) );
NAND3X1 NAND3X1_347 ( .A(_2321_), .B(_2332_), .C(_2334_), .Y(_2335_) );
INVX1 INVX1_268 ( .A(_2321_), .Y(_2336_) );
OAI21X1 OAI21X1_363 ( .A(gnd), .B(micro_ucr_hash1_a_20__3_), .C(micro_ucr_hash1_W_21__3_), .Y(_2337_) );
NAND2X1 NAND2X1_406 ( .A(_2331_), .B(_2333_), .Y(_2338_) );
NAND3X1 NAND3X1_348 ( .A(_2337_), .B(_2338_), .C(_2336_), .Y(_2339_) );
NAND2X1 NAND2X1_407 ( .A(_2335_), .B(_2339_), .Y(_2340_) );
XNOR2X1 XNOR2X1_164 ( .A(_2327_), .B(_2340_), .Y(micro_ucr_hash1_b_22__7_) );
INVX1 INVX1_269 ( .A(_2337_), .Y(_2341_) );
OAI21X1 OAI21X1_364 ( .A(micro_ucr_hash1_b_20__4_), .B(micro_ucr_hash1_a_20__4_), .C(micro_ucr_hash1_W_21__4_), .Y(_2342_) );
INVX1 INVX1_270 ( .A(micro_ucr_hash1_b_20__4_), .Y(_2343_) );
INVX1 INVX1_271 ( .A(micro_ucr_hash1_a_20__4_), .Y(_2344_) );
INVX1 INVX1_272 ( .A(micro_ucr_hash1_W_21__4_), .Y(_2345_) );
NAND3X1 NAND3X1_349 ( .A(_2343_), .B(_2344_), .C(_2345_), .Y(_2346_) );
AOI21X1 AOI21X1_235 ( .A(_2342_), .B(_2346_), .C(_2341_), .Y(_2252_) );
OAI21X1 OAI21X1_365 ( .A(micro_ucr_hash1_b_20__4_), .B(micro_ucr_hash1_a_20__4_), .C(_2345_), .Y(_2253_) );
NAND3X1 NAND3X1_350 ( .A(micro_ucr_hash1_W_21__4_), .B(_2343_), .C(_2344_), .Y(_2254_) );
AOI21X1 AOI21X1_236 ( .A(_2253_), .B(_2254_), .C(_2337_), .Y(_2255_) );
NOR2X1 NOR2X1_232 ( .A(_2255_), .B(_2252_), .Y(_2256_) );
AOI21X1 AOI21X1_237 ( .A(_2337_), .B(_2338_), .C(_2336_), .Y(_2257_) );
OAI21X1 OAI21X1_366 ( .A(_2257_), .B(_2326_), .C(_2339_), .Y(_2258_) );
NOR3X1 NOR3X1_65 ( .A(_2316_), .B(_2325_), .C(_2257_), .Y(_2259_) );
NOR2X1 NOR2X1_233 ( .A(_2258_), .B(_2259_), .Y(_2260_) );
XNOR2X1 XNOR2X1_165 ( .A(_2260_), .B(_2256_), .Y(micro_ucr_hash1_c_21__4_) );
NAND3X1 NAND3X1_351 ( .A(_2342_), .B(_2346_), .C(_2341_), .Y(_2261_) );
OAI21X1 OAI21X1_367 ( .A(_2260_), .B(_2252_), .C(_2261_), .Y(_2262_) );
INVX1 INVX1_273 ( .A(micro_ucr_hash1_W_21__5_), .Y(_2263_) );
OAI21X1 OAI21X1_368 ( .A(micro_ucr_hash1_b_20__5_), .B(micro_ucr_hash1_a_20__5_), .C(_2263_), .Y(_2264_) );
NOR2X1 NOR2X1_234 ( .A(micro_ucr_hash1_b_20__5_), .B(micro_ucr_hash1_a_20__5_), .Y(_2265_) );
NAND2X1 NAND2X1_408 ( .A(micro_ucr_hash1_W_21__5_), .B(_2265_), .Y(_2266_) );
NAND3X1 NAND3X1_352 ( .A(_2342_), .B(_2264_), .C(_2266_), .Y(_2267_) );
INVX1 INVX1_274 ( .A(_2342_), .Y(_2268_) );
NAND2X1 NAND2X1_409 ( .A(_2263_), .B(_2265_), .Y(_2269_) );
OAI21X1 OAI21X1_369 ( .A(micro_ucr_hash1_b_20__5_), .B(micro_ucr_hash1_a_20__5_), .C(micro_ucr_hash1_W_21__5_), .Y(_2270_) );
NAND3X1 NAND3X1_353 ( .A(_2270_), .B(_2269_), .C(_2268_), .Y(_2271_) );
NAND2X1 NAND2X1_410 ( .A(_2267_), .B(_2271_), .Y(_2272_) );
XOR2X1 XOR2X1_206 ( .A(_2262_), .B(_2272_), .Y(micro_ucr_hash1_c_21__5_) );
OAI21X1 OAI21X1_370 ( .A(gnd), .B(micro_ucr_hash1_a_20__2_), .C(_2322_), .Y(_2273_) );
NAND2X1 NAND2X1_411 ( .A(micro_ucr_hash1_W_21__2_), .B(_2323_), .Y(_2274_) );
AOI21X1 AOI21X1_238 ( .A(_2273_), .B(_2274_), .C(_2312_), .Y(_2275_) );
INVX1 INVX1_275 ( .A(_2339_), .Y(_2276_) );
AOI21X1 AOI21X1_239 ( .A(_2335_), .B(_2275_), .C(_2276_), .Y(_2277_) );
NOR3X1 NOR3X1_66 ( .A(_2317_), .B(_2318_), .C(_2319_), .Y(_2278_) );
NAND3X1 NAND3X1_354 ( .A(_2328_), .B(_2335_), .C(_2278_), .Y(_2279_) );
NAND2X1 NAND2X1_412 ( .A(_2272_), .B(_2256_), .Y(_2280_) );
AOI21X1 AOI21X1_240 ( .A(_2277_), .B(_2279_), .C(_2280_), .Y(_2281_) );
AOI22X1 AOI22X1_12 ( .A(_2269_), .B(_2270_), .C(_2261_), .D(_2342_), .Y(_2282_) );
INVX1 INVX1_276 ( .A(_2269_), .Y(_2283_) );
OAI21X1 OAI21X1_371 ( .A(micro_ucr_hash1_b_20__6_), .B(micro_ucr_hash1_a_20__6_), .C(micro_ucr_hash1_W_21__6_), .Y(_2284_) );
INVX1 INVX1_277 ( .A(micro_ucr_hash1_W_21__6_), .Y(_2285_) );
NOR2X1 NOR2X1_235 ( .A(micro_ucr_hash1_b_20__6_), .B(micro_ucr_hash1_a_20__6_), .Y(_2286_) );
NAND2X1 NAND2X1_413 ( .A(_2285_), .B(_2286_), .Y(_2287_) );
NAND2X1 NAND2X1_414 ( .A(_2284_), .B(_2287_), .Y(_2288_) );
NOR2X1 NOR2X1_236 ( .A(_2283_), .B(_2288_), .Y(_2289_) );
INVX1 INVX1_278 ( .A(_2289_), .Y(_2290_) );
NAND2X1 NAND2X1_415 ( .A(_2283_), .B(_2288_), .Y(_2291_) );
NAND2X1 NAND2X1_416 ( .A(_2291_), .B(_2290_), .Y(_2292_) );
INVX1 INVX1_279 ( .A(_2292_), .Y(_2293_) );
OAI21X1 OAI21X1_372 ( .A(_2281_), .B(_2282_), .C(_2293_), .Y(_2294_) );
NAND3X1 NAND3X1_355 ( .A(_2337_), .B(_2253_), .C(_2254_), .Y(_2295_) );
NAND2X1 NAND2X1_417 ( .A(_2295_), .B(_2261_), .Y(_2296_) );
AOI21X1 AOI21X1_241 ( .A(_2267_), .B(_2271_), .C(_2296_), .Y(_2297_) );
OAI21X1 OAI21X1_373 ( .A(_2258_), .B(_2259_), .C(_2297_), .Y(_2298_) );
INVX1 INVX1_280 ( .A(_2282_), .Y(_2299_) );
NAND3X1 NAND3X1_356 ( .A(_2299_), .B(_2292_), .C(_2298_), .Y(_2300_) );
AND2X2 AND2X2_117 ( .A(_2294_), .B(_2300_), .Y(micro_ucr_hash1_c_21__6_) );
AOI21X1 AOI21X1_242 ( .A(_2299_), .B(_2298_), .C(_2292_), .Y(_2301_) );
NOR2X1 NOR2X1_237 ( .A(micro_ucr_hash1_b_20__7_), .B(micro_ucr_hash1_a_20__7_), .Y(_2302_) );
XNOR2X1 XNOR2X1_166 ( .A(_2302_), .B(micro_ucr_hash1_W_21__7_), .Y(_2303_) );
XNOR2X1 XNOR2X1_167 ( .A(_2303_), .B(_2284_), .Y(_2304_) );
OAI21X1 OAI21X1_374 ( .A(_2301_), .B(_2289_), .C(_2304_), .Y(_2305_) );
INVX1 INVX1_281 ( .A(_2304_), .Y(_2306_) );
NAND3X1 NAND3X1_357 ( .A(_2290_), .B(_2306_), .C(_2294_), .Y(_2307_) );
NAND2X1 NAND2X1_418 ( .A(_2305_), .B(_2307_), .Y(micro_ucr_hash1_c_21__7_) );
XOR2X1 XOR2X1_207 ( .A(micro_ucr_hash1_b_22__4_), .B(gnd), .Y(micro_ucr_hash1_a_22__0_) );
XOR2X1 XOR2X1_208 ( .A(micro_ucr_hash1_b_22__5_), .B(gnd), .Y(micro_ucr_hash1_a_22__1_) );
XOR2X1 XOR2X1_209 ( .A(micro_ucr_hash1_b_22__6_), .B(gnd), .Y(micro_ucr_hash1_a_22__2_) );
XOR2X1 XOR2X1_210 ( .A(micro_ucr_hash1_b_22__7_), .B(gnd), .Y(micro_ucr_hash1_a_22__3_) );
XOR2X1 XOR2X1_211 ( .A(micro_ucr_hash1_c_21__4_), .B(micro_ucr_hash1_b_21__4_), .Y(micro_ucr_hash1_a_22__4_) );
XOR2X1 XOR2X1_212 ( .A(micro_ucr_hash1_c_21__5_), .B(micro_ucr_hash1_b_21__5_), .Y(micro_ucr_hash1_a_22__5_) );
XOR2X1 XOR2X1_213 ( .A(micro_ucr_hash1_c_21__6_), .B(micro_ucr_hash1_b_21__6_), .Y(micro_ucr_hash1_a_22__6_) );
XOR2X1 XOR2X1_214 ( .A(micro_ucr_hash1_c_21__7_), .B(micro_ucr_hash1_b_21__7_), .Y(micro_ucr_hash1_a_22__7_) );
INVX1 INVX1_282 ( .A(micro_ucr_hash1_W_22__0_), .Y(_2403_) );
NOR2X1 NOR2X1_238 ( .A(gnd), .B(micro_ucr_hash1_a_21__0_), .Y(_2404_) );
NAND2X1 NAND2X1_419 ( .A(_2403_), .B(_2404_), .Y(_2405_) );
OAI21X1 OAI21X1_375 ( .A(gnd), .B(micro_ucr_hash1_a_21__0_), .C(micro_ucr_hash1_W_22__0_), .Y(_2406_) );
NAND2X1 NAND2X1_420 ( .A(_2406_), .B(_2405_), .Y(micro_ucr_hash1_b_23__4_) );
OAI21X1 OAI21X1_376 ( .A(gnd), .B(micro_ucr_hash1_a_21__1_), .C(micro_ucr_hash1_W_22__1_), .Y(_2407_) );
INVX1 INVX1_283 ( .A(micro_ucr_hash1_W_22__1_), .Y(_2408_) );
NOR2X1 NOR2X1_239 ( .A(gnd), .B(micro_ucr_hash1_a_21__1_), .Y(_2409_) );
NAND2X1 NAND2X1_421 ( .A(_2408_), .B(_2409_), .Y(_2410_) );
NAND3X1 NAND3X1_358 ( .A(_2407_), .B(_2405_), .C(_2410_), .Y(_2411_) );
AND2X2 AND2X2_118 ( .A(_2404_), .B(_2403_), .Y(_2412_) );
INVX2 INVX2_64 ( .A(_2407_), .Y(_2413_) );
AND2X2 AND2X2_119 ( .A(_2409_), .B(_2408_), .Y(_2414_) );
OAI21X1 OAI21X1_377 ( .A(_2414_), .B(_2413_), .C(_2412_), .Y(_2415_) );
AND2X2 AND2X2_120 ( .A(_2415_), .B(_2411_), .Y(micro_ucr_hash1_b_23__5_) );
OAI21X1 OAI21X1_378 ( .A(gnd), .B(micro_ucr_hash1_a_21__2_), .C(micro_ucr_hash1_W_22__2_), .Y(_2416_) );
INVX1 INVX1_284 ( .A(micro_ucr_hash1_W_22__2_), .Y(_2417_) );
NOR2X1 NOR2X1_240 ( .A(gnd), .B(micro_ucr_hash1_a_21__2_), .Y(_2418_) );
NAND2X1 NAND2X1_422 ( .A(_2417_), .B(_2418_), .Y(_2419_) );
NAND2X1 NAND2X1_423 ( .A(_2416_), .B(_2419_), .Y(_2420_) );
NAND3X1 NAND3X1_359 ( .A(_2416_), .B(_2419_), .C(_2413_), .Y(_2421_) );
OAI21X1 OAI21X1_379 ( .A(_2411_), .B(_2420_), .C(_2421_), .Y(_2422_) );
INVX1 INVX1_285 ( .A(_2420_), .Y(_2423_) );
OAI21X1 OAI21X1_380 ( .A(_2412_), .B(_2414_), .C(_2407_), .Y(_2424_) );
NOR2X1 NOR2X1_241 ( .A(_2424_), .B(_2423_), .Y(_2425_) );
NOR2X1 NOR2X1_242 ( .A(_2422_), .B(_2425_), .Y(micro_ucr_hash1_b_23__6_) );
INVX1 INVX1_286 ( .A(micro_ucr_hash1_W_22__3_), .Y(_2426_) );
OAI21X1 OAI21X1_381 ( .A(gnd), .B(micro_ucr_hash1_a_21__3_), .C(_2426_), .Y(_2427_) );
NOR2X1 NOR2X1_243 ( .A(gnd), .B(micro_ucr_hash1_a_21__3_), .Y(_2428_) );
NAND2X1 NAND2X1_424 ( .A(micro_ucr_hash1_W_22__3_), .B(_2428_), .Y(_2429_) );
NAND3X1 NAND3X1_360 ( .A(_2416_), .B(_2427_), .C(_2429_), .Y(_2430_) );
INVX1 INVX1_287 ( .A(_2416_), .Y(_2431_) );
OAI21X1 OAI21X1_382 ( .A(gnd), .B(micro_ucr_hash1_a_21__3_), .C(micro_ucr_hash1_W_22__3_), .Y(_2432_) );
NAND2X1 NAND2X1_425 ( .A(_2426_), .B(_2428_), .Y(_2433_) );
NAND3X1 NAND3X1_361 ( .A(_2432_), .B(_2433_), .C(_2431_), .Y(_2434_) );
NAND2X1 NAND2X1_426 ( .A(_2430_), .B(_2434_), .Y(_2435_) );
XNOR2X1 XNOR2X1_168 ( .A(_2422_), .B(_2435_), .Y(micro_ucr_hash1_b_23__7_) );
INVX1 INVX1_288 ( .A(_2432_), .Y(_2436_) );
OAI21X1 OAI21X1_383 ( .A(micro_ucr_hash1_b_21__4_), .B(micro_ucr_hash1_a_21__4_), .C(micro_ucr_hash1_W_22__4_), .Y(_2437_) );
INVX1 INVX1_289 ( .A(micro_ucr_hash1_b_21__4_), .Y(_2438_) );
INVX1 INVX1_290 ( .A(micro_ucr_hash1_a_21__4_), .Y(_2439_) );
INVX1 INVX1_291 ( .A(micro_ucr_hash1_W_22__4_), .Y(_2440_) );
NAND3X1 NAND3X1_362 ( .A(_2438_), .B(_2439_), .C(_2440_), .Y(_2441_) );
AOI21X1 AOI21X1_243 ( .A(_2437_), .B(_2441_), .C(_2436_), .Y(_2347_) );
OAI21X1 OAI21X1_384 ( .A(micro_ucr_hash1_b_21__4_), .B(micro_ucr_hash1_a_21__4_), .C(_2440_), .Y(_2348_) );
NAND3X1 NAND3X1_363 ( .A(micro_ucr_hash1_W_22__4_), .B(_2438_), .C(_2439_), .Y(_2349_) );
AOI21X1 AOI21X1_244 ( .A(_2348_), .B(_2349_), .C(_2432_), .Y(_2350_) );
NOR2X1 NOR2X1_244 ( .A(_2350_), .B(_2347_), .Y(_2351_) );
AOI21X1 AOI21X1_245 ( .A(_2432_), .B(_2433_), .C(_2431_), .Y(_2352_) );
OAI21X1 OAI21X1_385 ( .A(_2352_), .B(_2421_), .C(_2434_), .Y(_2353_) );
NOR3X1 NOR3X1_67 ( .A(_2411_), .B(_2420_), .C(_2352_), .Y(_2354_) );
NOR2X1 NOR2X1_245 ( .A(_2353_), .B(_2354_), .Y(_2355_) );
XNOR2X1 XNOR2X1_169 ( .A(_2355_), .B(_2351_), .Y(micro_ucr_hash1_c_22__4_) );
NAND3X1 NAND3X1_364 ( .A(_2437_), .B(_2441_), .C(_2436_), .Y(_2356_) );
OAI21X1 OAI21X1_386 ( .A(_2355_), .B(_2347_), .C(_2356_), .Y(_2357_) );
INVX1 INVX1_292 ( .A(micro_ucr_hash1_W_22__5_), .Y(_2358_) );
OAI21X1 OAI21X1_387 ( .A(micro_ucr_hash1_b_21__5_), .B(micro_ucr_hash1_a_21__5_), .C(_2358_), .Y(_2359_) );
NOR2X1 NOR2X1_246 ( .A(micro_ucr_hash1_b_21__5_), .B(micro_ucr_hash1_a_21__5_), .Y(_2360_) );
NAND2X1 NAND2X1_427 ( .A(micro_ucr_hash1_W_22__5_), .B(_2360_), .Y(_2361_) );
NAND3X1 NAND3X1_365 ( .A(_2437_), .B(_2359_), .C(_2361_), .Y(_2362_) );
INVX1 INVX1_293 ( .A(_2437_), .Y(_2363_) );
NAND2X1 NAND2X1_428 ( .A(_2358_), .B(_2360_), .Y(_2364_) );
OAI21X1 OAI21X1_388 ( .A(micro_ucr_hash1_b_21__5_), .B(micro_ucr_hash1_a_21__5_), .C(micro_ucr_hash1_W_22__5_), .Y(_2365_) );
NAND3X1 NAND3X1_366 ( .A(_2365_), .B(_2364_), .C(_2363_), .Y(_2366_) );
NAND2X1 NAND2X1_429 ( .A(_2362_), .B(_2366_), .Y(_2367_) );
XOR2X1 XOR2X1_215 ( .A(_2357_), .B(_2367_), .Y(micro_ucr_hash1_c_22__5_) );
OAI21X1 OAI21X1_389 ( .A(gnd), .B(micro_ucr_hash1_a_21__2_), .C(_2417_), .Y(_2368_) );
NAND2X1 NAND2X1_430 ( .A(micro_ucr_hash1_W_22__2_), .B(_2418_), .Y(_2369_) );
AOI21X1 AOI21X1_246 ( .A(_2368_), .B(_2369_), .C(_2407_), .Y(_2370_) );
INVX1 INVX1_294 ( .A(_2434_), .Y(_2371_) );
AOI21X1 AOI21X1_247 ( .A(_2430_), .B(_2370_), .C(_2371_), .Y(_2372_) );
NOR3X1 NOR3X1_68 ( .A(_2412_), .B(_2413_), .C(_2414_), .Y(_2373_) );
NAND3X1 NAND3X1_367 ( .A(_2423_), .B(_2430_), .C(_2373_), .Y(_2374_) );
NAND2X1 NAND2X1_431 ( .A(_2367_), .B(_2351_), .Y(_2375_) );
AOI21X1 AOI21X1_248 ( .A(_2372_), .B(_2374_), .C(_2375_), .Y(_2376_) );
AOI22X1 AOI22X1_13 ( .A(_2364_), .B(_2365_), .C(_2356_), .D(_2437_), .Y(_2377_) );
INVX1 INVX1_295 ( .A(_2364_), .Y(_2378_) );
OAI21X1 OAI21X1_390 ( .A(micro_ucr_hash1_b_21__6_), .B(micro_ucr_hash1_a_21__6_), .C(micro_ucr_hash1_W_22__6_), .Y(_2379_) );
INVX1 INVX1_296 ( .A(micro_ucr_hash1_W_22__6_), .Y(_2380_) );
NOR2X1 NOR2X1_247 ( .A(micro_ucr_hash1_b_21__6_), .B(micro_ucr_hash1_a_21__6_), .Y(_2381_) );
NAND2X1 NAND2X1_432 ( .A(_2380_), .B(_2381_), .Y(_2382_) );
NAND2X1 NAND2X1_433 ( .A(_2379_), .B(_2382_), .Y(_2383_) );
NOR2X1 NOR2X1_248 ( .A(_2378_), .B(_2383_), .Y(_2384_) );
INVX1 INVX1_297 ( .A(_2384_), .Y(_2385_) );
NAND2X1 NAND2X1_434 ( .A(_2378_), .B(_2383_), .Y(_2386_) );
NAND2X1 NAND2X1_435 ( .A(_2386_), .B(_2385_), .Y(_2387_) );
INVX1 INVX1_298 ( .A(_2387_), .Y(_2388_) );
OAI21X1 OAI21X1_391 ( .A(_2376_), .B(_2377_), .C(_2388_), .Y(_2389_) );
NAND3X1 NAND3X1_368 ( .A(_2432_), .B(_2348_), .C(_2349_), .Y(_2390_) );
NAND2X1 NAND2X1_436 ( .A(_2390_), .B(_2356_), .Y(_2391_) );
AOI21X1 AOI21X1_249 ( .A(_2362_), .B(_2366_), .C(_2391_), .Y(_2392_) );
OAI21X1 OAI21X1_392 ( .A(_2353_), .B(_2354_), .C(_2392_), .Y(_2393_) );
INVX1 INVX1_299 ( .A(_2377_), .Y(_2394_) );
NAND3X1 NAND3X1_369 ( .A(_2394_), .B(_2387_), .C(_2393_), .Y(_2395_) );
AND2X2 AND2X2_121 ( .A(_2389_), .B(_2395_), .Y(micro_ucr_hash1_c_22__6_) );
AOI21X1 AOI21X1_250 ( .A(_2394_), .B(_2393_), .C(_2387_), .Y(_2396_) );
NOR2X1 NOR2X1_249 ( .A(micro_ucr_hash1_b_21__7_), .B(micro_ucr_hash1_a_21__7_), .Y(_2397_) );
XNOR2X1 XNOR2X1_170 ( .A(_2397_), .B(micro_ucr_hash1_W_22__7_), .Y(_2398_) );
XNOR2X1 XNOR2X1_171 ( .A(_2398_), .B(_2379_), .Y(_2399_) );
OAI21X1 OAI21X1_393 ( .A(_2396_), .B(_2384_), .C(_2399_), .Y(_2400_) );
INVX1 INVX1_300 ( .A(_2399_), .Y(_2401_) );
NAND3X1 NAND3X1_370 ( .A(_2385_), .B(_2401_), .C(_2389_), .Y(_2402_) );
NAND2X1 NAND2X1_437 ( .A(_2400_), .B(_2402_), .Y(micro_ucr_hash1_c_22__7_) );
XOR2X1 XOR2X1_216 ( .A(micro_ucr_hash1_b_23__4_), .B(gnd), .Y(micro_ucr_hash1_a_23__0_) );
XOR2X1 XOR2X1_217 ( .A(micro_ucr_hash1_b_23__5_), .B(gnd), .Y(micro_ucr_hash1_a_23__1_) );
XOR2X1 XOR2X1_218 ( .A(micro_ucr_hash1_b_23__6_), .B(gnd), .Y(micro_ucr_hash1_a_23__2_) );
XOR2X1 XOR2X1_219 ( .A(micro_ucr_hash1_b_23__7_), .B(gnd), .Y(micro_ucr_hash1_a_23__3_) );
XOR2X1 XOR2X1_220 ( .A(micro_ucr_hash1_c_22__4_), .B(micro_ucr_hash1_b_22__4_), .Y(micro_ucr_hash1_a_23__4_) );
XOR2X1 XOR2X1_221 ( .A(micro_ucr_hash1_c_22__5_), .B(micro_ucr_hash1_b_22__5_), .Y(micro_ucr_hash1_a_23__5_) );
XOR2X1 XOR2X1_222 ( .A(micro_ucr_hash1_c_22__6_), .B(micro_ucr_hash1_b_22__6_), .Y(micro_ucr_hash1_a_23__6_) );
XOR2X1 XOR2X1_223 ( .A(micro_ucr_hash1_c_22__7_), .B(micro_ucr_hash1_b_22__7_), .Y(micro_ucr_hash1_a_23__7_) );
INVX1 INVX1_301 ( .A(micro_ucr_hash1_W_23__0_), .Y(_2498_) );
NOR2X1 NOR2X1_250 ( .A(gnd), .B(micro_ucr_hash1_a_22__0_), .Y(_2499_) );
NAND2X1 NAND2X1_438 ( .A(_2498_), .B(_2499_), .Y(_2500_) );
OAI21X1 OAI21X1_394 ( .A(gnd), .B(micro_ucr_hash1_a_22__0_), .C(micro_ucr_hash1_W_23__0_), .Y(_2501_) );
NAND2X1 NAND2X1_439 ( .A(_2501_), .B(_2500_), .Y(micro_ucr_hash1_b_24__4_) );
OAI21X1 OAI21X1_395 ( .A(gnd), .B(micro_ucr_hash1_a_22__1_), .C(micro_ucr_hash1_W_23__1_), .Y(_2502_) );
INVX1 INVX1_302 ( .A(micro_ucr_hash1_W_23__1_), .Y(_2503_) );
NOR2X1 NOR2X1_251 ( .A(gnd), .B(micro_ucr_hash1_a_22__1_), .Y(_2504_) );
NAND2X1 NAND2X1_440 ( .A(_2503_), .B(_2504_), .Y(_2505_) );
NAND3X1 NAND3X1_371 ( .A(_2502_), .B(_2500_), .C(_2505_), .Y(_2506_) );
AND2X2 AND2X2_122 ( .A(_2499_), .B(_2498_), .Y(_2507_) );
INVX2 INVX2_65 ( .A(_2502_), .Y(_2508_) );
AND2X2 AND2X2_123 ( .A(_2504_), .B(_2503_), .Y(_2509_) );
OAI21X1 OAI21X1_396 ( .A(_2509_), .B(_2508_), .C(_2507_), .Y(_2510_) );
AND2X2 AND2X2_124 ( .A(_2510_), .B(_2506_), .Y(micro_ucr_hash1_b_24__5_) );
OAI21X1 OAI21X1_397 ( .A(gnd), .B(micro_ucr_hash1_a_22__2_), .C(micro_ucr_hash1_W_23__2_), .Y(_2511_) );
INVX1 INVX1_303 ( .A(micro_ucr_hash1_W_23__2_), .Y(_2512_) );
NOR2X1 NOR2X1_252 ( .A(gnd), .B(micro_ucr_hash1_a_22__2_), .Y(_2513_) );
NAND2X1 NAND2X1_441 ( .A(_2512_), .B(_2513_), .Y(_2514_) );
NAND2X1 NAND2X1_442 ( .A(_2511_), .B(_2514_), .Y(_2515_) );
NAND3X1 NAND3X1_372 ( .A(_2511_), .B(_2514_), .C(_2508_), .Y(_2516_) );
OAI21X1 OAI21X1_398 ( .A(_2506_), .B(_2515_), .C(_2516_), .Y(_2517_) );
INVX1 INVX1_304 ( .A(_2515_), .Y(_2518_) );
OAI21X1 OAI21X1_399 ( .A(_2507_), .B(_2509_), .C(_2502_), .Y(_2519_) );
NOR2X1 NOR2X1_253 ( .A(_2519_), .B(_2518_), .Y(_2520_) );
NOR2X1 NOR2X1_254 ( .A(_2517_), .B(_2520_), .Y(micro_ucr_hash1_b_24__6_) );
INVX1 INVX1_305 ( .A(micro_ucr_hash1_W_23__3_), .Y(_2521_) );
OAI21X1 OAI21X1_400 ( .A(gnd), .B(micro_ucr_hash1_a_22__3_), .C(_2521_), .Y(_2522_) );
NOR2X1 NOR2X1_255 ( .A(gnd), .B(micro_ucr_hash1_a_22__3_), .Y(_2523_) );
NAND2X1 NAND2X1_443 ( .A(micro_ucr_hash1_W_23__3_), .B(_2523_), .Y(_2524_) );
NAND3X1 NAND3X1_373 ( .A(_2511_), .B(_2522_), .C(_2524_), .Y(_2525_) );
INVX1 INVX1_306 ( .A(_2511_), .Y(_2526_) );
OAI21X1 OAI21X1_401 ( .A(gnd), .B(micro_ucr_hash1_a_22__3_), .C(micro_ucr_hash1_W_23__3_), .Y(_2527_) );
NAND2X1 NAND2X1_444 ( .A(_2521_), .B(_2523_), .Y(_2528_) );
NAND3X1 NAND3X1_374 ( .A(_2527_), .B(_2528_), .C(_2526_), .Y(_2529_) );
NAND2X1 NAND2X1_445 ( .A(_2525_), .B(_2529_), .Y(_2530_) );
XNOR2X1 XNOR2X1_172 ( .A(_2517_), .B(_2530_), .Y(micro_ucr_hash1_b_24__7_) );
INVX1 INVX1_307 ( .A(_2527_), .Y(_2531_) );
OAI21X1 OAI21X1_402 ( .A(micro_ucr_hash1_b_22__4_), .B(micro_ucr_hash1_a_22__4_), .C(micro_ucr_hash1_W_23__4_), .Y(_2532_) );
INVX1 INVX1_308 ( .A(micro_ucr_hash1_b_22__4_), .Y(_2533_) );
INVX1 INVX1_309 ( .A(micro_ucr_hash1_a_22__4_), .Y(_2534_) );
INVX1 INVX1_310 ( .A(micro_ucr_hash1_W_23__4_), .Y(_2535_) );
NAND3X1 NAND3X1_375 ( .A(_2533_), .B(_2534_), .C(_2535_), .Y(_2536_) );
AOI21X1 AOI21X1_251 ( .A(_2532_), .B(_2536_), .C(_2531_), .Y(_2442_) );
OAI21X1 OAI21X1_403 ( .A(micro_ucr_hash1_b_22__4_), .B(micro_ucr_hash1_a_22__4_), .C(_2535_), .Y(_2443_) );
NAND3X1 NAND3X1_376 ( .A(micro_ucr_hash1_W_23__4_), .B(_2533_), .C(_2534_), .Y(_2444_) );
AOI21X1 AOI21X1_252 ( .A(_2443_), .B(_2444_), .C(_2527_), .Y(_2445_) );
NOR2X1 NOR2X1_256 ( .A(_2445_), .B(_2442_), .Y(_2446_) );
AOI21X1 AOI21X1_253 ( .A(_2527_), .B(_2528_), .C(_2526_), .Y(_2447_) );
OAI21X1 OAI21X1_404 ( .A(_2447_), .B(_2516_), .C(_2529_), .Y(_2448_) );
NOR3X1 NOR3X1_69 ( .A(_2506_), .B(_2515_), .C(_2447_), .Y(_2449_) );
NOR2X1 NOR2X1_257 ( .A(_2448_), .B(_2449_), .Y(_2450_) );
XNOR2X1 XNOR2X1_173 ( .A(_2450_), .B(_2446_), .Y(micro_ucr_hash1_c_23__4_) );
NAND3X1 NAND3X1_377 ( .A(_2532_), .B(_2536_), .C(_2531_), .Y(_2451_) );
OAI21X1 OAI21X1_405 ( .A(_2450_), .B(_2442_), .C(_2451_), .Y(_2452_) );
INVX1 INVX1_311 ( .A(micro_ucr_hash1_W_23__5_), .Y(_2453_) );
OAI21X1 OAI21X1_406 ( .A(micro_ucr_hash1_b_22__5_), .B(micro_ucr_hash1_a_22__5_), .C(_2453_), .Y(_2454_) );
NOR2X1 NOR2X1_258 ( .A(micro_ucr_hash1_b_22__5_), .B(micro_ucr_hash1_a_22__5_), .Y(_2455_) );
NAND2X1 NAND2X1_446 ( .A(micro_ucr_hash1_W_23__5_), .B(_2455_), .Y(_2456_) );
NAND3X1 NAND3X1_378 ( .A(_2532_), .B(_2454_), .C(_2456_), .Y(_2457_) );
INVX1 INVX1_312 ( .A(_2532_), .Y(_2458_) );
NAND2X1 NAND2X1_447 ( .A(_2453_), .B(_2455_), .Y(_2459_) );
OAI21X1 OAI21X1_407 ( .A(micro_ucr_hash1_b_22__5_), .B(micro_ucr_hash1_a_22__5_), .C(micro_ucr_hash1_W_23__5_), .Y(_2460_) );
NAND3X1 NAND3X1_379 ( .A(_2460_), .B(_2459_), .C(_2458_), .Y(_2461_) );
NAND2X1 NAND2X1_448 ( .A(_2457_), .B(_2461_), .Y(_2462_) );
XOR2X1 XOR2X1_224 ( .A(_2452_), .B(_2462_), .Y(micro_ucr_hash1_c_23__5_) );
OAI21X1 OAI21X1_408 ( .A(gnd), .B(micro_ucr_hash1_a_22__2_), .C(_2512_), .Y(_2463_) );
NAND2X1 NAND2X1_449 ( .A(micro_ucr_hash1_W_23__2_), .B(_2513_), .Y(_2464_) );
AOI21X1 AOI21X1_254 ( .A(_2463_), .B(_2464_), .C(_2502_), .Y(_2465_) );
INVX1 INVX1_313 ( .A(_2529_), .Y(_2466_) );
AOI21X1 AOI21X1_255 ( .A(_2525_), .B(_2465_), .C(_2466_), .Y(_2467_) );
NOR3X1 NOR3X1_70 ( .A(_2507_), .B(_2508_), .C(_2509_), .Y(_2468_) );
NAND3X1 NAND3X1_380 ( .A(_2518_), .B(_2525_), .C(_2468_), .Y(_2469_) );
NAND2X1 NAND2X1_450 ( .A(_2462_), .B(_2446_), .Y(_2470_) );
AOI21X1 AOI21X1_256 ( .A(_2467_), .B(_2469_), .C(_2470_), .Y(_2471_) );
AOI22X1 AOI22X1_14 ( .A(_2459_), .B(_2460_), .C(_2451_), .D(_2532_), .Y(_2472_) );
INVX1 INVX1_314 ( .A(_2459_), .Y(_2473_) );
OAI21X1 OAI21X1_409 ( .A(micro_ucr_hash1_b_22__6_), .B(micro_ucr_hash1_a_22__6_), .C(micro_ucr_hash1_W_23__6_), .Y(_2474_) );
INVX1 INVX1_315 ( .A(micro_ucr_hash1_W_23__6_), .Y(_2475_) );
NOR2X1 NOR2X1_259 ( .A(micro_ucr_hash1_b_22__6_), .B(micro_ucr_hash1_a_22__6_), .Y(_2476_) );
NAND2X1 NAND2X1_451 ( .A(_2475_), .B(_2476_), .Y(_2477_) );
NAND2X1 NAND2X1_452 ( .A(_2474_), .B(_2477_), .Y(_2478_) );
NOR2X1 NOR2X1_260 ( .A(_2473_), .B(_2478_), .Y(_2479_) );
INVX1 INVX1_316 ( .A(_2479_), .Y(_2480_) );
NAND2X1 NAND2X1_453 ( .A(_2473_), .B(_2478_), .Y(_2481_) );
NAND2X1 NAND2X1_454 ( .A(_2481_), .B(_2480_), .Y(_2482_) );
INVX1 INVX1_317 ( .A(_2482_), .Y(_2483_) );
OAI21X1 OAI21X1_410 ( .A(_2471_), .B(_2472_), .C(_2483_), .Y(_2484_) );
NAND3X1 NAND3X1_381 ( .A(_2527_), .B(_2443_), .C(_2444_), .Y(_2485_) );
NAND2X1 NAND2X1_455 ( .A(_2485_), .B(_2451_), .Y(_2486_) );
AOI21X1 AOI21X1_257 ( .A(_2457_), .B(_2461_), .C(_2486_), .Y(_2487_) );
OAI21X1 OAI21X1_411 ( .A(_2448_), .B(_2449_), .C(_2487_), .Y(_2488_) );
INVX1 INVX1_318 ( .A(_2472_), .Y(_2489_) );
NAND3X1 NAND3X1_382 ( .A(_2489_), .B(_2482_), .C(_2488_), .Y(_2490_) );
AND2X2 AND2X2_125 ( .A(_2484_), .B(_2490_), .Y(micro_ucr_hash1_c_23__6_) );
AOI21X1 AOI21X1_258 ( .A(_2489_), .B(_2488_), .C(_2482_), .Y(_2491_) );
NOR2X1 NOR2X1_261 ( .A(micro_ucr_hash1_b_22__7_), .B(micro_ucr_hash1_a_22__7_), .Y(_2492_) );
XNOR2X1 XNOR2X1_174 ( .A(_2492_), .B(micro_ucr_hash1_W_23__7_), .Y(_2493_) );
XNOR2X1 XNOR2X1_175 ( .A(_2493_), .B(_2474_), .Y(_2494_) );
OAI21X1 OAI21X1_412 ( .A(_2491_), .B(_2479_), .C(_2494_), .Y(_2495_) );
INVX1 INVX1_319 ( .A(_2494_), .Y(_2496_) );
NAND3X1 NAND3X1_383 ( .A(_2480_), .B(_2496_), .C(_2484_), .Y(_2497_) );
NAND2X1 NAND2X1_456 ( .A(_2495_), .B(_2497_), .Y(micro_ucr_hash1_c_23__7_) );
XOR2X1 XOR2X1_225 ( .A(micro_ucr_hash1_b_24__4_), .B(gnd), .Y(micro_ucr_hash1_a_24__0_) );
XOR2X1 XOR2X1_226 ( .A(micro_ucr_hash1_b_24__5_), .B(gnd), .Y(micro_ucr_hash1_a_24__1_) );
XOR2X1 XOR2X1_227 ( .A(micro_ucr_hash1_b_24__6_), .B(gnd), .Y(micro_ucr_hash1_a_24__2_) );
XOR2X1 XOR2X1_228 ( .A(micro_ucr_hash1_b_24__7_), .B(gnd), .Y(micro_ucr_hash1_a_24__3_) );
XOR2X1 XOR2X1_229 ( .A(micro_ucr_hash1_c_23__4_), .B(micro_ucr_hash1_b_23__4_), .Y(micro_ucr_hash1_a_24__4_) );
XOR2X1 XOR2X1_230 ( .A(micro_ucr_hash1_c_23__5_), .B(micro_ucr_hash1_b_23__5_), .Y(micro_ucr_hash1_a_24__5_) );
XOR2X1 XOR2X1_231 ( .A(micro_ucr_hash1_c_23__6_), .B(micro_ucr_hash1_b_23__6_), .Y(micro_ucr_hash1_a_24__6_) );
XOR2X1 XOR2X1_232 ( .A(micro_ucr_hash1_c_23__7_), .B(micro_ucr_hash1_b_23__7_), .Y(micro_ucr_hash1_a_24__7_) );
INVX1 INVX1_320 ( .A(micro_ucr_hash1_W_24__0_), .Y(_2593_) );
NOR2X1 NOR2X1_262 ( .A(gnd), .B(micro_ucr_hash1_a_23__0_), .Y(_2594_) );
NAND2X1 NAND2X1_457 ( .A(_2593_), .B(_2594_), .Y(_2595_) );
OAI21X1 OAI21X1_413 ( .A(gnd), .B(micro_ucr_hash1_a_23__0_), .C(micro_ucr_hash1_W_24__0_), .Y(_2596_) );
NAND2X1 NAND2X1_458 ( .A(_2596_), .B(_2595_), .Y(micro_ucr_hash1_b_25__4_) );
OAI21X1 OAI21X1_414 ( .A(gnd), .B(micro_ucr_hash1_a_23__1_), .C(micro_ucr_hash1_W_24__1_), .Y(_2597_) );
INVX1 INVX1_321 ( .A(micro_ucr_hash1_W_24__1_), .Y(_2598_) );
NOR2X1 NOR2X1_263 ( .A(gnd), .B(micro_ucr_hash1_a_23__1_), .Y(_2599_) );
NAND2X1 NAND2X1_459 ( .A(_2598_), .B(_2599_), .Y(_2600_) );
NAND3X1 NAND3X1_384 ( .A(_2597_), .B(_2595_), .C(_2600_), .Y(_2601_) );
AND2X2 AND2X2_126 ( .A(_2594_), .B(_2593_), .Y(_2602_) );
INVX2 INVX2_66 ( .A(_2597_), .Y(_2603_) );
AND2X2 AND2X2_127 ( .A(_2599_), .B(_2598_), .Y(_2604_) );
OAI21X1 OAI21X1_415 ( .A(_2604_), .B(_2603_), .C(_2602_), .Y(_2605_) );
AND2X2 AND2X2_128 ( .A(_2605_), .B(_2601_), .Y(micro_ucr_hash1_b_25__5_) );
OAI21X1 OAI21X1_416 ( .A(gnd), .B(micro_ucr_hash1_a_23__2_), .C(micro_ucr_hash1_W_24__2_), .Y(_2606_) );
INVX1 INVX1_322 ( .A(micro_ucr_hash1_W_24__2_), .Y(_2607_) );
NOR2X1 NOR2X1_264 ( .A(gnd), .B(micro_ucr_hash1_a_23__2_), .Y(_2608_) );
NAND2X1 NAND2X1_460 ( .A(_2607_), .B(_2608_), .Y(_2609_) );
NAND2X1 NAND2X1_461 ( .A(_2606_), .B(_2609_), .Y(_2610_) );
NAND3X1 NAND3X1_385 ( .A(_2606_), .B(_2609_), .C(_2603_), .Y(_2611_) );
OAI21X1 OAI21X1_417 ( .A(_2601_), .B(_2610_), .C(_2611_), .Y(_2612_) );
INVX1 INVX1_323 ( .A(_2610_), .Y(_2613_) );
OAI21X1 OAI21X1_418 ( .A(_2602_), .B(_2604_), .C(_2597_), .Y(_2614_) );
NOR2X1 NOR2X1_265 ( .A(_2614_), .B(_2613_), .Y(_2615_) );
NOR2X1 NOR2X1_266 ( .A(_2612_), .B(_2615_), .Y(micro_ucr_hash1_b_25__6_) );
INVX1 INVX1_324 ( .A(micro_ucr_hash1_W_24__3_), .Y(_2616_) );
OAI21X1 OAI21X1_419 ( .A(gnd), .B(micro_ucr_hash1_a_23__3_), .C(_2616_), .Y(_2617_) );
NOR2X1 NOR2X1_267 ( .A(gnd), .B(micro_ucr_hash1_a_23__3_), .Y(_2618_) );
NAND2X1 NAND2X1_462 ( .A(micro_ucr_hash1_W_24__3_), .B(_2618_), .Y(_2619_) );
NAND3X1 NAND3X1_386 ( .A(_2606_), .B(_2617_), .C(_2619_), .Y(_2620_) );
INVX1 INVX1_325 ( .A(_2606_), .Y(_2621_) );
OAI21X1 OAI21X1_420 ( .A(gnd), .B(micro_ucr_hash1_a_23__3_), .C(micro_ucr_hash1_W_24__3_), .Y(_2622_) );
NAND2X1 NAND2X1_463 ( .A(_2616_), .B(_2618_), .Y(_2623_) );
NAND3X1 NAND3X1_387 ( .A(_2622_), .B(_2623_), .C(_2621_), .Y(_2624_) );
NAND2X1 NAND2X1_464 ( .A(_2620_), .B(_2624_), .Y(_2625_) );
XNOR2X1 XNOR2X1_176 ( .A(_2612_), .B(_2625_), .Y(micro_ucr_hash1_b_25__7_) );
INVX1 INVX1_326 ( .A(_2622_), .Y(_2626_) );
OAI21X1 OAI21X1_421 ( .A(micro_ucr_hash1_b_23__4_), .B(micro_ucr_hash1_a_23__4_), .C(micro_ucr_hash1_W_24__4_), .Y(_2627_) );
INVX1 INVX1_327 ( .A(micro_ucr_hash1_b_23__4_), .Y(_2628_) );
INVX1 INVX1_328 ( .A(micro_ucr_hash1_a_23__4_), .Y(_2629_) );
INVX1 INVX1_329 ( .A(micro_ucr_hash1_W_24__4_), .Y(_2630_) );
NAND3X1 NAND3X1_388 ( .A(_2628_), .B(_2629_), .C(_2630_), .Y(_2631_) );
AOI21X1 AOI21X1_259 ( .A(_2627_), .B(_2631_), .C(_2626_), .Y(_2537_) );
OAI21X1 OAI21X1_422 ( .A(micro_ucr_hash1_b_23__4_), .B(micro_ucr_hash1_a_23__4_), .C(_2630_), .Y(_2538_) );
NAND3X1 NAND3X1_389 ( .A(micro_ucr_hash1_W_24__4_), .B(_2628_), .C(_2629_), .Y(_2539_) );
AOI21X1 AOI21X1_260 ( .A(_2538_), .B(_2539_), .C(_2622_), .Y(_2540_) );
NOR2X1 NOR2X1_268 ( .A(_2540_), .B(_2537_), .Y(_2541_) );
AOI21X1 AOI21X1_261 ( .A(_2622_), .B(_2623_), .C(_2621_), .Y(_2542_) );
OAI21X1 OAI21X1_423 ( .A(_2542_), .B(_2611_), .C(_2624_), .Y(_2543_) );
NOR3X1 NOR3X1_71 ( .A(_2601_), .B(_2610_), .C(_2542_), .Y(_2544_) );
NOR2X1 NOR2X1_269 ( .A(_2543_), .B(_2544_), .Y(_2545_) );
XNOR2X1 XNOR2X1_177 ( .A(_2545_), .B(_2541_), .Y(micro_ucr_hash1_c_24__4_) );
NAND3X1 NAND3X1_390 ( .A(_2627_), .B(_2631_), .C(_2626_), .Y(_2546_) );
OAI21X1 OAI21X1_424 ( .A(_2545_), .B(_2537_), .C(_2546_), .Y(_2547_) );
INVX1 INVX1_330 ( .A(micro_ucr_hash1_W_24__5_), .Y(_2548_) );
OAI21X1 OAI21X1_425 ( .A(micro_ucr_hash1_b_23__5_), .B(micro_ucr_hash1_a_23__5_), .C(_2548_), .Y(_2549_) );
NOR2X1 NOR2X1_270 ( .A(micro_ucr_hash1_b_23__5_), .B(micro_ucr_hash1_a_23__5_), .Y(_2550_) );
NAND2X1 NAND2X1_465 ( .A(micro_ucr_hash1_W_24__5_), .B(_2550_), .Y(_2551_) );
NAND3X1 NAND3X1_391 ( .A(_2627_), .B(_2549_), .C(_2551_), .Y(_2552_) );
INVX1 INVX1_331 ( .A(_2627_), .Y(_2553_) );
NAND2X1 NAND2X1_466 ( .A(_2548_), .B(_2550_), .Y(_2554_) );
OAI21X1 OAI21X1_426 ( .A(micro_ucr_hash1_b_23__5_), .B(micro_ucr_hash1_a_23__5_), .C(micro_ucr_hash1_W_24__5_), .Y(_2555_) );
NAND3X1 NAND3X1_392 ( .A(_2555_), .B(_2554_), .C(_2553_), .Y(_2556_) );
NAND2X1 NAND2X1_467 ( .A(_2552_), .B(_2556_), .Y(_2557_) );
XOR2X1 XOR2X1_233 ( .A(_2547_), .B(_2557_), .Y(micro_ucr_hash1_c_24__5_) );
OAI21X1 OAI21X1_427 ( .A(gnd), .B(micro_ucr_hash1_a_23__2_), .C(_2607_), .Y(_2558_) );
NAND2X1 NAND2X1_468 ( .A(micro_ucr_hash1_W_24__2_), .B(_2608_), .Y(_2559_) );
AOI21X1 AOI21X1_262 ( .A(_2558_), .B(_2559_), .C(_2597_), .Y(_2560_) );
INVX1 INVX1_332 ( .A(_2624_), .Y(_2561_) );
AOI21X1 AOI21X1_263 ( .A(_2620_), .B(_2560_), .C(_2561_), .Y(_2562_) );
NOR3X1 NOR3X1_72 ( .A(_2602_), .B(_2603_), .C(_2604_), .Y(_2563_) );
NAND3X1 NAND3X1_393 ( .A(_2613_), .B(_2620_), .C(_2563_), .Y(_2564_) );
NAND2X1 NAND2X1_469 ( .A(_2557_), .B(_2541_), .Y(_2565_) );
AOI21X1 AOI21X1_264 ( .A(_2562_), .B(_2564_), .C(_2565_), .Y(_2566_) );
AOI22X1 AOI22X1_15 ( .A(_2554_), .B(_2555_), .C(_2546_), .D(_2627_), .Y(_2567_) );
INVX1 INVX1_333 ( .A(_2554_), .Y(_2568_) );
OAI21X1 OAI21X1_428 ( .A(micro_ucr_hash1_b_23__6_), .B(micro_ucr_hash1_a_23__6_), .C(micro_ucr_hash1_W_24__6_), .Y(_2569_) );
INVX1 INVX1_334 ( .A(micro_ucr_hash1_W_24__6_), .Y(_2570_) );
NOR2X1 NOR2X1_271 ( .A(micro_ucr_hash1_b_23__6_), .B(micro_ucr_hash1_a_23__6_), .Y(_2571_) );
NAND2X1 NAND2X1_470 ( .A(_2570_), .B(_2571_), .Y(_2572_) );
NAND2X1 NAND2X1_471 ( .A(_2569_), .B(_2572_), .Y(_2573_) );
NOR2X1 NOR2X1_272 ( .A(_2568_), .B(_2573_), .Y(_2574_) );
INVX1 INVX1_335 ( .A(_2574_), .Y(_2575_) );
NAND2X1 NAND2X1_472 ( .A(_2568_), .B(_2573_), .Y(_2576_) );
NAND2X1 NAND2X1_473 ( .A(_2576_), .B(_2575_), .Y(_2577_) );
INVX1 INVX1_336 ( .A(_2577_), .Y(_2578_) );
OAI21X1 OAI21X1_429 ( .A(_2566_), .B(_2567_), .C(_2578_), .Y(_2579_) );
NAND3X1 NAND3X1_394 ( .A(_2622_), .B(_2538_), .C(_2539_), .Y(_2580_) );
NAND2X1 NAND2X1_474 ( .A(_2580_), .B(_2546_), .Y(_2581_) );
AOI21X1 AOI21X1_265 ( .A(_2552_), .B(_2556_), .C(_2581_), .Y(_2582_) );
OAI21X1 OAI21X1_430 ( .A(_2543_), .B(_2544_), .C(_2582_), .Y(_2583_) );
INVX1 INVX1_337 ( .A(_2567_), .Y(_2584_) );
NAND3X1 NAND3X1_395 ( .A(_2584_), .B(_2577_), .C(_2583_), .Y(_2585_) );
AND2X2 AND2X2_129 ( .A(_2579_), .B(_2585_), .Y(micro_ucr_hash1_c_24__6_) );
AOI21X1 AOI21X1_266 ( .A(_2584_), .B(_2583_), .C(_2577_), .Y(_2586_) );
NOR2X1 NOR2X1_273 ( .A(micro_ucr_hash1_b_23__7_), .B(micro_ucr_hash1_a_23__7_), .Y(_2587_) );
XNOR2X1 XNOR2X1_178 ( .A(_2587_), .B(micro_ucr_hash1_W_24__7_), .Y(_2588_) );
XNOR2X1 XNOR2X1_179 ( .A(_2588_), .B(_2569_), .Y(_2589_) );
OAI21X1 OAI21X1_431 ( .A(_2586_), .B(_2574_), .C(_2589_), .Y(_2590_) );
INVX1 INVX1_338 ( .A(_2589_), .Y(_2591_) );
NAND3X1 NAND3X1_396 ( .A(_2575_), .B(_2591_), .C(_2579_), .Y(_2592_) );
NAND2X1 NAND2X1_475 ( .A(_2590_), .B(_2592_), .Y(micro_ucr_hash1_c_24__7_) );
XOR2X1 XOR2X1_234 ( .A(micro_ucr_hash1_b_25__4_), .B(gnd), .Y(micro_ucr_hash1_a_25__0_) );
XOR2X1 XOR2X1_235 ( .A(micro_ucr_hash1_b_25__5_), .B(gnd), .Y(micro_ucr_hash1_a_25__1_) );
XOR2X1 XOR2X1_236 ( .A(micro_ucr_hash1_b_25__6_), .B(gnd), .Y(micro_ucr_hash1_a_25__2_) );
XOR2X1 XOR2X1_237 ( .A(micro_ucr_hash1_b_25__7_), .B(gnd), .Y(micro_ucr_hash1_a_25__3_) );
XOR2X1 XOR2X1_238 ( .A(micro_ucr_hash1_c_24__4_), .B(micro_ucr_hash1_b_24__4_), .Y(micro_ucr_hash1_a_25__4_) );
XOR2X1 XOR2X1_239 ( .A(micro_ucr_hash1_c_24__5_), .B(micro_ucr_hash1_b_24__5_), .Y(micro_ucr_hash1_a_25__5_) );
XOR2X1 XOR2X1_240 ( .A(micro_ucr_hash1_c_24__6_), .B(micro_ucr_hash1_b_24__6_), .Y(micro_ucr_hash1_a_25__6_) );
XOR2X1 XOR2X1_241 ( .A(micro_ucr_hash1_c_24__7_), .B(micro_ucr_hash1_b_24__7_), .Y(micro_ucr_hash1_a_25__7_) );
INVX1 INVX1_339 ( .A(micro_ucr_hash1_W_25__0_), .Y(_2688_) );
NOR2X1 NOR2X1_274 ( .A(gnd), .B(micro_ucr_hash1_a_24__0_), .Y(_2689_) );
NAND2X1 NAND2X1_476 ( .A(_2688_), .B(_2689_), .Y(_2690_) );
OAI21X1 OAI21X1_432 ( .A(gnd), .B(micro_ucr_hash1_a_24__0_), .C(micro_ucr_hash1_W_25__0_), .Y(_2691_) );
NAND2X1 NAND2X1_477 ( .A(_2691_), .B(_2690_), .Y(micro_ucr_hash1_b_26__4_) );
OAI21X1 OAI21X1_433 ( .A(gnd), .B(micro_ucr_hash1_a_24__1_), .C(micro_ucr_hash1_W_25__1_), .Y(_2692_) );
INVX1 INVX1_340 ( .A(micro_ucr_hash1_W_25__1_), .Y(_2693_) );
NOR2X1 NOR2X1_275 ( .A(gnd), .B(micro_ucr_hash1_a_24__1_), .Y(_2694_) );
NAND2X1 NAND2X1_478 ( .A(_2693_), .B(_2694_), .Y(_2695_) );
NAND3X1 NAND3X1_397 ( .A(_2692_), .B(_2690_), .C(_2695_), .Y(_2696_) );
AND2X2 AND2X2_130 ( .A(_2689_), .B(_2688_), .Y(_2697_) );
INVX2 INVX2_67 ( .A(_2692_), .Y(_2698_) );
AND2X2 AND2X2_131 ( .A(_2694_), .B(_2693_), .Y(_2699_) );
OAI21X1 OAI21X1_434 ( .A(_2699_), .B(_2698_), .C(_2697_), .Y(_2700_) );
AND2X2 AND2X2_132 ( .A(_2700_), .B(_2696_), .Y(micro_ucr_hash1_b_26__5_) );
OAI21X1 OAI21X1_435 ( .A(gnd), .B(micro_ucr_hash1_a_24__2_), .C(micro_ucr_hash1_W_25__2_), .Y(_2701_) );
INVX1 INVX1_341 ( .A(micro_ucr_hash1_W_25__2_), .Y(_2702_) );
NOR2X1 NOR2X1_276 ( .A(gnd), .B(micro_ucr_hash1_a_24__2_), .Y(_2703_) );
NAND2X1 NAND2X1_479 ( .A(_2702_), .B(_2703_), .Y(_2704_) );
NAND2X1 NAND2X1_480 ( .A(_2701_), .B(_2704_), .Y(_2705_) );
NAND3X1 NAND3X1_398 ( .A(_2701_), .B(_2704_), .C(_2698_), .Y(_2706_) );
OAI21X1 OAI21X1_436 ( .A(_2696_), .B(_2705_), .C(_2706_), .Y(_2707_) );
INVX1 INVX1_342 ( .A(_2705_), .Y(_2708_) );
OAI21X1 OAI21X1_437 ( .A(_2697_), .B(_2699_), .C(_2692_), .Y(_2709_) );
NOR2X1 NOR2X1_277 ( .A(_2709_), .B(_2708_), .Y(_2710_) );
NOR2X1 NOR2X1_278 ( .A(_2707_), .B(_2710_), .Y(micro_ucr_hash1_b_26__6_) );
INVX1 INVX1_343 ( .A(micro_ucr_hash1_W_25__3_), .Y(_2711_) );
OAI21X1 OAI21X1_438 ( .A(gnd), .B(micro_ucr_hash1_a_24__3_), .C(_2711_), .Y(_2712_) );
NOR2X1 NOR2X1_279 ( .A(gnd), .B(micro_ucr_hash1_a_24__3_), .Y(_2713_) );
NAND2X1 NAND2X1_481 ( .A(micro_ucr_hash1_W_25__3_), .B(_2713_), .Y(_2714_) );
NAND3X1 NAND3X1_399 ( .A(_2701_), .B(_2712_), .C(_2714_), .Y(_2715_) );
INVX1 INVX1_344 ( .A(_2701_), .Y(_2716_) );
OAI21X1 OAI21X1_439 ( .A(gnd), .B(micro_ucr_hash1_a_24__3_), .C(micro_ucr_hash1_W_25__3_), .Y(_2717_) );
NAND2X1 NAND2X1_482 ( .A(_2711_), .B(_2713_), .Y(_2718_) );
NAND3X1 NAND3X1_400 ( .A(_2717_), .B(_2718_), .C(_2716_), .Y(_2719_) );
NAND2X1 NAND2X1_483 ( .A(_2715_), .B(_2719_), .Y(_2720_) );
XNOR2X1 XNOR2X1_180 ( .A(_2707_), .B(_2720_), .Y(micro_ucr_hash1_b_26__7_) );
INVX1 INVX1_345 ( .A(_2717_), .Y(_2721_) );
OAI21X1 OAI21X1_440 ( .A(micro_ucr_hash1_b_24__4_), .B(micro_ucr_hash1_a_24__4_), .C(micro_ucr_hash1_W_25__4_), .Y(_2722_) );
INVX1 INVX1_346 ( .A(micro_ucr_hash1_b_24__4_), .Y(_2723_) );
INVX1 INVX1_347 ( .A(micro_ucr_hash1_a_24__4_), .Y(_2724_) );
INVX1 INVX1_348 ( .A(micro_ucr_hash1_W_25__4_), .Y(_2725_) );
NAND3X1 NAND3X1_401 ( .A(_2723_), .B(_2724_), .C(_2725_), .Y(_2726_) );
AOI21X1 AOI21X1_267 ( .A(_2722_), .B(_2726_), .C(_2721_), .Y(_2632_) );
OAI21X1 OAI21X1_441 ( .A(micro_ucr_hash1_b_24__4_), .B(micro_ucr_hash1_a_24__4_), .C(_2725_), .Y(_2633_) );
NAND3X1 NAND3X1_402 ( .A(micro_ucr_hash1_W_25__4_), .B(_2723_), .C(_2724_), .Y(_2634_) );
AOI21X1 AOI21X1_268 ( .A(_2633_), .B(_2634_), .C(_2717_), .Y(_2635_) );
NOR2X1 NOR2X1_280 ( .A(_2635_), .B(_2632_), .Y(_2636_) );
AOI21X1 AOI21X1_269 ( .A(_2717_), .B(_2718_), .C(_2716_), .Y(_2637_) );
OAI21X1 OAI21X1_442 ( .A(_2637_), .B(_2706_), .C(_2719_), .Y(_2638_) );
NOR3X1 NOR3X1_73 ( .A(_2696_), .B(_2705_), .C(_2637_), .Y(_2639_) );
NOR2X1 NOR2X1_281 ( .A(_2638_), .B(_2639_), .Y(_2640_) );
XNOR2X1 XNOR2X1_181 ( .A(_2640_), .B(_2636_), .Y(micro_ucr_hash1_c_25__4_) );
NAND3X1 NAND3X1_403 ( .A(_2722_), .B(_2726_), .C(_2721_), .Y(_2641_) );
OAI21X1 OAI21X1_443 ( .A(_2640_), .B(_2632_), .C(_2641_), .Y(_2642_) );
INVX1 INVX1_349 ( .A(micro_ucr_hash1_W_25__5_), .Y(_2643_) );
OAI21X1 OAI21X1_444 ( .A(micro_ucr_hash1_b_24__5_), .B(micro_ucr_hash1_a_24__5_), .C(_2643_), .Y(_2644_) );
NOR2X1 NOR2X1_282 ( .A(micro_ucr_hash1_b_24__5_), .B(micro_ucr_hash1_a_24__5_), .Y(_2645_) );
NAND2X1 NAND2X1_484 ( .A(micro_ucr_hash1_W_25__5_), .B(_2645_), .Y(_2646_) );
NAND3X1 NAND3X1_404 ( .A(_2722_), .B(_2644_), .C(_2646_), .Y(_2647_) );
INVX1 INVX1_350 ( .A(_2722_), .Y(_2648_) );
NAND2X1 NAND2X1_485 ( .A(_2643_), .B(_2645_), .Y(_2649_) );
OAI21X1 OAI21X1_445 ( .A(micro_ucr_hash1_b_24__5_), .B(micro_ucr_hash1_a_24__5_), .C(micro_ucr_hash1_W_25__5_), .Y(_2650_) );
NAND3X1 NAND3X1_405 ( .A(_2650_), .B(_2649_), .C(_2648_), .Y(_2651_) );
NAND2X1 NAND2X1_486 ( .A(_2647_), .B(_2651_), .Y(_2652_) );
XOR2X1 XOR2X1_242 ( .A(_2642_), .B(_2652_), .Y(micro_ucr_hash1_c_25__5_) );
OAI21X1 OAI21X1_446 ( .A(gnd), .B(micro_ucr_hash1_a_24__2_), .C(_2702_), .Y(_2653_) );
NAND2X1 NAND2X1_487 ( .A(micro_ucr_hash1_W_25__2_), .B(_2703_), .Y(_2654_) );
AOI21X1 AOI21X1_270 ( .A(_2653_), .B(_2654_), .C(_2692_), .Y(_2655_) );
INVX1 INVX1_351 ( .A(_2719_), .Y(_2656_) );
AOI21X1 AOI21X1_271 ( .A(_2715_), .B(_2655_), .C(_2656_), .Y(_2657_) );
NOR3X1 NOR3X1_74 ( .A(_2697_), .B(_2698_), .C(_2699_), .Y(_2658_) );
NAND3X1 NAND3X1_406 ( .A(_2708_), .B(_2715_), .C(_2658_), .Y(_2659_) );
NAND2X1 NAND2X1_488 ( .A(_2652_), .B(_2636_), .Y(_2660_) );
AOI21X1 AOI21X1_272 ( .A(_2657_), .B(_2659_), .C(_2660_), .Y(_2661_) );
AOI22X1 AOI22X1_16 ( .A(_2649_), .B(_2650_), .C(_2641_), .D(_2722_), .Y(_2662_) );
INVX1 INVX1_352 ( .A(_2649_), .Y(_2663_) );
OAI21X1 OAI21X1_447 ( .A(micro_ucr_hash1_b_24__6_), .B(micro_ucr_hash1_a_24__6_), .C(micro_ucr_hash1_W_25__6_), .Y(_2664_) );
INVX1 INVX1_353 ( .A(micro_ucr_hash1_W_25__6_), .Y(_2665_) );
NOR2X1 NOR2X1_283 ( .A(micro_ucr_hash1_b_24__6_), .B(micro_ucr_hash1_a_24__6_), .Y(_2666_) );
NAND2X1 NAND2X1_489 ( .A(_2665_), .B(_2666_), .Y(_2667_) );
NAND2X1 NAND2X1_490 ( .A(_2664_), .B(_2667_), .Y(_2668_) );
NOR2X1 NOR2X1_284 ( .A(_2663_), .B(_2668_), .Y(_2669_) );
INVX1 INVX1_354 ( .A(_2669_), .Y(_2670_) );
NAND2X1 NAND2X1_491 ( .A(_2663_), .B(_2668_), .Y(_2671_) );
NAND2X1 NAND2X1_492 ( .A(_2671_), .B(_2670_), .Y(_2672_) );
INVX1 INVX1_355 ( .A(_2672_), .Y(_2673_) );
OAI21X1 OAI21X1_448 ( .A(_2661_), .B(_2662_), .C(_2673_), .Y(_2674_) );
NAND3X1 NAND3X1_407 ( .A(_2717_), .B(_2633_), .C(_2634_), .Y(_2675_) );
NAND2X1 NAND2X1_493 ( .A(_2675_), .B(_2641_), .Y(_2676_) );
AOI21X1 AOI21X1_273 ( .A(_2647_), .B(_2651_), .C(_2676_), .Y(_2677_) );
OAI21X1 OAI21X1_449 ( .A(_2638_), .B(_2639_), .C(_2677_), .Y(_2678_) );
INVX1 INVX1_356 ( .A(_2662_), .Y(_2679_) );
NAND3X1 NAND3X1_408 ( .A(_2679_), .B(_2672_), .C(_2678_), .Y(_2680_) );
AND2X2 AND2X2_133 ( .A(_2674_), .B(_2680_), .Y(micro_ucr_hash1_c_25__6_) );
AOI21X1 AOI21X1_274 ( .A(_2679_), .B(_2678_), .C(_2672_), .Y(_2681_) );
NOR2X1 NOR2X1_285 ( .A(micro_ucr_hash1_b_24__7_), .B(micro_ucr_hash1_a_24__7_), .Y(_2682_) );
XNOR2X1 XNOR2X1_182 ( .A(_2682_), .B(micro_ucr_hash1_W_25__7_), .Y(_2683_) );
XNOR2X1 XNOR2X1_183 ( .A(_2683_), .B(_2664_), .Y(_2684_) );
OAI21X1 OAI21X1_450 ( .A(_2681_), .B(_2669_), .C(_2684_), .Y(_2685_) );
INVX1 INVX1_357 ( .A(_2684_), .Y(_2686_) );
NAND3X1 NAND3X1_409 ( .A(_2670_), .B(_2686_), .C(_2674_), .Y(_2687_) );
NAND2X1 NAND2X1_494 ( .A(_2685_), .B(_2687_), .Y(micro_ucr_hash1_c_25__7_) );
XOR2X1 XOR2X1_243 ( .A(micro_ucr_hash1_b_26__4_), .B(gnd), .Y(micro_ucr_hash1_a_26__0_) );
XOR2X1 XOR2X1_244 ( .A(micro_ucr_hash1_b_26__5_), .B(gnd), .Y(micro_ucr_hash1_a_26__1_) );
XOR2X1 XOR2X1_245 ( .A(micro_ucr_hash1_b_26__6_), .B(gnd), .Y(micro_ucr_hash1_a_26__2_) );
XOR2X1 XOR2X1_246 ( .A(micro_ucr_hash1_b_26__7_), .B(gnd), .Y(micro_ucr_hash1_a_26__3_) );
XOR2X1 XOR2X1_247 ( .A(micro_ucr_hash1_c_25__4_), .B(micro_ucr_hash1_b_25__4_), .Y(micro_ucr_hash1_a_26__4_) );
XOR2X1 XOR2X1_248 ( .A(micro_ucr_hash1_c_25__5_), .B(micro_ucr_hash1_b_25__5_), .Y(micro_ucr_hash1_a_26__5_) );
XOR2X1 XOR2X1_249 ( .A(micro_ucr_hash1_c_25__6_), .B(micro_ucr_hash1_b_25__6_), .Y(micro_ucr_hash1_a_26__6_) );
XOR2X1 XOR2X1_250 ( .A(micro_ucr_hash1_c_25__7_), .B(micro_ucr_hash1_b_25__7_), .Y(micro_ucr_hash1_a_26__7_) );
INVX1 INVX1_358 ( .A(micro_ucr_hash1_W_26__0_), .Y(_2783_) );
NOR2X1 NOR2X1_286 ( .A(gnd), .B(micro_ucr_hash1_a_25__0_), .Y(_2784_) );
NAND2X1 NAND2X1_495 ( .A(_2783_), .B(_2784_), .Y(_2785_) );
OAI21X1 OAI21X1_451 ( .A(gnd), .B(micro_ucr_hash1_a_25__0_), .C(micro_ucr_hash1_W_26__0_), .Y(_2786_) );
NAND2X1 NAND2X1_496 ( .A(_2786_), .B(_2785_), .Y(micro_ucr_hash1_b_27__4_) );
OAI21X1 OAI21X1_452 ( .A(gnd), .B(micro_ucr_hash1_a_25__1_), .C(micro_ucr_hash1_W_26__1_), .Y(_2787_) );
INVX1 INVX1_359 ( .A(micro_ucr_hash1_W_26__1_), .Y(_2788_) );
NOR2X1 NOR2X1_287 ( .A(gnd), .B(micro_ucr_hash1_a_25__1_), .Y(_2789_) );
NAND2X1 NAND2X1_497 ( .A(_2788_), .B(_2789_), .Y(_2790_) );
NAND3X1 NAND3X1_410 ( .A(_2787_), .B(_2785_), .C(_2790_), .Y(_2791_) );
AND2X2 AND2X2_134 ( .A(_2784_), .B(_2783_), .Y(_2792_) );
INVX2 INVX2_68 ( .A(_2787_), .Y(_2793_) );
AND2X2 AND2X2_135 ( .A(_2789_), .B(_2788_), .Y(_2794_) );
OAI21X1 OAI21X1_453 ( .A(_2794_), .B(_2793_), .C(_2792_), .Y(_2795_) );
AND2X2 AND2X2_136 ( .A(_2795_), .B(_2791_), .Y(micro_ucr_hash1_b_27__5_) );
OAI21X1 OAI21X1_454 ( .A(gnd), .B(micro_ucr_hash1_a_25__2_), .C(micro_ucr_hash1_W_26__2_), .Y(_2796_) );
INVX1 INVX1_360 ( .A(micro_ucr_hash1_W_26__2_), .Y(_2797_) );
NOR2X1 NOR2X1_288 ( .A(gnd), .B(micro_ucr_hash1_a_25__2_), .Y(_2798_) );
NAND2X1 NAND2X1_498 ( .A(_2797_), .B(_2798_), .Y(_2799_) );
NAND2X1 NAND2X1_499 ( .A(_2796_), .B(_2799_), .Y(_2800_) );
NAND3X1 NAND3X1_411 ( .A(_2796_), .B(_2799_), .C(_2793_), .Y(_2801_) );
OAI21X1 OAI21X1_455 ( .A(_2791_), .B(_2800_), .C(_2801_), .Y(_2802_) );
INVX1 INVX1_361 ( .A(_2800_), .Y(_2803_) );
OAI21X1 OAI21X1_456 ( .A(_2792_), .B(_2794_), .C(_2787_), .Y(_2804_) );
NOR2X1 NOR2X1_289 ( .A(_2804_), .B(_2803_), .Y(_2805_) );
NOR2X1 NOR2X1_290 ( .A(_2802_), .B(_2805_), .Y(micro_ucr_hash1_b_27__6_) );
INVX1 INVX1_362 ( .A(micro_ucr_hash1_W_26__3_), .Y(_2806_) );
OAI21X1 OAI21X1_457 ( .A(gnd), .B(micro_ucr_hash1_a_25__3_), .C(_2806_), .Y(_2807_) );
NOR2X1 NOR2X1_291 ( .A(gnd), .B(micro_ucr_hash1_a_25__3_), .Y(_2808_) );
NAND2X1 NAND2X1_500 ( .A(micro_ucr_hash1_W_26__3_), .B(_2808_), .Y(_2809_) );
NAND3X1 NAND3X1_412 ( .A(_2796_), .B(_2807_), .C(_2809_), .Y(_2810_) );
INVX1 INVX1_363 ( .A(_2796_), .Y(_2811_) );
OAI21X1 OAI21X1_458 ( .A(gnd), .B(micro_ucr_hash1_a_25__3_), .C(micro_ucr_hash1_W_26__3_), .Y(_2812_) );
NAND2X1 NAND2X1_501 ( .A(_2806_), .B(_2808_), .Y(_2813_) );
NAND3X1 NAND3X1_413 ( .A(_2812_), .B(_2813_), .C(_2811_), .Y(_2814_) );
NAND2X1 NAND2X1_502 ( .A(_2810_), .B(_2814_), .Y(_2815_) );
XNOR2X1 XNOR2X1_184 ( .A(_2802_), .B(_2815_), .Y(micro_ucr_hash1_b_27__7_) );
INVX1 INVX1_364 ( .A(_2812_), .Y(_2816_) );
OAI21X1 OAI21X1_459 ( .A(micro_ucr_hash1_b_25__4_), .B(micro_ucr_hash1_a_25__4_), .C(micro_ucr_hash1_W_26__4_), .Y(_2817_) );
INVX1 INVX1_365 ( .A(micro_ucr_hash1_b_25__4_), .Y(_2818_) );
INVX1 INVX1_366 ( .A(micro_ucr_hash1_a_25__4_), .Y(_2819_) );
INVX1 INVX1_367 ( .A(micro_ucr_hash1_W_26__4_), .Y(_2820_) );
NAND3X1 NAND3X1_414 ( .A(_2818_), .B(_2819_), .C(_2820_), .Y(_2821_) );
AOI21X1 AOI21X1_275 ( .A(_2817_), .B(_2821_), .C(_2816_), .Y(_2727_) );
OAI21X1 OAI21X1_460 ( .A(micro_ucr_hash1_b_25__4_), .B(micro_ucr_hash1_a_25__4_), .C(_2820_), .Y(_2728_) );
NAND3X1 NAND3X1_415 ( .A(micro_ucr_hash1_W_26__4_), .B(_2818_), .C(_2819_), .Y(_2729_) );
AOI21X1 AOI21X1_276 ( .A(_2728_), .B(_2729_), .C(_2812_), .Y(_2730_) );
NOR2X1 NOR2X1_292 ( .A(_2730_), .B(_2727_), .Y(_2731_) );
AOI21X1 AOI21X1_277 ( .A(_2812_), .B(_2813_), .C(_2811_), .Y(_2732_) );
OAI21X1 OAI21X1_461 ( .A(_2732_), .B(_2801_), .C(_2814_), .Y(_2733_) );
NOR3X1 NOR3X1_75 ( .A(_2791_), .B(_2800_), .C(_2732_), .Y(_2734_) );
NOR2X1 NOR2X1_293 ( .A(_2733_), .B(_2734_), .Y(_2735_) );
XNOR2X1 XNOR2X1_185 ( .A(_2735_), .B(_2731_), .Y(micro_ucr_hash1_c_26__4_) );
NAND3X1 NAND3X1_416 ( .A(_2817_), .B(_2821_), .C(_2816_), .Y(_2736_) );
OAI21X1 OAI21X1_462 ( .A(_2735_), .B(_2727_), .C(_2736_), .Y(_2737_) );
INVX1 INVX1_368 ( .A(micro_ucr_hash1_W_26__5_), .Y(_2738_) );
OAI21X1 OAI21X1_463 ( .A(micro_ucr_hash1_b_25__5_), .B(micro_ucr_hash1_a_25__5_), .C(_2738_), .Y(_2739_) );
NOR2X1 NOR2X1_294 ( .A(micro_ucr_hash1_b_25__5_), .B(micro_ucr_hash1_a_25__5_), .Y(_2740_) );
NAND2X1 NAND2X1_503 ( .A(micro_ucr_hash1_W_26__5_), .B(_2740_), .Y(_2741_) );
NAND3X1 NAND3X1_417 ( .A(_2817_), .B(_2739_), .C(_2741_), .Y(_2742_) );
INVX1 INVX1_369 ( .A(_2817_), .Y(_2743_) );
NAND2X1 NAND2X1_504 ( .A(_2738_), .B(_2740_), .Y(_2744_) );
OAI21X1 OAI21X1_464 ( .A(micro_ucr_hash1_b_25__5_), .B(micro_ucr_hash1_a_25__5_), .C(micro_ucr_hash1_W_26__5_), .Y(_2745_) );
NAND3X1 NAND3X1_418 ( .A(_2745_), .B(_2744_), .C(_2743_), .Y(_2746_) );
NAND2X1 NAND2X1_505 ( .A(_2742_), .B(_2746_), .Y(_2747_) );
XOR2X1 XOR2X1_251 ( .A(_2737_), .B(_2747_), .Y(micro_ucr_hash1_c_26__5_) );
OAI21X1 OAI21X1_465 ( .A(gnd), .B(micro_ucr_hash1_a_25__2_), .C(_2797_), .Y(_2748_) );
NAND2X1 NAND2X1_506 ( .A(micro_ucr_hash1_W_26__2_), .B(_2798_), .Y(_2749_) );
AOI21X1 AOI21X1_278 ( .A(_2748_), .B(_2749_), .C(_2787_), .Y(_2750_) );
INVX1 INVX1_370 ( .A(_2814_), .Y(_2751_) );
AOI21X1 AOI21X1_279 ( .A(_2810_), .B(_2750_), .C(_2751_), .Y(_2752_) );
NOR3X1 NOR3X1_76 ( .A(_2792_), .B(_2793_), .C(_2794_), .Y(_2753_) );
NAND3X1 NAND3X1_419 ( .A(_2803_), .B(_2810_), .C(_2753_), .Y(_2754_) );
NAND2X1 NAND2X1_507 ( .A(_2747_), .B(_2731_), .Y(_2755_) );
AOI21X1 AOI21X1_280 ( .A(_2752_), .B(_2754_), .C(_2755_), .Y(_2756_) );
AOI22X1 AOI22X1_17 ( .A(_2744_), .B(_2745_), .C(_2736_), .D(_2817_), .Y(_2757_) );
INVX1 INVX1_371 ( .A(_2744_), .Y(_2758_) );
OAI21X1 OAI21X1_466 ( .A(micro_ucr_hash1_b_25__6_), .B(micro_ucr_hash1_a_25__6_), .C(micro_ucr_hash1_W_26__6_), .Y(_2759_) );
INVX1 INVX1_372 ( .A(micro_ucr_hash1_W_26__6_), .Y(_2760_) );
NOR2X1 NOR2X1_295 ( .A(micro_ucr_hash1_b_25__6_), .B(micro_ucr_hash1_a_25__6_), .Y(_2761_) );
NAND2X1 NAND2X1_508 ( .A(_2760_), .B(_2761_), .Y(_2762_) );
NAND2X1 NAND2X1_509 ( .A(_2759_), .B(_2762_), .Y(_2763_) );
NOR2X1 NOR2X1_296 ( .A(_2758_), .B(_2763_), .Y(_2764_) );
INVX1 INVX1_373 ( .A(_2764_), .Y(_2765_) );
NAND2X1 NAND2X1_510 ( .A(_2758_), .B(_2763_), .Y(_2766_) );
NAND2X1 NAND2X1_511 ( .A(_2766_), .B(_2765_), .Y(_2767_) );
INVX1 INVX1_374 ( .A(_2767_), .Y(_2768_) );
OAI21X1 OAI21X1_467 ( .A(_2756_), .B(_2757_), .C(_2768_), .Y(_2769_) );
NAND3X1 NAND3X1_420 ( .A(_2812_), .B(_2728_), .C(_2729_), .Y(_2770_) );
NAND2X1 NAND2X1_512 ( .A(_2770_), .B(_2736_), .Y(_2771_) );
AOI21X1 AOI21X1_281 ( .A(_2742_), .B(_2746_), .C(_2771_), .Y(_2772_) );
OAI21X1 OAI21X1_468 ( .A(_2733_), .B(_2734_), .C(_2772_), .Y(_2773_) );
INVX1 INVX1_375 ( .A(_2757_), .Y(_2774_) );
NAND3X1 NAND3X1_421 ( .A(_2774_), .B(_2767_), .C(_2773_), .Y(_2775_) );
AND2X2 AND2X2_137 ( .A(_2769_), .B(_2775_), .Y(micro_ucr_hash1_c_26__6_) );
AOI21X1 AOI21X1_282 ( .A(_2774_), .B(_2773_), .C(_2767_), .Y(_2776_) );
NOR2X1 NOR2X1_297 ( .A(micro_ucr_hash1_b_25__7_), .B(micro_ucr_hash1_a_25__7_), .Y(_2777_) );
XNOR2X1 XNOR2X1_186 ( .A(_2777_), .B(micro_ucr_hash1_W_26__7_), .Y(_2778_) );
XNOR2X1 XNOR2X1_187 ( .A(_2778_), .B(_2759_), .Y(_2779_) );
OAI21X1 OAI21X1_469 ( .A(_2776_), .B(_2764_), .C(_2779_), .Y(_2780_) );
INVX1 INVX1_376 ( .A(_2779_), .Y(_2781_) );
NAND3X1 NAND3X1_422 ( .A(_2765_), .B(_2781_), .C(_2769_), .Y(_2782_) );
NAND2X1 NAND2X1_513 ( .A(_2780_), .B(_2782_), .Y(micro_ucr_hash1_c_26__7_) );
XOR2X1 XOR2X1_252 ( .A(micro_ucr_hash1_b_27__4_), .B(gnd), .Y(micro_ucr_hash1_a_27__0_) );
XOR2X1 XOR2X1_253 ( .A(micro_ucr_hash1_b_27__5_), .B(gnd), .Y(micro_ucr_hash1_a_27__1_) );
XOR2X1 XOR2X1_254 ( .A(micro_ucr_hash1_b_27__6_), .B(gnd), .Y(micro_ucr_hash1_a_27__2_) );
XOR2X1 XOR2X1_255 ( .A(micro_ucr_hash1_b_27__7_), .B(gnd), .Y(micro_ucr_hash1_a_27__3_) );
XOR2X1 XOR2X1_256 ( .A(micro_ucr_hash1_c_26__4_), .B(micro_ucr_hash1_b_26__4_), .Y(micro_ucr_hash1_a_27__4_) );
XOR2X1 XOR2X1_257 ( .A(micro_ucr_hash1_c_26__5_), .B(micro_ucr_hash1_b_26__5_), .Y(micro_ucr_hash1_a_27__5_) );
XOR2X1 XOR2X1_258 ( .A(micro_ucr_hash1_c_26__6_), .B(micro_ucr_hash1_b_26__6_), .Y(micro_ucr_hash1_a_27__6_) );
XOR2X1 XOR2X1_259 ( .A(micro_ucr_hash1_c_26__7_), .B(micro_ucr_hash1_b_26__7_), .Y(micro_ucr_hash1_a_27__7_) );
INVX1 INVX1_377 ( .A(micro_ucr_hash1_W_27__0_), .Y(_2878_) );
NOR2X1 NOR2X1_298 ( .A(gnd), .B(micro_ucr_hash1_a_26__0_), .Y(_2879_) );
NAND2X1 NAND2X1_514 ( .A(_2878_), .B(_2879_), .Y(_2880_) );
OAI21X1 OAI21X1_470 ( .A(gnd), .B(micro_ucr_hash1_a_26__0_), .C(micro_ucr_hash1_W_27__0_), .Y(_2881_) );
NAND2X1 NAND2X1_515 ( .A(_2881_), .B(_2880_), .Y(micro_ucr_hash1_b_28__4_) );
OAI21X1 OAI21X1_471 ( .A(gnd), .B(micro_ucr_hash1_a_26__1_), .C(micro_ucr_hash1_W_27__1_), .Y(_2882_) );
INVX1 INVX1_378 ( .A(micro_ucr_hash1_W_27__1_), .Y(_2883_) );
NOR2X1 NOR2X1_299 ( .A(gnd), .B(micro_ucr_hash1_a_26__1_), .Y(_2884_) );
NAND2X1 NAND2X1_516 ( .A(_2883_), .B(_2884_), .Y(_2885_) );
NAND3X1 NAND3X1_423 ( .A(_2882_), .B(_2880_), .C(_2885_), .Y(_2886_) );
AND2X2 AND2X2_138 ( .A(_2879_), .B(_2878_), .Y(_2887_) );
INVX2 INVX2_69 ( .A(_2882_), .Y(_2888_) );
AND2X2 AND2X2_139 ( .A(_2884_), .B(_2883_), .Y(_2889_) );
OAI21X1 OAI21X1_472 ( .A(_2889_), .B(_2888_), .C(_2887_), .Y(_2890_) );
AND2X2 AND2X2_140 ( .A(_2890_), .B(_2886_), .Y(micro_ucr_hash1_b_28__5_) );
OAI21X1 OAI21X1_473 ( .A(gnd), .B(micro_ucr_hash1_a_26__2_), .C(micro_ucr_hash1_W_27__2_), .Y(_2891_) );
INVX1 INVX1_379 ( .A(micro_ucr_hash1_W_27__2_), .Y(_2892_) );
NOR2X1 NOR2X1_300 ( .A(gnd), .B(micro_ucr_hash1_a_26__2_), .Y(_2893_) );
NAND2X1 NAND2X1_517 ( .A(_2892_), .B(_2893_), .Y(_2894_) );
NAND2X1 NAND2X1_518 ( .A(_2891_), .B(_2894_), .Y(_2895_) );
NAND3X1 NAND3X1_424 ( .A(_2891_), .B(_2894_), .C(_2888_), .Y(_2896_) );
OAI21X1 OAI21X1_474 ( .A(_2886_), .B(_2895_), .C(_2896_), .Y(_2897_) );
INVX1 INVX1_380 ( .A(_2895_), .Y(_2898_) );
OAI21X1 OAI21X1_475 ( .A(_2887_), .B(_2889_), .C(_2882_), .Y(_2899_) );
NOR2X1 NOR2X1_301 ( .A(_2899_), .B(_2898_), .Y(_2900_) );
NOR2X1 NOR2X1_302 ( .A(_2897_), .B(_2900_), .Y(micro_ucr_hash1_b_28__6_) );
INVX1 INVX1_381 ( .A(micro_ucr_hash1_W_27__3_), .Y(_2901_) );
OAI21X1 OAI21X1_476 ( .A(gnd), .B(micro_ucr_hash1_a_26__3_), .C(_2901_), .Y(_2902_) );
NOR2X1 NOR2X1_303 ( .A(gnd), .B(micro_ucr_hash1_a_26__3_), .Y(_2903_) );
NAND2X1 NAND2X1_519 ( .A(micro_ucr_hash1_W_27__3_), .B(_2903_), .Y(_2904_) );
NAND3X1 NAND3X1_425 ( .A(_2891_), .B(_2902_), .C(_2904_), .Y(_2905_) );
INVX1 INVX1_382 ( .A(_2891_), .Y(_2906_) );
OAI21X1 OAI21X1_477 ( .A(gnd), .B(micro_ucr_hash1_a_26__3_), .C(micro_ucr_hash1_W_27__3_), .Y(_2907_) );
NAND2X1 NAND2X1_520 ( .A(_2901_), .B(_2903_), .Y(_2908_) );
NAND3X1 NAND3X1_426 ( .A(_2907_), .B(_2908_), .C(_2906_), .Y(_2909_) );
NAND2X1 NAND2X1_521 ( .A(_2905_), .B(_2909_), .Y(_2910_) );
XNOR2X1 XNOR2X1_188 ( .A(_2897_), .B(_2910_), .Y(micro_ucr_hash1_b_28__7_) );
INVX1 INVX1_383 ( .A(_2907_), .Y(_2911_) );
OAI21X1 OAI21X1_478 ( .A(micro_ucr_hash1_b_26__4_), .B(micro_ucr_hash1_a_26__4_), .C(micro_ucr_hash1_W_27__4_), .Y(_2912_) );
INVX1 INVX1_384 ( .A(micro_ucr_hash1_b_26__4_), .Y(_2913_) );
INVX1 INVX1_385 ( .A(micro_ucr_hash1_a_26__4_), .Y(_2914_) );
INVX1 INVX1_386 ( .A(micro_ucr_hash1_W_27__4_), .Y(_2915_) );
NAND3X1 NAND3X1_427 ( .A(_2913_), .B(_2914_), .C(_2915_), .Y(_2916_) );
AOI21X1 AOI21X1_283 ( .A(_2912_), .B(_2916_), .C(_2911_), .Y(_2822_) );
OAI21X1 OAI21X1_479 ( .A(micro_ucr_hash1_b_26__4_), .B(micro_ucr_hash1_a_26__4_), .C(_2915_), .Y(_2823_) );
NAND3X1 NAND3X1_428 ( .A(micro_ucr_hash1_W_27__4_), .B(_2913_), .C(_2914_), .Y(_2824_) );
AOI21X1 AOI21X1_284 ( .A(_2823_), .B(_2824_), .C(_2907_), .Y(_2825_) );
NOR2X1 NOR2X1_304 ( .A(_2825_), .B(_2822_), .Y(_2826_) );
AOI21X1 AOI21X1_285 ( .A(_2907_), .B(_2908_), .C(_2906_), .Y(_2827_) );
OAI21X1 OAI21X1_480 ( .A(_2827_), .B(_2896_), .C(_2909_), .Y(_2828_) );
NOR3X1 NOR3X1_77 ( .A(_2886_), .B(_2895_), .C(_2827_), .Y(_2829_) );
NOR2X1 NOR2X1_305 ( .A(_2828_), .B(_2829_), .Y(_2830_) );
XNOR2X1 XNOR2X1_189 ( .A(_2830_), .B(_2826_), .Y(micro_ucr_hash1_c_27__4_) );
NAND3X1 NAND3X1_429 ( .A(_2912_), .B(_2916_), .C(_2911_), .Y(_2831_) );
OAI21X1 OAI21X1_481 ( .A(_2830_), .B(_2822_), .C(_2831_), .Y(_2832_) );
INVX1 INVX1_387 ( .A(micro_ucr_hash1_W_27__5_), .Y(_2833_) );
OAI21X1 OAI21X1_482 ( .A(micro_ucr_hash1_b_26__5_), .B(micro_ucr_hash1_a_26__5_), .C(_2833_), .Y(_2834_) );
NOR2X1 NOR2X1_306 ( .A(micro_ucr_hash1_b_26__5_), .B(micro_ucr_hash1_a_26__5_), .Y(_2835_) );
NAND2X1 NAND2X1_522 ( .A(micro_ucr_hash1_W_27__5_), .B(_2835_), .Y(_2836_) );
NAND3X1 NAND3X1_430 ( .A(_2912_), .B(_2834_), .C(_2836_), .Y(_2837_) );
INVX1 INVX1_388 ( .A(_2912_), .Y(_2838_) );
NAND2X1 NAND2X1_523 ( .A(_2833_), .B(_2835_), .Y(_2839_) );
OAI21X1 OAI21X1_483 ( .A(micro_ucr_hash1_b_26__5_), .B(micro_ucr_hash1_a_26__5_), .C(micro_ucr_hash1_W_27__5_), .Y(_2840_) );
NAND3X1 NAND3X1_431 ( .A(_2840_), .B(_2839_), .C(_2838_), .Y(_2841_) );
NAND2X1 NAND2X1_524 ( .A(_2837_), .B(_2841_), .Y(_2842_) );
XOR2X1 XOR2X1_260 ( .A(_2832_), .B(_2842_), .Y(micro_ucr_hash1_c_27__5_) );
OAI21X1 OAI21X1_484 ( .A(gnd), .B(micro_ucr_hash1_a_26__2_), .C(_2892_), .Y(_2843_) );
NAND2X1 NAND2X1_525 ( .A(micro_ucr_hash1_W_27__2_), .B(_2893_), .Y(_2844_) );
AOI21X1 AOI21X1_286 ( .A(_2843_), .B(_2844_), .C(_2882_), .Y(_2845_) );
INVX1 INVX1_389 ( .A(_2909_), .Y(_2846_) );
AOI21X1 AOI21X1_287 ( .A(_2905_), .B(_2845_), .C(_2846_), .Y(_2847_) );
NOR3X1 NOR3X1_78 ( .A(_2887_), .B(_2888_), .C(_2889_), .Y(_2848_) );
NAND3X1 NAND3X1_432 ( .A(_2898_), .B(_2905_), .C(_2848_), .Y(_2849_) );
NAND2X1 NAND2X1_526 ( .A(_2842_), .B(_2826_), .Y(_2850_) );
AOI21X1 AOI21X1_288 ( .A(_2847_), .B(_2849_), .C(_2850_), .Y(_2851_) );
AOI22X1 AOI22X1_18 ( .A(_2839_), .B(_2840_), .C(_2831_), .D(_2912_), .Y(_2852_) );
INVX1 INVX1_390 ( .A(_2839_), .Y(_2853_) );
OAI21X1 OAI21X1_485 ( .A(micro_ucr_hash1_b_26__6_), .B(micro_ucr_hash1_a_26__6_), .C(micro_ucr_hash1_W_27__6_), .Y(_2854_) );
INVX1 INVX1_391 ( .A(micro_ucr_hash1_W_27__6_), .Y(_2855_) );
NOR2X1 NOR2X1_307 ( .A(micro_ucr_hash1_b_26__6_), .B(micro_ucr_hash1_a_26__6_), .Y(_2856_) );
NAND2X1 NAND2X1_527 ( .A(_2855_), .B(_2856_), .Y(_2857_) );
NAND2X1 NAND2X1_528 ( .A(_2854_), .B(_2857_), .Y(_2858_) );
NOR2X1 NOR2X1_308 ( .A(_2853_), .B(_2858_), .Y(_2859_) );
INVX1 INVX1_392 ( .A(_2859_), .Y(_2860_) );
NAND2X1 NAND2X1_529 ( .A(_2853_), .B(_2858_), .Y(_2861_) );
NAND2X1 NAND2X1_530 ( .A(_2861_), .B(_2860_), .Y(_2862_) );
INVX1 INVX1_393 ( .A(_2862_), .Y(_2863_) );
OAI21X1 OAI21X1_486 ( .A(_2851_), .B(_2852_), .C(_2863_), .Y(_2864_) );
NAND3X1 NAND3X1_433 ( .A(_2907_), .B(_2823_), .C(_2824_), .Y(_2865_) );
NAND2X1 NAND2X1_531 ( .A(_2865_), .B(_2831_), .Y(_2866_) );
AOI21X1 AOI21X1_289 ( .A(_2837_), .B(_2841_), .C(_2866_), .Y(_2867_) );
OAI21X1 OAI21X1_487 ( .A(_2828_), .B(_2829_), .C(_2867_), .Y(_2868_) );
INVX1 INVX1_394 ( .A(_2852_), .Y(_2869_) );
NAND3X1 NAND3X1_434 ( .A(_2869_), .B(_2862_), .C(_2868_), .Y(_2870_) );
AND2X2 AND2X2_141 ( .A(_2864_), .B(_2870_), .Y(micro_ucr_hash1_c_27__6_) );
AOI21X1 AOI21X1_290 ( .A(_2869_), .B(_2868_), .C(_2862_), .Y(_2871_) );
NOR2X1 NOR2X1_309 ( .A(micro_ucr_hash1_b_26__7_), .B(micro_ucr_hash1_a_26__7_), .Y(_2872_) );
XNOR2X1 XNOR2X1_190 ( .A(_2872_), .B(micro_ucr_hash1_W_27__7_), .Y(_2873_) );
XNOR2X1 XNOR2X1_191 ( .A(_2873_), .B(_2854_), .Y(_2874_) );
OAI21X1 OAI21X1_488 ( .A(_2871_), .B(_2859_), .C(_2874_), .Y(_2875_) );
INVX1 INVX1_395 ( .A(_2874_), .Y(_2876_) );
NAND3X1 NAND3X1_435 ( .A(_2860_), .B(_2876_), .C(_2864_), .Y(_2877_) );
NAND2X1 NAND2X1_532 ( .A(_2875_), .B(_2877_), .Y(micro_ucr_hash1_c_27__7_) );
XOR2X1 XOR2X1_261 ( .A(micro_ucr_hash1_b_28__4_), .B(gnd), .Y(micro_ucr_hash1_a_28__0_) );
XOR2X1 XOR2X1_262 ( .A(micro_ucr_hash1_b_28__5_), .B(gnd), .Y(micro_ucr_hash1_a_28__1_) );
XOR2X1 XOR2X1_263 ( .A(micro_ucr_hash1_b_28__6_), .B(gnd), .Y(micro_ucr_hash1_a_28__2_) );
XOR2X1 XOR2X1_264 ( .A(micro_ucr_hash1_b_28__7_), .B(gnd), .Y(micro_ucr_hash1_a_28__3_) );
XOR2X1 XOR2X1_265 ( .A(micro_ucr_hash1_c_27__4_), .B(micro_ucr_hash1_b_27__4_), .Y(micro_ucr_hash1_a_28__4_) );
XOR2X1 XOR2X1_266 ( .A(micro_ucr_hash1_c_27__5_), .B(micro_ucr_hash1_b_27__5_), .Y(micro_ucr_hash1_a_28__5_) );
XOR2X1 XOR2X1_267 ( .A(micro_ucr_hash1_c_27__6_), .B(micro_ucr_hash1_b_27__6_), .Y(micro_ucr_hash1_a_28__6_) );
XOR2X1 XOR2X1_268 ( .A(micro_ucr_hash1_c_27__7_), .B(micro_ucr_hash1_b_27__7_), .Y(micro_ucr_hash1_a_28__7_) );
INVX1 INVX1_396 ( .A(micro_ucr_hash1_W_28__0_), .Y(_2973_) );
NOR2X1 NOR2X1_310 ( .A(gnd), .B(micro_ucr_hash1_a_27__0_), .Y(_2974_) );
NAND2X1 NAND2X1_533 ( .A(_2973_), .B(_2974_), .Y(_2975_) );
OAI21X1 OAI21X1_489 ( .A(gnd), .B(micro_ucr_hash1_a_27__0_), .C(micro_ucr_hash1_W_28__0_), .Y(_2976_) );
NAND2X1 NAND2X1_534 ( .A(_2976_), .B(_2975_), .Y(micro_ucr_hash1_b_29__4_) );
OAI21X1 OAI21X1_490 ( .A(gnd), .B(micro_ucr_hash1_a_27__1_), .C(micro_ucr_hash1_W_28__1_), .Y(_2977_) );
INVX1 INVX1_397 ( .A(micro_ucr_hash1_W_28__1_), .Y(_2978_) );
NOR2X1 NOR2X1_311 ( .A(gnd), .B(micro_ucr_hash1_a_27__1_), .Y(_2979_) );
NAND2X1 NAND2X1_535 ( .A(_2978_), .B(_2979_), .Y(_2980_) );
NAND3X1 NAND3X1_436 ( .A(_2977_), .B(_2975_), .C(_2980_), .Y(_2981_) );
AND2X2 AND2X2_142 ( .A(_2974_), .B(_2973_), .Y(_2982_) );
INVX2 INVX2_70 ( .A(_2977_), .Y(_2983_) );
AND2X2 AND2X2_143 ( .A(_2979_), .B(_2978_), .Y(_2984_) );
OAI21X1 OAI21X1_491 ( .A(_2984_), .B(_2983_), .C(_2982_), .Y(_2985_) );
AND2X2 AND2X2_144 ( .A(_2985_), .B(_2981_), .Y(micro_ucr_hash1_b_29__5_) );
OAI21X1 OAI21X1_492 ( .A(gnd), .B(micro_ucr_hash1_a_27__2_), .C(micro_ucr_hash1_W_28__2_), .Y(_2986_) );
INVX1 INVX1_398 ( .A(micro_ucr_hash1_W_28__2_), .Y(_2987_) );
NOR2X1 NOR2X1_312 ( .A(gnd), .B(micro_ucr_hash1_a_27__2_), .Y(_2988_) );
NAND2X1 NAND2X1_536 ( .A(_2987_), .B(_2988_), .Y(_2989_) );
NAND2X1 NAND2X1_537 ( .A(_2986_), .B(_2989_), .Y(_2990_) );
NAND3X1 NAND3X1_437 ( .A(_2986_), .B(_2989_), .C(_2983_), .Y(_2991_) );
OAI21X1 OAI21X1_493 ( .A(_2981_), .B(_2990_), .C(_2991_), .Y(_2992_) );
INVX1 INVX1_399 ( .A(_2990_), .Y(_2993_) );
OAI21X1 OAI21X1_494 ( .A(_2982_), .B(_2984_), .C(_2977_), .Y(_2994_) );
NOR2X1 NOR2X1_313 ( .A(_2994_), .B(_2993_), .Y(_2995_) );
NOR2X1 NOR2X1_314 ( .A(_2992_), .B(_2995_), .Y(micro_ucr_hash1_b_29__6_) );
INVX1 INVX1_400 ( .A(micro_ucr_hash1_W_28__3_), .Y(_2996_) );
OAI21X1 OAI21X1_495 ( .A(gnd), .B(micro_ucr_hash1_a_27__3_), .C(_2996_), .Y(_2997_) );
NOR2X1 NOR2X1_315 ( .A(gnd), .B(micro_ucr_hash1_a_27__3_), .Y(_2998_) );
NAND2X1 NAND2X1_538 ( .A(micro_ucr_hash1_W_28__3_), .B(_2998_), .Y(_2999_) );
NAND3X1 NAND3X1_438 ( .A(_2986_), .B(_2997_), .C(_2999_), .Y(_3000_) );
INVX1 INVX1_401 ( .A(_2986_), .Y(_3001_) );
OAI21X1 OAI21X1_496 ( .A(gnd), .B(micro_ucr_hash1_a_27__3_), .C(micro_ucr_hash1_W_28__3_), .Y(_3002_) );
NAND2X1 NAND2X1_539 ( .A(_2996_), .B(_2998_), .Y(_3003_) );
NAND3X1 NAND3X1_439 ( .A(_3002_), .B(_3003_), .C(_3001_), .Y(_3004_) );
NAND2X1 NAND2X1_540 ( .A(_3000_), .B(_3004_), .Y(_3005_) );
XNOR2X1 XNOR2X1_192 ( .A(_2992_), .B(_3005_), .Y(micro_ucr_hash1_b_29__7_) );
INVX1 INVX1_402 ( .A(_3002_), .Y(_3006_) );
OAI21X1 OAI21X1_497 ( .A(micro_ucr_hash1_b_27__4_), .B(micro_ucr_hash1_a_27__4_), .C(micro_ucr_hash1_W_28__4_), .Y(_3007_) );
INVX1 INVX1_403 ( .A(micro_ucr_hash1_b_27__4_), .Y(_3008_) );
INVX1 INVX1_404 ( .A(micro_ucr_hash1_a_27__4_), .Y(_3009_) );
INVX1 INVX1_405 ( .A(micro_ucr_hash1_W_28__4_), .Y(_3010_) );
NAND3X1 NAND3X1_440 ( .A(_3008_), .B(_3009_), .C(_3010_), .Y(_3011_) );
AOI21X1 AOI21X1_291 ( .A(_3007_), .B(_3011_), .C(_3006_), .Y(_2917_) );
OAI21X1 OAI21X1_498 ( .A(micro_ucr_hash1_b_27__4_), .B(micro_ucr_hash1_a_27__4_), .C(_3010_), .Y(_2918_) );
NAND3X1 NAND3X1_441 ( .A(micro_ucr_hash1_W_28__4_), .B(_3008_), .C(_3009_), .Y(_2919_) );
AOI21X1 AOI21X1_292 ( .A(_2918_), .B(_2919_), .C(_3002_), .Y(_2920_) );
NOR2X1 NOR2X1_316 ( .A(_2920_), .B(_2917_), .Y(_2921_) );
AOI21X1 AOI21X1_293 ( .A(_3002_), .B(_3003_), .C(_3001_), .Y(_2922_) );
OAI21X1 OAI21X1_499 ( .A(_2922_), .B(_2991_), .C(_3004_), .Y(_2923_) );
NOR3X1 NOR3X1_79 ( .A(_2981_), .B(_2990_), .C(_2922_), .Y(_2924_) );
NOR2X1 NOR2X1_317 ( .A(_2923_), .B(_2924_), .Y(_2925_) );
XNOR2X1 XNOR2X1_193 ( .A(_2925_), .B(_2921_), .Y(micro_ucr_hash1_c_28__4_) );
NAND3X1 NAND3X1_442 ( .A(_3007_), .B(_3011_), .C(_3006_), .Y(_2926_) );
OAI21X1 OAI21X1_500 ( .A(_2925_), .B(_2917_), .C(_2926_), .Y(_2927_) );
INVX1 INVX1_406 ( .A(micro_ucr_hash1_W_28__5_), .Y(_2928_) );
OAI21X1 OAI21X1_501 ( .A(micro_ucr_hash1_b_27__5_), .B(micro_ucr_hash1_a_27__5_), .C(_2928_), .Y(_2929_) );
NOR2X1 NOR2X1_318 ( .A(micro_ucr_hash1_b_27__5_), .B(micro_ucr_hash1_a_27__5_), .Y(_2930_) );
NAND2X1 NAND2X1_541 ( .A(micro_ucr_hash1_W_28__5_), .B(_2930_), .Y(_2931_) );
NAND3X1 NAND3X1_443 ( .A(_3007_), .B(_2929_), .C(_2931_), .Y(_2932_) );
INVX1 INVX1_407 ( .A(_3007_), .Y(_2933_) );
NAND2X1 NAND2X1_542 ( .A(_2928_), .B(_2930_), .Y(_2934_) );
OAI21X1 OAI21X1_502 ( .A(micro_ucr_hash1_b_27__5_), .B(micro_ucr_hash1_a_27__5_), .C(micro_ucr_hash1_W_28__5_), .Y(_2935_) );
NAND3X1 NAND3X1_444 ( .A(_2935_), .B(_2934_), .C(_2933_), .Y(_2936_) );
NAND2X1 NAND2X1_543 ( .A(_2932_), .B(_2936_), .Y(_2937_) );
XOR2X1 XOR2X1_269 ( .A(_2927_), .B(_2937_), .Y(micro_ucr_hash1_c_28__5_) );
OAI21X1 OAI21X1_503 ( .A(gnd), .B(micro_ucr_hash1_a_27__2_), .C(_2987_), .Y(_2938_) );
NAND2X1 NAND2X1_544 ( .A(micro_ucr_hash1_W_28__2_), .B(_2988_), .Y(_2939_) );
AOI21X1 AOI21X1_294 ( .A(_2938_), .B(_2939_), .C(_2977_), .Y(_2940_) );
INVX1 INVX1_408 ( .A(_3004_), .Y(_2941_) );
AOI21X1 AOI21X1_295 ( .A(_3000_), .B(_2940_), .C(_2941_), .Y(_2942_) );
NOR3X1 NOR3X1_80 ( .A(_2982_), .B(_2983_), .C(_2984_), .Y(_2943_) );
NAND3X1 NAND3X1_445 ( .A(_2993_), .B(_3000_), .C(_2943_), .Y(_2944_) );
NAND2X1 NAND2X1_545 ( .A(_2937_), .B(_2921_), .Y(_2945_) );
AOI21X1 AOI21X1_296 ( .A(_2942_), .B(_2944_), .C(_2945_), .Y(_2946_) );
AOI22X1 AOI22X1_19 ( .A(_2934_), .B(_2935_), .C(_2926_), .D(_3007_), .Y(_2947_) );
INVX1 INVX1_409 ( .A(_2934_), .Y(_2948_) );
OAI21X1 OAI21X1_504 ( .A(micro_ucr_hash1_b_27__6_), .B(micro_ucr_hash1_a_27__6_), .C(micro_ucr_hash1_W_28__6_), .Y(_2949_) );
INVX1 INVX1_410 ( .A(micro_ucr_hash1_W_28__6_), .Y(_2950_) );
NOR2X1 NOR2X1_319 ( .A(micro_ucr_hash1_b_27__6_), .B(micro_ucr_hash1_a_27__6_), .Y(_2951_) );
NAND2X1 NAND2X1_546 ( .A(_2950_), .B(_2951_), .Y(_2952_) );
NAND2X1 NAND2X1_547 ( .A(_2949_), .B(_2952_), .Y(_2953_) );
NOR2X1 NOR2X1_320 ( .A(_2948_), .B(_2953_), .Y(_2954_) );
INVX1 INVX1_411 ( .A(_2954_), .Y(_2955_) );
NAND2X1 NAND2X1_548 ( .A(_2948_), .B(_2953_), .Y(_2956_) );
NAND2X1 NAND2X1_549 ( .A(_2956_), .B(_2955_), .Y(_2957_) );
INVX1 INVX1_412 ( .A(_2957_), .Y(_2958_) );
OAI21X1 OAI21X1_505 ( .A(_2946_), .B(_2947_), .C(_2958_), .Y(_2959_) );
NAND3X1 NAND3X1_446 ( .A(_3002_), .B(_2918_), .C(_2919_), .Y(_2960_) );
NAND2X1 NAND2X1_550 ( .A(_2960_), .B(_2926_), .Y(_2961_) );
AOI21X1 AOI21X1_297 ( .A(_2932_), .B(_2936_), .C(_2961_), .Y(_2962_) );
OAI21X1 OAI21X1_506 ( .A(_2923_), .B(_2924_), .C(_2962_), .Y(_2963_) );
INVX1 INVX1_413 ( .A(_2947_), .Y(_2964_) );
NAND3X1 NAND3X1_447 ( .A(_2964_), .B(_2957_), .C(_2963_), .Y(_2965_) );
AND2X2 AND2X2_145 ( .A(_2959_), .B(_2965_), .Y(micro_ucr_hash1_c_28__6_) );
AOI21X1 AOI21X1_298 ( .A(_2964_), .B(_2963_), .C(_2957_), .Y(_2966_) );
NOR2X1 NOR2X1_321 ( .A(micro_ucr_hash1_b_27__7_), .B(micro_ucr_hash1_a_27__7_), .Y(_2967_) );
XNOR2X1 XNOR2X1_194 ( .A(_2967_), .B(micro_ucr_hash1_W_28__7_), .Y(_2968_) );
XNOR2X1 XNOR2X1_195 ( .A(_2968_), .B(_2949_), .Y(_2969_) );
OAI21X1 OAI21X1_507 ( .A(_2966_), .B(_2954_), .C(_2969_), .Y(_2970_) );
INVX1 INVX1_414 ( .A(_2969_), .Y(_2971_) );
NAND3X1 NAND3X1_448 ( .A(_2955_), .B(_2971_), .C(_2959_), .Y(_2972_) );
NAND2X1 NAND2X1_551 ( .A(_2970_), .B(_2972_), .Y(micro_ucr_hash1_c_28__7_) );
XOR2X1 XOR2X1_270 ( .A(micro_ucr_hash1_b_29__4_), .B(gnd), .Y(micro_ucr_hash1_a_29__0_) );
XOR2X1 XOR2X1_271 ( .A(micro_ucr_hash1_b_29__5_), .B(gnd), .Y(micro_ucr_hash1_a_29__1_) );
XOR2X1 XOR2X1_272 ( .A(micro_ucr_hash1_b_29__6_), .B(gnd), .Y(micro_ucr_hash1_a_29__2_) );
XOR2X1 XOR2X1_273 ( .A(micro_ucr_hash1_b_29__7_), .B(gnd), .Y(micro_ucr_hash1_a_29__3_) );
XOR2X1 XOR2X1_274 ( .A(micro_ucr_hash1_c_28__4_), .B(micro_ucr_hash1_b_28__4_), .Y(micro_ucr_hash1_a_29__4_) );
XOR2X1 XOR2X1_275 ( .A(micro_ucr_hash1_c_28__5_), .B(micro_ucr_hash1_b_28__5_), .Y(micro_ucr_hash1_a_29__5_) );
XOR2X1 XOR2X1_276 ( .A(micro_ucr_hash1_c_28__6_), .B(micro_ucr_hash1_b_28__6_), .Y(micro_ucr_hash1_a_29__6_) );
XOR2X1 XOR2X1_277 ( .A(micro_ucr_hash1_c_28__7_), .B(micro_ucr_hash1_b_28__7_), .Y(micro_ucr_hash1_a_29__7_) );
INVX1 INVX1_415 ( .A(micro_ucr_hash1_W_29__0_), .Y(_3068_) );
NOR2X1 NOR2X1_322 ( .A(gnd), .B(micro_ucr_hash1_a_28__0_), .Y(_3069_) );
NAND2X1 NAND2X1_552 ( .A(_3068_), .B(_3069_), .Y(_3070_) );
OAI21X1 OAI21X1_508 ( .A(gnd), .B(micro_ucr_hash1_a_28__0_), .C(micro_ucr_hash1_W_29__0_), .Y(_3071_) );
NAND2X1 NAND2X1_553 ( .A(_3071_), .B(_3070_), .Y(micro_ucr_hash1_b_30__4_) );
OAI21X1 OAI21X1_509 ( .A(gnd), .B(micro_ucr_hash1_a_28__1_), .C(micro_ucr_hash1_W_29__1_), .Y(_3072_) );
INVX1 INVX1_416 ( .A(micro_ucr_hash1_W_29__1_), .Y(_3073_) );
NOR2X1 NOR2X1_323 ( .A(gnd), .B(micro_ucr_hash1_a_28__1_), .Y(_3074_) );
NAND2X1 NAND2X1_554 ( .A(_3073_), .B(_3074_), .Y(_3075_) );
NAND3X1 NAND3X1_449 ( .A(_3072_), .B(_3070_), .C(_3075_), .Y(_3076_) );
AND2X2 AND2X2_146 ( .A(_3069_), .B(_3068_), .Y(_3077_) );
INVX2 INVX2_71 ( .A(_3072_), .Y(_3078_) );
AND2X2 AND2X2_147 ( .A(_3074_), .B(_3073_), .Y(_3079_) );
OAI21X1 OAI21X1_510 ( .A(_3079_), .B(_3078_), .C(_3077_), .Y(_3080_) );
AND2X2 AND2X2_148 ( .A(_3080_), .B(_3076_), .Y(micro_ucr_hash1_b_30__5_) );
OAI21X1 OAI21X1_511 ( .A(gnd), .B(micro_ucr_hash1_a_28__2_), .C(micro_ucr_hash1_W_29__2_), .Y(_3081_) );
INVX1 INVX1_417 ( .A(micro_ucr_hash1_W_29__2_), .Y(_3082_) );
NOR2X1 NOR2X1_324 ( .A(gnd), .B(micro_ucr_hash1_a_28__2_), .Y(_3083_) );
NAND2X1 NAND2X1_555 ( .A(_3082_), .B(_3083_), .Y(_3084_) );
NAND2X1 NAND2X1_556 ( .A(_3081_), .B(_3084_), .Y(_3085_) );
NAND3X1 NAND3X1_450 ( .A(_3081_), .B(_3084_), .C(_3078_), .Y(_3086_) );
OAI21X1 OAI21X1_512 ( .A(_3076_), .B(_3085_), .C(_3086_), .Y(_3087_) );
INVX1 INVX1_418 ( .A(_3085_), .Y(_3088_) );
OAI21X1 OAI21X1_513 ( .A(_3077_), .B(_3079_), .C(_3072_), .Y(_3089_) );
NOR2X1 NOR2X1_325 ( .A(_3089_), .B(_3088_), .Y(_3090_) );
NOR2X1 NOR2X1_326 ( .A(_3087_), .B(_3090_), .Y(micro_ucr_hash1_b_30__6_) );
INVX1 INVX1_419 ( .A(micro_ucr_hash1_W_29__3_), .Y(_3091_) );
OAI21X1 OAI21X1_514 ( .A(gnd), .B(micro_ucr_hash1_a_28__3_), .C(_3091_), .Y(_3092_) );
NOR2X1 NOR2X1_327 ( .A(gnd), .B(micro_ucr_hash1_a_28__3_), .Y(_3093_) );
NAND2X1 NAND2X1_557 ( .A(micro_ucr_hash1_W_29__3_), .B(_3093_), .Y(_3094_) );
NAND3X1 NAND3X1_451 ( .A(_3081_), .B(_3092_), .C(_3094_), .Y(_3095_) );
INVX1 INVX1_420 ( .A(_3081_), .Y(_3096_) );
OAI21X1 OAI21X1_515 ( .A(gnd), .B(micro_ucr_hash1_a_28__3_), .C(micro_ucr_hash1_W_29__3_), .Y(_3097_) );
NAND2X1 NAND2X1_558 ( .A(_3091_), .B(_3093_), .Y(_3098_) );
NAND3X1 NAND3X1_452 ( .A(_3097_), .B(_3098_), .C(_3096_), .Y(_3099_) );
NAND2X1 NAND2X1_559 ( .A(_3095_), .B(_3099_), .Y(_3100_) );
XNOR2X1 XNOR2X1_196 ( .A(_3087_), .B(_3100_), .Y(micro_ucr_hash1_b_30__7_) );
INVX1 INVX1_421 ( .A(_3097_), .Y(_3101_) );
OAI21X1 OAI21X1_516 ( .A(micro_ucr_hash1_b_28__4_), .B(micro_ucr_hash1_a_28__4_), .C(micro_ucr_hash1_W_29__4_), .Y(_3102_) );
INVX1 INVX1_422 ( .A(micro_ucr_hash1_b_28__4_), .Y(_3103_) );
INVX1 INVX1_423 ( .A(micro_ucr_hash1_a_28__4_), .Y(_3104_) );
INVX1 INVX1_424 ( .A(micro_ucr_hash1_W_29__4_), .Y(_3105_) );
NAND3X1 NAND3X1_453 ( .A(_3103_), .B(_3104_), .C(_3105_), .Y(_3106_) );
AOI21X1 AOI21X1_299 ( .A(_3102_), .B(_3106_), .C(_3101_), .Y(_3012_) );
OAI21X1 OAI21X1_517 ( .A(micro_ucr_hash1_b_28__4_), .B(micro_ucr_hash1_a_28__4_), .C(_3105_), .Y(_3013_) );
NAND3X1 NAND3X1_454 ( .A(micro_ucr_hash1_W_29__4_), .B(_3103_), .C(_3104_), .Y(_3014_) );
AOI21X1 AOI21X1_300 ( .A(_3013_), .B(_3014_), .C(_3097_), .Y(_3015_) );
NOR2X1 NOR2X1_328 ( .A(_3015_), .B(_3012_), .Y(_3016_) );
AOI21X1 AOI21X1_301 ( .A(_3097_), .B(_3098_), .C(_3096_), .Y(_3017_) );
OAI21X1 OAI21X1_518 ( .A(_3017_), .B(_3086_), .C(_3099_), .Y(_3018_) );
NOR3X1 NOR3X1_81 ( .A(_3076_), .B(_3085_), .C(_3017_), .Y(_3019_) );
NOR2X1 NOR2X1_329 ( .A(_3018_), .B(_3019_), .Y(_3020_) );
XNOR2X1 XNOR2X1_197 ( .A(_3020_), .B(_3016_), .Y(micro_ucr_hash1_c_29__4_) );
NAND3X1 NAND3X1_455 ( .A(_3102_), .B(_3106_), .C(_3101_), .Y(_3021_) );
OAI21X1 OAI21X1_519 ( .A(_3020_), .B(_3012_), .C(_3021_), .Y(_3022_) );
INVX1 INVX1_425 ( .A(micro_ucr_hash1_W_29__5_), .Y(_3023_) );
OAI21X1 OAI21X1_520 ( .A(micro_ucr_hash1_b_28__5_), .B(micro_ucr_hash1_a_28__5_), .C(_3023_), .Y(_3024_) );
NOR2X1 NOR2X1_330 ( .A(micro_ucr_hash1_b_28__5_), .B(micro_ucr_hash1_a_28__5_), .Y(_3025_) );
NAND2X1 NAND2X1_560 ( .A(micro_ucr_hash1_W_29__5_), .B(_3025_), .Y(_3026_) );
NAND3X1 NAND3X1_456 ( .A(_3102_), .B(_3024_), .C(_3026_), .Y(_3027_) );
INVX1 INVX1_426 ( .A(_3102_), .Y(_3028_) );
NAND2X1 NAND2X1_561 ( .A(_3023_), .B(_3025_), .Y(_3029_) );
OAI21X1 OAI21X1_521 ( .A(micro_ucr_hash1_b_28__5_), .B(micro_ucr_hash1_a_28__5_), .C(micro_ucr_hash1_W_29__5_), .Y(_3030_) );
NAND3X1 NAND3X1_457 ( .A(_3030_), .B(_3029_), .C(_3028_), .Y(_3031_) );
NAND2X1 NAND2X1_562 ( .A(_3027_), .B(_3031_), .Y(_3032_) );
XOR2X1 XOR2X1_278 ( .A(_3022_), .B(_3032_), .Y(micro_ucr_hash1_c_29__5_) );
OAI21X1 OAI21X1_522 ( .A(gnd), .B(micro_ucr_hash1_a_28__2_), .C(_3082_), .Y(_3033_) );
NAND2X1 NAND2X1_563 ( .A(micro_ucr_hash1_W_29__2_), .B(_3083_), .Y(_3034_) );
AOI21X1 AOI21X1_302 ( .A(_3033_), .B(_3034_), .C(_3072_), .Y(_3035_) );
INVX1 INVX1_427 ( .A(_3099_), .Y(_3036_) );
AOI21X1 AOI21X1_303 ( .A(_3095_), .B(_3035_), .C(_3036_), .Y(_3037_) );
NOR3X1 NOR3X1_82 ( .A(_3077_), .B(_3078_), .C(_3079_), .Y(_3038_) );
NAND3X1 NAND3X1_458 ( .A(_3088_), .B(_3095_), .C(_3038_), .Y(_3039_) );
NAND2X1 NAND2X1_564 ( .A(_3032_), .B(_3016_), .Y(_3040_) );
AOI21X1 AOI21X1_304 ( .A(_3037_), .B(_3039_), .C(_3040_), .Y(_3041_) );
AOI22X1 AOI22X1_20 ( .A(_3029_), .B(_3030_), .C(_3021_), .D(_3102_), .Y(_3042_) );
INVX1 INVX1_428 ( .A(_3029_), .Y(_3043_) );
OAI21X1 OAI21X1_523 ( .A(micro_ucr_hash1_b_28__6_), .B(micro_ucr_hash1_a_28__6_), .C(micro_ucr_hash1_W_29__6_), .Y(_3044_) );
INVX1 INVX1_429 ( .A(micro_ucr_hash1_W_29__6_), .Y(_3045_) );
NOR2X1 NOR2X1_331 ( .A(micro_ucr_hash1_b_28__6_), .B(micro_ucr_hash1_a_28__6_), .Y(_3046_) );
NAND2X1 NAND2X1_565 ( .A(_3045_), .B(_3046_), .Y(_3047_) );
NAND2X1 NAND2X1_566 ( .A(_3044_), .B(_3047_), .Y(_3048_) );
NOR2X1 NOR2X1_332 ( .A(_3043_), .B(_3048_), .Y(_3049_) );
INVX1 INVX1_430 ( .A(_3049_), .Y(_3050_) );
NAND2X1 NAND2X1_567 ( .A(_3043_), .B(_3048_), .Y(_3051_) );
NAND2X1 NAND2X1_568 ( .A(_3051_), .B(_3050_), .Y(_3052_) );
INVX1 INVX1_431 ( .A(_3052_), .Y(_3053_) );
OAI21X1 OAI21X1_524 ( .A(_3041_), .B(_3042_), .C(_3053_), .Y(_3054_) );
NAND3X1 NAND3X1_459 ( .A(_3097_), .B(_3013_), .C(_3014_), .Y(_3055_) );
NAND2X1 NAND2X1_569 ( .A(_3055_), .B(_3021_), .Y(_3056_) );
AOI21X1 AOI21X1_305 ( .A(_3027_), .B(_3031_), .C(_3056_), .Y(_3057_) );
OAI21X1 OAI21X1_525 ( .A(_3018_), .B(_3019_), .C(_3057_), .Y(_3058_) );
INVX1 INVX1_432 ( .A(_3042_), .Y(_3059_) );
NAND3X1 NAND3X1_460 ( .A(_3059_), .B(_3052_), .C(_3058_), .Y(_3060_) );
AND2X2 AND2X2_149 ( .A(_3054_), .B(_3060_), .Y(micro_ucr_hash1_c_29__6_) );
AOI21X1 AOI21X1_306 ( .A(_3059_), .B(_3058_), .C(_3052_), .Y(_3061_) );
NOR2X1 NOR2X1_333 ( .A(micro_ucr_hash1_b_28__7_), .B(micro_ucr_hash1_a_28__7_), .Y(_3062_) );
XNOR2X1 XNOR2X1_198 ( .A(_3062_), .B(micro_ucr_hash1_W_29__7_), .Y(_3063_) );
XNOR2X1 XNOR2X1_199 ( .A(_3063_), .B(_3044_), .Y(_3064_) );
OAI21X1 OAI21X1_526 ( .A(_3061_), .B(_3049_), .C(_3064_), .Y(_3065_) );
INVX1 INVX1_433 ( .A(_3064_), .Y(_3066_) );
NAND3X1 NAND3X1_461 ( .A(_3050_), .B(_3066_), .C(_3054_), .Y(_3067_) );
NAND2X1 NAND2X1_570 ( .A(_3065_), .B(_3067_), .Y(micro_ucr_hash1_c_29__7_) );
XOR2X1 XOR2X1_279 ( .A(micro_ucr_hash1_b_30__4_), .B(gnd), .Y(micro_ucr_hash1_a_30__0_) );
XOR2X1 XOR2X1_280 ( .A(micro_ucr_hash1_b_30__5_), .B(gnd), .Y(micro_ucr_hash1_a_30__1_) );
XOR2X1 XOR2X1_281 ( .A(micro_ucr_hash1_b_30__6_), .B(gnd), .Y(micro_ucr_hash1_a_30__2_) );
XOR2X1 XOR2X1_282 ( .A(micro_ucr_hash1_b_30__7_), .B(gnd), .Y(micro_ucr_hash1_a_30__3_) );
XOR2X1 XOR2X1_283 ( .A(micro_ucr_hash1_c_29__4_), .B(micro_ucr_hash1_b_29__4_), .Y(micro_ucr_hash1_a_30__4_) );
XOR2X1 XOR2X1_284 ( .A(micro_ucr_hash1_c_29__5_), .B(micro_ucr_hash1_b_29__5_), .Y(micro_ucr_hash1_a_30__5_) );
XOR2X1 XOR2X1_285 ( .A(micro_ucr_hash1_c_29__6_), .B(micro_ucr_hash1_b_29__6_), .Y(micro_ucr_hash1_a_30__6_) );
XOR2X1 XOR2X1_286 ( .A(micro_ucr_hash1_c_29__7_), .B(micro_ucr_hash1_b_29__7_), .Y(micro_ucr_hash1_a_30__7_) );
INVX1 INVX1_434 ( .A(micro_ucr_hash1_W_30__0_), .Y(_3163_) );
NOR2X1 NOR2X1_334 ( .A(gnd), .B(micro_ucr_hash1_a_29__0_), .Y(_3164_) );
NAND2X1 NAND2X1_571 ( .A(_3163_), .B(_3164_), .Y(_3165_) );
OAI21X1 OAI21X1_527 ( .A(gnd), .B(micro_ucr_hash1_a_29__0_), .C(micro_ucr_hash1_W_30__0_), .Y(_3166_) );
NAND2X1 NAND2X1_572 ( .A(_3166_), .B(_3165_), .Y(micro_ucr_hash1_b_31__4_) );
OAI21X1 OAI21X1_528 ( .A(gnd), .B(micro_ucr_hash1_a_29__1_), .C(micro_ucr_hash1_W_30__1_), .Y(_3167_) );
INVX1 INVX1_435 ( .A(micro_ucr_hash1_W_30__1_), .Y(_3168_) );
NOR2X1 NOR2X1_335 ( .A(gnd), .B(micro_ucr_hash1_a_29__1_), .Y(_3169_) );
NAND2X1 NAND2X1_573 ( .A(_3168_), .B(_3169_), .Y(_3170_) );
NAND3X1 NAND3X1_462 ( .A(_3167_), .B(_3165_), .C(_3170_), .Y(_3171_) );
AND2X2 AND2X2_150 ( .A(_3164_), .B(_3163_), .Y(_3172_) );
INVX2 INVX2_72 ( .A(_3167_), .Y(_3173_) );
AND2X2 AND2X2_151 ( .A(_3169_), .B(_3168_), .Y(_3174_) );
OAI21X1 OAI21X1_529 ( .A(_3174_), .B(_3173_), .C(_3172_), .Y(_3175_) );
AND2X2 AND2X2_152 ( .A(_3175_), .B(_3171_), .Y(micro_ucr_hash1_b_31__5_) );
OAI21X1 OAI21X1_530 ( .A(gnd), .B(micro_ucr_hash1_a_29__2_), .C(micro_ucr_hash1_W_30__2_), .Y(_3176_) );
INVX1 INVX1_436 ( .A(micro_ucr_hash1_W_30__2_), .Y(_3177_) );
NOR2X1 NOR2X1_336 ( .A(gnd), .B(micro_ucr_hash1_a_29__2_), .Y(_3178_) );
NAND2X1 NAND2X1_574 ( .A(_3177_), .B(_3178_), .Y(_3179_) );
NAND2X1 NAND2X1_575 ( .A(_3176_), .B(_3179_), .Y(_3180_) );
NAND3X1 NAND3X1_463 ( .A(_3176_), .B(_3179_), .C(_3173_), .Y(_3181_) );
OAI21X1 OAI21X1_531 ( .A(_3171_), .B(_3180_), .C(_3181_), .Y(_3182_) );
INVX1 INVX1_437 ( .A(_3180_), .Y(_3183_) );
OAI21X1 OAI21X1_532 ( .A(_3172_), .B(_3174_), .C(_3167_), .Y(_3184_) );
NOR2X1 NOR2X1_337 ( .A(_3184_), .B(_3183_), .Y(_3185_) );
NOR2X1 NOR2X1_338 ( .A(_3182_), .B(_3185_), .Y(micro_ucr_hash1_b_31__6_) );
INVX1 INVX1_438 ( .A(micro_ucr_hash1_W_30__3_), .Y(_3186_) );
OAI21X1 OAI21X1_533 ( .A(gnd), .B(micro_ucr_hash1_a_29__3_), .C(_3186_), .Y(_3187_) );
NOR2X1 NOR2X1_339 ( .A(gnd), .B(micro_ucr_hash1_a_29__3_), .Y(_3188_) );
NAND2X1 NAND2X1_576 ( .A(micro_ucr_hash1_W_30__3_), .B(_3188_), .Y(_3189_) );
NAND3X1 NAND3X1_464 ( .A(_3176_), .B(_3187_), .C(_3189_), .Y(_3190_) );
INVX1 INVX1_439 ( .A(_3176_), .Y(_3191_) );
OAI21X1 OAI21X1_534 ( .A(gnd), .B(micro_ucr_hash1_a_29__3_), .C(micro_ucr_hash1_W_30__3_), .Y(_3192_) );
NAND2X1 NAND2X1_577 ( .A(_3186_), .B(_3188_), .Y(_3193_) );
NAND3X1 NAND3X1_465 ( .A(_3192_), .B(_3193_), .C(_3191_), .Y(_3194_) );
NAND2X1 NAND2X1_578 ( .A(_3190_), .B(_3194_), .Y(_3195_) );
XNOR2X1 XNOR2X1_200 ( .A(_3182_), .B(_3195_), .Y(micro_ucr_hash1_b_31__7_) );
INVX1 INVX1_440 ( .A(_3192_), .Y(_3196_) );
OAI21X1 OAI21X1_535 ( .A(micro_ucr_hash1_b_29__4_), .B(micro_ucr_hash1_a_29__4_), .C(micro_ucr_hash1_W_30__4_), .Y(_3197_) );
INVX1 INVX1_441 ( .A(micro_ucr_hash1_b_29__4_), .Y(_3198_) );
INVX1 INVX1_442 ( .A(micro_ucr_hash1_a_29__4_), .Y(_3199_) );
INVX1 INVX1_443 ( .A(micro_ucr_hash1_W_30__4_), .Y(_3200_) );
NAND3X1 NAND3X1_466 ( .A(_3198_), .B(_3199_), .C(_3200_), .Y(_3201_) );
AOI21X1 AOI21X1_307 ( .A(_3197_), .B(_3201_), .C(_3196_), .Y(_3107_) );
OAI21X1 OAI21X1_536 ( .A(micro_ucr_hash1_b_29__4_), .B(micro_ucr_hash1_a_29__4_), .C(_3200_), .Y(_3108_) );
NAND3X1 NAND3X1_467 ( .A(micro_ucr_hash1_W_30__4_), .B(_3198_), .C(_3199_), .Y(_3109_) );
AOI21X1 AOI21X1_308 ( .A(_3108_), .B(_3109_), .C(_3192_), .Y(_3110_) );
NOR2X1 NOR2X1_340 ( .A(_3110_), .B(_3107_), .Y(_3111_) );
AOI21X1 AOI21X1_309 ( .A(_3192_), .B(_3193_), .C(_3191_), .Y(_3112_) );
OAI21X1 OAI21X1_537 ( .A(_3112_), .B(_3181_), .C(_3194_), .Y(_3113_) );
NOR3X1 NOR3X1_83 ( .A(_3171_), .B(_3180_), .C(_3112_), .Y(_3114_) );
NOR2X1 NOR2X1_341 ( .A(_3113_), .B(_3114_), .Y(_3115_) );
XNOR2X1 XNOR2X1_201 ( .A(_3115_), .B(_3111_), .Y(micro_ucr_hash1_c_30__4_) );
NAND3X1 NAND3X1_468 ( .A(_3197_), .B(_3201_), .C(_3196_), .Y(_3116_) );
OAI21X1 OAI21X1_538 ( .A(_3115_), .B(_3107_), .C(_3116_), .Y(_3117_) );
INVX1 INVX1_444 ( .A(micro_ucr_hash1_W_30__5_), .Y(_3118_) );
OAI21X1 OAI21X1_539 ( .A(micro_ucr_hash1_b_29__5_), .B(micro_ucr_hash1_a_29__5_), .C(_3118_), .Y(_3119_) );
NOR2X1 NOR2X1_342 ( .A(micro_ucr_hash1_b_29__5_), .B(micro_ucr_hash1_a_29__5_), .Y(_3120_) );
NAND2X1 NAND2X1_579 ( .A(micro_ucr_hash1_W_30__5_), .B(_3120_), .Y(_3121_) );
NAND3X1 NAND3X1_469 ( .A(_3197_), .B(_3119_), .C(_3121_), .Y(_3122_) );
INVX1 INVX1_445 ( .A(_3197_), .Y(_3123_) );
NAND2X1 NAND2X1_580 ( .A(_3118_), .B(_3120_), .Y(_3124_) );
OAI21X1 OAI21X1_540 ( .A(micro_ucr_hash1_b_29__5_), .B(micro_ucr_hash1_a_29__5_), .C(micro_ucr_hash1_W_30__5_), .Y(_3125_) );
NAND3X1 NAND3X1_470 ( .A(_3125_), .B(_3124_), .C(_3123_), .Y(_3126_) );
NAND2X1 NAND2X1_581 ( .A(_3122_), .B(_3126_), .Y(_3127_) );
XOR2X1 XOR2X1_287 ( .A(_3117_), .B(_3127_), .Y(micro_ucr_hash1_c_30__5_) );
OAI21X1 OAI21X1_541 ( .A(gnd), .B(micro_ucr_hash1_a_29__2_), .C(_3177_), .Y(_3128_) );
NAND2X1 NAND2X1_582 ( .A(micro_ucr_hash1_W_30__2_), .B(_3178_), .Y(_3129_) );
AOI21X1 AOI21X1_310 ( .A(_3128_), .B(_3129_), .C(_3167_), .Y(_3130_) );
INVX1 INVX1_446 ( .A(_3194_), .Y(_3131_) );
AOI21X1 AOI21X1_311 ( .A(_3190_), .B(_3130_), .C(_3131_), .Y(_3132_) );
NOR3X1 NOR3X1_84 ( .A(_3172_), .B(_3173_), .C(_3174_), .Y(_3133_) );
NAND3X1 NAND3X1_471 ( .A(_3183_), .B(_3190_), .C(_3133_), .Y(_3134_) );
NAND2X1 NAND2X1_583 ( .A(_3127_), .B(_3111_), .Y(_3135_) );
AOI21X1 AOI21X1_312 ( .A(_3132_), .B(_3134_), .C(_3135_), .Y(_3136_) );
AOI22X1 AOI22X1_21 ( .A(_3124_), .B(_3125_), .C(_3116_), .D(_3197_), .Y(_3137_) );
INVX1 INVX1_447 ( .A(_3124_), .Y(_3138_) );
OAI21X1 OAI21X1_542 ( .A(micro_ucr_hash1_b_29__6_), .B(micro_ucr_hash1_a_29__6_), .C(micro_ucr_hash1_W_30__6_), .Y(_3139_) );
INVX1 INVX1_448 ( .A(micro_ucr_hash1_W_30__6_), .Y(_3140_) );
NOR2X1 NOR2X1_343 ( .A(micro_ucr_hash1_b_29__6_), .B(micro_ucr_hash1_a_29__6_), .Y(_3141_) );
NAND2X1 NAND2X1_584 ( .A(_3140_), .B(_3141_), .Y(_3142_) );
NAND2X1 NAND2X1_585 ( .A(_3139_), .B(_3142_), .Y(_3143_) );
NOR2X1 NOR2X1_344 ( .A(_3138_), .B(_3143_), .Y(_3144_) );
INVX1 INVX1_449 ( .A(_3144_), .Y(_3145_) );
NAND2X1 NAND2X1_586 ( .A(_3138_), .B(_3143_), .Y(_3146_) );
NAND2X1 NAND2X1_587 ( .A(_3146_), .B(_3145_), .Y(_3147_) );
INVX1 INVX1_450 ( .A(_3147_), .Y(_3148_) );
OAI21X1 OAI21X1_543 ( .A(_3136_), .B(_3137_), .C(_3148_), .Y(_3149_) );
NAND3X1 NAND3X1_472 ( .A(_3192_), .B(_3108_), .C(_3109_), .Y(_3150_) );
NAND2X1 NAND2X1_588 ( .A(_3150_), .B(_3116_), .Y(_3151_) );
AOI21X1 AOI21X1_313 ( .A(_3122_), .B(_3126_), .C(_3151_), .Y(_3152_) );
OAI21X1 OAI21X1_544 ( .A(_3113_), .B(_3114_), .C(_3152_), .Y(_3153_) );
INVX1 INVX1_451 ( .A(_3137_), .Y(_3154_) );
NAND3X1 NAND3X1_473 ( .A(_3154_), .B(_3147_), .C(_3153_), .Y(_3155_) );
AND2X2 AND2X2_153 ( .A(_3149_), .B(_3155_), .Y(micro_ucr_hash1_c_30__6_) );
AOI21X1 AOI21X1_314 ( .A(_3154_), .B(_3153_), .C(_3147_), .Y(_3156_) );
NOR2X1 NOR2X1_345 ( .A(micro_ucr_hash1_b_29__7_), .B(micro_ucr_hash1_a_29__7_), .Y(_3157_) );
XNOR2X1 XNOR2X1_202 ( .A(_3157_), .B(micro_ucr_hash1_W_30__7_), .Y(_3158_) );
XNOR2X1 XNOR2X1_203 ( .A(_3158_), .B(_3139_), .Y(_3159_) );
OAI21X1 OAI21X1_545 ( .A(_3156_), .B(_3144_), .C(_3159_), .Y(_3160_) );
INVX1 INVX1_452 ( .A(_3159_), .Y(_3161_) );
NAND3X1 NAND3X1_474 ( .A(_3145_), .B(_3161_), .C(_3149_), .Y(_3162_) );
NAND2X1 NAND2X1_589 ( .A(_3160_), .B(_3162_), .Y(micro_ucr_hash1_c_30__7_) );
XOR2X1 XOR2X1_288 ( .A(micro_ucr_hash1_b_31__4_), .B(gnd), .Y(micro_ucr_hash1_a_31__0_) );
XOR2X1 XOR2X1_289 ( .A(micro_ucr_hash1_b_31__5_), .B(gnd), .Y(micro_ucr_hash1_a_31__1_) );
XOR2X1 XOR2X1_290 ( .A(micro_ucr_hash1_b_31__6_), .B(gnd), .Y(micro_ucr_hash1_a_31__2_) );
XOR2X1 XOR2X1_291 ( .A(micro_ucr_hash1_b_31__7_), .B(gnd), .Y(micro_ucr_hash1_a_31__3_) );
XOR2X1 XOR2X1_292 ( .A(micro_ucr_hash1_c_30__4_), .B(micro_ucr_hash1_b_30__4_), .Y(micro_ucr_hash1_a_31__4_) );
XOR2X1 XOR2X1_293 ( .A(micro_ucr_hash1_c_30__5_), .B(micro_ucr_hash1_b_30__5_), .Y(micro_ucr_hash1_a_31__5_) );
XOR2X1 XOR2X1_294 ( .A(micro_ucr_hash1_c_30__6_), .B(micro_ucr_hash1_b_30__6_), .Y(micro_ucr_hash1_a_31__6_) );
XOR2X1 XOR2X1_295 ( .A(micro_ucr_hash1_c_30__7_), .B(micro_ucr_hash1_b_30__7_), .Y(micro_ucr_hash1_a_31__7_) );
INVX1 INVX1_453 ( .A(micro_ucr_hash1_W_31__0_), .Y(_3258_) );
NOR2X1 NOR2X1_346 ( .A(gnd), .B(micro_ucr_hash1_a_30__0_), .Y(_3259_) );
NAND2X1 NAND2X1_590 ( .A(_3258_), .B(_3259_), .Y(_3260_) );
OAI21X1 OAI21X1_546 ( .A(gnd), .B(micro_ucr_hash1_a_30__0_), .C(micro_ucr_hash1_W_31__0_), .Y(_3261_) );
NAND2X1 NAND2X1_591 ( .A(_3261_), .B(_3260_), .Y(micro_ucr_hash1_c_31__0_) );
OAI21X1 OAI21X1_547 ( .A(gnd), .B(micro_ucr_hash1_a_30__1_), .C(micro_ucr_hash1_W_31__1_), .Y(_3262_) );
INVX1 INVX1_454 ( .A(micro_ucr_hash1_W_31__1_), .Y(_3263_) );
NOR2X1 NOR2X1_347 ( .A(gnd), .B(micro_ucr_hash1_a_30__1_), .Y(_3264_) );
NAND2X1 NAND2X1_592 ( .A(_3263_), .B(_3264_), .Y(_3265_) );
NAND3X1 NAND3X1_475 ( .A(_3262_), .B(_3260_), .C(_3265_), .Y(_3266_) );
AND2X2 AND2X2_154 ( .A(_3259_), .B(_3258_), .Y(_3267_) );
INVX2 INVX2_73 ( .A(_3262_), .Y(_3268_) );
AND2X2 AND2X2_155 ( .A(_3264_), .B(_3263_), .Y(_3269_) );
OAI21X1 OAI21X1_548 ( .A(_3269_), .B(_3268_), .C(_3267_), .Y(_3270_) );
AND2X2 AND2X2_156 ( .A(_3270_), .B(_3266_), .Y(micro_ucr_hash1_c_31__1_) );
OAI21X1 OAI21X1_549 ( .A(gnd), .B(micro_ucr_hash1_a_30__2_), .C(micro_ucr_hash1_W_31__2_), .Y(_3271_) );
INVX1 INVX1_455 ( .A(micro_ucr_hash1_W_31__2_), .Y(_3272_) );
NOR2X1 NOR2X1_348 ( .A(gnd), .B(micro_ucr_hash1_a_30__2_), .Y(_3273_) );
NAND2X1 NAND2X1_593 ( .A(_3272_), .B(_3273_), .Y(_3274_) );
NAND2X1 NAND2X1_594 ( .A(_3271_), .B(_3274_), .Y(_3275_) );
NAND3X1 NAND3X1_476 ( .A(_3271_), .B(_3274_), .C(_3268_), .Y(_3276_) );
OAI21X1 OAI21X1_550 ( .A(_3266_), .B(_3275_), .C(_3276_), .Y(_3277_) );
INVX1 INVX1_456 ( .A(_3275_), .Y(_3278_) );
OAI21X1 OAI21X1_551 ( .A(_3267_), .B(_3269_), .C(_3262_), .Y(_3279_) );
NOR2X1 NOR2X1_349 ( .A(_3279_), .B(_3278_), .Y(_3280_) );
NOR2X1 NOR2X1_350 ( .A(_3277_), .B(_3280_), .Y(micro_ucr_hash1_c_31__2_) );
INVX1 INVX1_457 ( .A(micro_ucr_hash1_W_31__3_), .Y(_3281_) );
OAI21X1 OAI21X1_552 ( .A(gnd), .B(micro_ucr_hash1_a_30__3_), .C(_3281_), .Y(_3282_) );
NOR2X1 NOR2X1_351 ( .A(gnd), .B(micro_ucr_hash1_a_30__3_), .Y(_3283_) );
NAND2X1 NAND2X1_595 ( .A(micro_ucr_hash1_W_31__3_), .B(_3283_), .Y(_3284_) );
NAND3X1 NAND3X1_477 ( .A(_3271_), .B(_3282_), .C(_3284_), .Y(_3285_) );
INVX1 INVX1_458 ( .A(_3271_), .Y(_3286_) );
OAI21X1 OAI21X1_553 ( .A(gnd), .B(micro_ucr_hash1_a_30__3_), .C(micro_ucr_hash1_W_31__3_), .Y(_3287_) );
NAND2X1 NAND2X1_596 ( .A(_3281_), .B(_3283_), .Y(_3288_) );
NAND3X1 NAND3X1_478 ( .A(_3287_), .B(_3288_), .C(_3286_), .Y(_3289_) );
NAND2X1 NAND2X1_597 ( .A(_3285_), .B(_3289_), .Y(_3290_) );
XNOR2X1 XNOR2X1_204 ( .A(_3277_), .B(_3290_), .Y(micro_ucr_hash1_c_31__3_) );
INVX1 INVX1_459 ( .A(_3287_), .Y(_3291_) );
OAI21X1 OAI21X1_554 ( .A(micro_ucr_hash1_b_30__4_), .B(micro_ucr_hash1_a_30__4_), .C(micro_ucr_hash1_W_31__4_), .Y(_3292_) );
INVX1 INVX1_460 ( .A(micro_ucr_hash1_b_30__4_), .Y(_3293_) );
INVX1 INVX1_461 ( .A(micro_ucr_hash1_a_30__4_), .Y(_3294_) );
INVX1 INVX1_462 ( .A(micro_ucr_hash1_W_31__4_), .Y(_3295_) );
NAND3X1 NAND3X1_479 ( .A(_3293_), .B(_3294_), .C(_3295_), .Y(_3296_) );
AOI21X1 AOI21X1_315 ( .A(_3292_), .B(_3296_), .C(_3291_), .Y(_3202_) );
OAI21X1 OAI21X1_555 ( .A(micro_ucr_hash1_b_30__4_), .B(micro_ucr_hash1_a_30__4_), .C(_3295_), .Y(_3203_) );
NAND3X1 NAND3X1_480 ( .A(micro_ucr_hash1_W_31__4_), .B(_3293_), .C(_3294_), .Y(_3204_) );
AOI21X1 AOI21X1_316 ( .A(_3203_), .B(_3204_), .C(_3287_), .Y(_3205_) );
NOR2X1 NOR2X1_352 ( .A(_3205_), .B(_3202_), .Y(_3206_) );
AOI21X1 AOI21X1_317 ( .A(_3287_), .B(_3288_), .C(_3286_), .Y(_3207_) );
OAI21X1 OAI21X1_556 ( .A(_3207_), .B(_3276_), .C(_3289_), .Y(_3208_) );
NOR3X1 NOR3X1_85 ( .A(_3266_), .B(_3275_), .C(_3207_), .Y(_3209_) );
NOR2X1 NOR2X1_353 ( .A(_3208_), .B(_3209_), .Y(_3210_) );
XNOR2X1 XNOR2X1_205 ( .A(_3210_), .B(_3206_), .Y(micro_ucr_hash1_c_31__4_) );
NAND3X1 NAND3X1_481 ( .A(_3292_), .B(_3296_), .C(_3291_), .Y(_3211_) );
OAI21X1 OAI21X1_557 ( .A(_3210_), .B(_3202_), .C(_3211_), .Y(_3212_) );
INVX1 INVX1_463 ( .A(micro_ucr_hash1_W_31__5_), .Y(_3213_) );
OAI21X1 OAI21X1_558 ( .A(micro_ucr_hash1_b_30__5_), .B(micro_ucr_hash1_a_30__5_), .C(_3213_), .Y(_3214_) );
NOR2X1 NOR2X1_354 ( .A(micro_ucr_hash1_b_30__5_), .B(micro_ucr_hash1_a_30__5_), .Y(_3215_) );
NAND2X1 NAND2X1_598 ( .A(micro_ucr_hash1_W_31__5_), .B(_3215_), .Y(_3216_) );
NAND3X1 NAND3X1_482 ( .A(_3292_), .B(_3214_), .C(_3216_), .Y(_3217_) );
INVX1 INVX1_464 ( .A(_3292_), .Y(_3218_) );
NAND2X1 NAND2X1_599 ( .A(_3213_), .B(_3215_), .Y(_3219_) );
OAI21X1 OAI21X1_559 ( .A(micro_ucr_hash1_b_30__5_), .B(micro_ucr_hash1_a_30__5_), .C(micro_ucr_hash1_W_31__5_), .Y(_3220_) );
NAND3X1 NAND3X1_483 ( .A(_3220_), .B(_3219_), .C(_3218_), .Y(_3221_) );
NAND2X1 NAND2X1_600 ( .A(_3217_), .B(_3221_), .Y(_3222_) );
XOR2X1 XOR2X1_296 ( .A(_3212_), .B(_3222_), .Y(micro_ucr_hash1_c_31__5_) );
OAI21X1 OAI21X1_560 ( .A(gnd), .B(micro_ucr_hash1_a_30__2_), .C(_3272_), .Y(_3223_) );
NAND2X1 NAND2X1_601 ( .A(micro_ucr_hash1_W_31__2_), .B(_3273_), .Y(_3224_) );
AOI21X1 AOI21X1_318 ( .A(_3223_), .B(_3224_), .C(_3262_), .Y(_3225_) );
INVX1 INVX1_465 ( .A(_3289_), .Y(_3226_) );
AOI21X1 AOI21X1_319 ( .A(_3285_), .B(_3225_), .C(_3226_), .Y(_3227_) );
NOR3X1 NOR3X1_86 ( .A(_3267_), .B(_3268_), .C(_3269_), .Y(_3228_) );
NAND3X1 NAND3X1_484 ( .A(_3278_), .B(_3285_), .C(_3228_), .Y(_3229_) );
NAND2X1 NAND2X1_602 ( .A(_3222_), .B(_3206_), .Y(_3230_) );
AOI21X1 AOI21X1_320 ( .A(_3227_), .B(_3229_), .C(_3230_), .Y(_3231_) );
AOI22X1 AOI22X1_22 ( .A(_3219_), .B(_3220_), .C(_3211_), .D(_3292_), .Y(_3232_) );
INVX1 INVX1_466 ( .A(_3219_), .Y(_3233_) );
OAI21X1 OAI21X1_561 ( .A(micro_ucr_hash1_b_30__6_), .B(micro_ucr_hash1_a_30__6_), .C(micro_ucr_hash1_W_31__6_), .Y(_3234_) );
INVX1 INVX1_467 ( .A(micro_ucr_hash1_W_31__6_), .Y(_3235_) );
NOR2X1 NOR2X1_355 ( .A(micro_ucr_hash1_b_30__6_), .B(micro_ucr_hash1_a_30__6_), .Y(_3236_) );
NAND2X1 NAND2X1_603 ( .A(_3235_), .B(_3236_), .Y(_3237_) );
NAND2X1 NAND2X1_604 ( .A(_3234_), .B(_3237_), .Y(_3238_) );
NOR2X1 NOR2X1_356 ( .A(_3233_), .B(_3238_), .Y(_3239_) );
INVX1 INVX1_468 ( .A(_3239_), .Y(_3240_) );
NAND2X1 NAND2X1_605 ( .A(_3233_), .B(_3238_), .Y(_3241_) );
NAND2X1 NAND2X1_606 ( .A(_3241_), .B(_3240_), .Y(_3242_) );
INVX1 INVX1_469 ( .A(_3242_), .Y(_3243_) );
OAI21X1 OAI21X1_562 ( .A(_3231_), .B(_3232_), .C(_3243_), .Y(_3244_) );
NAND3X1 NAND3X1_485 ( .A(_3287_), .B(_3203_), .C(_3204_), .Y(_3245_) );
NAND2X1 NAND2X1_607 ( .A(_3245_), .B(_3211_), .Y(_3246_) );
AOI21X1 AOI21X1_321 ( .A(_3217_), .B(_3221_), .C(_3246_), .Y(_3247_) );
OAI21X1 OAI21X1_563 ( .A(_3208_), .B(_3209_), .C(_3247_), .Y(_3248_) );
INVX1 INVX1_470 ( .A(_3232_), .Y(_3249_) );
NAND3X1 NAND3X1_486 ( .A(_3249_), .B(_3242_), .C(_3248_), .Y(_3250_) );
AND2X2 AND2X2_157 ( .A(_3244_), .B(_3250_), .Y(micro_ucr_hash1_c_31__6_) );
AOI21X1 AOI21X1_322 ( .A(_3249_), .B(_3248_), .C(_3242_), .Y(_3251_) );
NOR2X1 NOR2X1_357 ( .A(micro_ucr_hash1_b_30__7_), .B(micro_ucr_hash1_a_30__7_), .Y(_3252_) );
XNOR2X1 XNOR2X1_206 ( .A(_3252_), .B(micro_ucr_hash1_W_31__7_), .Y(_3253_) );
XNOR2X1 XNOR2X1_207 ( .A(_3253_), .B(_3234_), .Y(_3254_) );
OAI21X1 OAI21X1_564 ( .A(_3251_), .B(_3239_), .C(_3254_), .Y(_3255_) );
INVX1 INVX1_471 ( .A(_3254_), .Y(_3256_) );
NAND3X1 NAND3X1_487 ( .A(_3240_), .B(_3256_), .C(_3244_), .Y(_3257_) );
NAND2X1 NAND2X1_608 ( .A(_3255_), .B(_3257_), .Y(micro_ucr_hash1_c_31__7_) );
INVX8 INVX8_2 ( .A(reset_bF_buf4), .Y(_3299_) );
INVX1 INVX1_472 ( .A(entrada_hash1_contadores_0_), .Y(_3300_) );
NOR2X1 NOR2X1_358 ( .A(_3299__bF_buf4), .B(_3300_), .Y(_3298__0_) );
AND2X2 AND2X2_158 ( .A(reset_bF_buf2), .B(entrada_hash1_contadores_1_), .Y(_3298__1_) );
AND2X2 AND2X2_159 ( .A(reset_bF_buf0), .B(entrada_hash1_contadores_2_), .Y(_3298__2_) );
INVX2 INVX2_74 ( .A(entrada_hash1_contadores_3_), .Y(_3301_) );
NOR2X1 NOR2X1_359 ( .A(_3299__bF_buf4), .B(_3301_), .Y(_3298__3_) );
INVX1 INVX1_473 ( .A(entrada_hash1_contadores_4_), .Y(_3302_) );
NOR2X1 NOR2X1_360 ( .A(_3299__bF_buf4), .B(_3302_), .Y(_3298__4_) );
INVX1 INVX1_474 ( .A(entrada_hash1_contadores_5_), .Y(_3303_) );
NOR2X1 NOR2X1_361 ( .A(_3299__bF_buf3), .B(_3303_), .Y(_3298__5_) );
AND2X2 AND2X2_160 ( .A(reset_bF_buf3), .B(entrada_hash1_contadores_6_), .Y(_3298__6_) );
INVX1 INVX1_475 ( .A(entrada_hash1_contadores_7_), .Y(_3304_) );
NOR2X1 NOR2X1_362 ( .A(_3299__bF_buf2), .B(_3304_), .Y(_3298__7_) );
AND2X2 AND2X2_161 ( .A(reset_bF_buf2), .B(entrada_hash1_contadores_8_), .Y(_3298__8_) );
INVX1 INVX1_476 ( .A(entrada_hash1_contadores_9_), .Y(_3305_) );
NOR2X1 NOR2X1_363 ( .A(_3299__bF_buf0), .B(_3305_), .Y(_3298__9_) );
AND2X2 AND2X2_162 ( .A(reset_bF_buf2), .B(entrada_hash1_contadores_10_), .Y(_3298__10_) );
AND2X2 AND2X2_163 ( .A(reset_bF_buf2), .B(entrada_hash1_contadores_11_), .Y(_3298__11_) );
INVX1 INVX1_477 ( .A(entrada_hash1_contadores_12_), .Y(_3306_) );
NOR2X1 NOR2X1_364 ( .A(_3299__bF_buf0), .B(_3306_), .Y(_3298__12_) );
AND2X2 AND2X2_164 ( .A(reset_bF_buf4), .B(entrada_hash1_contadores_13_), .Y(_3298__13_) );
INVX1 INVX1_478 ( .A(entrada_hash1_contadores_14_), .Y(_3307_) );
NOR2X1 NOR2X1_365 ( .A(_3299__bF_buf0), .B(_3307_), .Y(_3298__14_) );
INVX2 INVX2_75 ( .A(entrada_hash1_contadores_15_), .Y(_3308_) );
NOR2X1 NOR2X1_366 ( .A(_3299__bF_buf0), .B(_3308_), .Y(_3298__15_) );
INVX2 INVX2_76 ( .A(entrada_hash1_contadores_16_), .Y(_3309_) );
NOR2X1 NOR2X1_367 ( .A(_3299__bF_buf1), .B(_3309_), .Y(_3298__16_) );
AND2X2 AND2X2_165 ( .A(reset_bF_buf1), .B(entrada_hash1_contadores_17_), .Y(_3298__17_) );
AND2X2 AND2X2_166 ( .A(reset_bF_buf4), .B(entrada_hash1_contadores_18_), .Y(_3298__18_) );
INVX1 INVX1_479 ( .A(entrada_hash1_contadores_19_), .Y(_3310_) );
NOR2X1 NOR2X1_368 ( .A(_3299__bF_buf1), .B(_3310_), .Y(_3298__19_) );
INVX1 INVX1_480 ( .A(entrada_hash1_contadores_20_), .Y(_3311_) );
NOR2X1 NOR2X1_369 ( .A(_3299__bF_buf1), .B(_3311_), .Y(_3298__20_) );
INVX2 INVX2_77 ( .A(entrada_hash1_contadores_21_), .Y(_3312_) );
NOR2X1 NOR2X1_370 ( .A(_3299__bF_buf1), .B(_3312_), .Y(_3298__21_) );
INVX1 INVX1_481 ( .A(entrada_hash1_contadores_22_), .Y(_3313_) );
NOR2X1 NOR2X1_371 ( .A(_3299__bF_buf4), .B(_3313_), .Y(_3298__22_) );
INVX1 INVX1_482 ( .A(entrada_hash1_contadores_23_), .Y(_3314_) );
NOR2X1 NOR2X1_372 ( .A(_3299__bF_buf1), .B(_3314_), .Y(_3298__23_) );
INVX2 INVX2_78 ( .A(entrada_hash1_contadores_24_), .Y(_3315_) );
NOR2X1 NOR2X1_373 ( .A(_3299__bF_buf3), .B(_3315_), .Y(_3298__24_) );
INVX2 INVX2_79 ( .A(entrada_hash1_contadores_25_), .Y(_3316_) );
NOR2X1 NOR2X1_374 ( .A(_3299__bF_buf3), .B(_3316_), .Y(_3298__25_) );
AND2X2 AND2X2_167 ( .A(reset_bF_buf3), .B(entrada_hash1_contadores_26_), .Y(_3298__26_) );
INVX1 INVX1_483 ( .A(entrada_hash1_contadores_27_), .Y(_3317_) );
NOR2X1 NOR2X1_375 ( .A(_3299__bF_buf2), .B(_3317_), .Y(_3298__27_) );
INVX1 INVX1_484 ( .A(entrada_hash1_contadores_28_), .Y(_3318_) );
NOR2X1 NOR2X1_376 ( .A(_3299__bF_buf2), .B(_3318_), .Y(_3298__28_) );
INVX2 INVX2_80 ( .A(entrada_hash1_contadores_29_), .Y(_3319_) );
NOR2X1 NOR2X1_377 ( .A(_3299__bF_buf2), .B(_3319_), .Y(_3298__29_) );
INVX2 INVX2_81 ( .A(entrada_hash1_contadores_30_), .Y(_3320_) );
NOR2X1 NOR2X1_378 ( .A(_3299__bF_buf2), .B(_3320_), .Y(_3298__30_) );
INVX1 INVX1_485 ( .A(entrada_hash1_contadores_31_), .Y(_3321_) );
NOR2X1 NOR2X1_379 ( .A(_3299__bF_buf2), .B(_3321_), .Y(_3298__31_) );
INVX1 INVX1_486 ( .A(_127__bF_buf0), .Y(_3322_) );
NAND2X1 NAND2X1_609 ( .A(inicio), .B(_3322_), .Y(_3323_) );
NOR2X1 NOR2X1_380 ( .A(_3300_), .B(_3323_), .Y(_3324_) );
INVX1 INVX1_487 ( .A(inicio), .Y(_3325_) );
NOR2X1 NOR2X1_381 ( .A(_127__bF_buf0), .B(_3325_), .Y(_3326_) );
OAI21X1 OAI21X1_565 ( .A(_3326_), .B(entrada_hash1_contadores_0_), .C(reset_bF_buf5), .Y(_3327_) );
NOR2X1 NOR2X1_382 ( .A(_3324_), .B(_3327_), .Y(_3297__0_) );
NAND2X1 NAND2X1_610 ( .A(entrada_hash1_contadores_0_), .B(entrada_hash1_contadores_1_), .Y(_3328_) );
NOR2X1 NOR2X1_383 ( .A(_3328_), .B(_3323_), .Y(_3329_) );
OAI21X1 OAI21X1_566 ( .A(_3324_), .B(entrada_hash1_contadores_1_), .C(reset_bF_buf5), .Y(_3330_) );
NOR2X1 NOR2X1_384 ( .A(_3329_), .B(_3330_), .Y(_3297__1_) );
OAI21X1 OAI21X1_567 ( .A(_3329_), .B(entrada_hash1_contadores_2_), .C(reset_bF_buf5), .Y(_3331_) );
AOI21X1 AOI21X1_323 ( .A(entrada_hash1_contadores_2_), .B(_3329_), .C(_3331_), .Y(_3297__2_) );
NAND2X1 NAND2X1_611 ( .A(entrada_hash1_contadores_2_), .B(_3329_), .Y(_3332_) );
OAI21X1 OAI21X1_568 ( .A(_3332_), .B(_3301_), .C(reset_bF_buf0), .Y(_3333_) );
AOI21X1 AOI21X1_324 ( .A(_3301_), .B(_3332_), .C(_3333_), .Y(_3297__3_) );
AND2X2 AND2X2_168 ( .A(entrada_hash1_contadores_2_), .B(entrada_hash1_contadores_3_), .Y(_3334_) );
NAND3X1 NAND3X1_488 ( .A(entrada_hash1_contadores_4_), .B(_3334_), .C(_3329_), .Y(_3335_) );
INVX4 INVX4_2 ( .A(_3335_), .Y(_3336_) );
OAI21X1 OAI21X1_569 ( .A(_3332_), .B(_3301_), .C(_3302_), .Y(_3337_) );
NAND2X1 NAND2X1_612 ( .A(reset_bF_buf0), .B(_3337_), .Y(_3338_) );
NOR2X1 NOR2X1_385 ( .A(_3336_), .B(_3338_), .Y(_3297__4_) );
OAI21X1 OAI21X1_570 ( .A(_3336_), .B(entrada_hash1_contadores_5_), .C(reset_bF_buf0), .Y(_3339_) );
AOI21X1 AOI21X1_325 ( .A(entrada_hash1_contadores_5_), .B(_3336_), .C(_3339_), .Y(_3297__5_) );
AOI21X1 AOI21X1_326 ( .A(entrada_hash1_contadores_5_), .B(_3336_), .C(entrada_hash1_contadores_6_), .Y(_3340_) );
NAND2X1 NAND2X1_613 ( .A(entrada_hash1_contadores_5_), .B(entrada_hash1_contadores_6_), .Y(_3341_) );
OAI21X1 OAI21X1_571 ( .A(_3335_), .B(_3341_), .C(reset_bF_buf3), .Y(_3342_) );
NOR2X1 NOR2X1_386 ( .A(_3342_), .B(_3340_), .Y(_3297__6_) );
OAI21X1 OAI21X1_572 ( .A(_3335_), .B(_3341_), .C(entrada_hash1_contadores_7_), .Y(_3343_) );
AND2X2 AND2X2_169 ( .A(entrada_hash1_contadores_5_), .B(entrada_hash1_contadores_6_), .Y(_3344_) );
NAND3X1 NAND3X1_489 ( .A(_3304_), .B(_3344_), .C(_3336_), .Y(_3345_) );
AOI21X1 AOI21X1_327 ( .A(_3343_), .B(_3345_), .C(_3299__bF_buf3), .Y(_3297__7_) );
NAND2X1 NAND2X1_614 ( .A(entrada_hash1_contadores_4_), .B(entrada_hash1_contadores_7_), .Y(_3346_) );
NOR2X1 NOR2X1_387 ( .A(_3328_), .B(_3346_), .Y(_3347_) );
NAND2X1 NAND2X1_615 ( .A(entrada_hash1_contadores_2_), .B(entrada_hash1_contadores_3_), .Y(_3348_) );
NOR2X1 NOR2X1_388 ( .A(_3348_), .B(_3341_), .Y(_3349_) );
NAND3X1 NAND3X1_490 ( .A(_3326_), .B(_3347_), .C(_3349_), .Y(_3350_) );
INVX2 INVX2_82 ( .A(_3350_), .Y(_3351_) );
OAI21X1 OAI21X1_573 ( .A(_3351_), .B(entrada_hash1_contadores_8_), .C(reset_bF_buf1), .Y(_3352_) );
AOI21X1 AOI21X1_328 ( .A(entrada_hash1_contadores_8_), .B(_3351_), .C(_3352_), .Y(_3297__8_) );
NAND2X1 NAND2X1_616 ( .A(entrada_hash1_contadores_8_), .B(_3351_), .Y(_3353_) );
NAND2X1 NAND2X1_617 ( .A(entrada_hash1_contadores_8_), .B(entrada_hash1_contadores_9_), .Y(_3354_) );
OAI21X1 OAI21X1_574 ( .A(_3350_), .B(_3354_), .C(reset_bF_buf1), .Y(_3355_) );
AOI21X1 AOI21X1_329 ( .A(_3305_), .B(_3353_), .C(_3355_), .Y(_3297__9_) );
NOR2X1 NOR2X1_389 ( .A(_3354_), .B(_3350_), .Y(_3356_) );
OAI21X1 OAI21X1_575 ( .A(_3356_), .B(entrada_hash1_contadores_10_), .C(reset_bF_buf1), .Y(_3357_) );
AOI21X1 AOI21X1_330 ( .A(entrada_hash1_contadores_10_), .B(_3356_), .C(_3357_), .Y(_3297__10_) );
NAND3X1 NAND3X1_491 ( .A(entrada_hash1_contadores_8_), .B(entrada_hash1_contadores_9_), .C(entrada_hash1_contadores_10_), .Y(_3358_) );
NOR2X1 NOR2X1_390 ( .A(_3358_), .B(_3350_), .Y(_3359_) );
NOR2X1 NOR2X1_391 ( .A(entrada_hash1_contadores_11_), .B(_3359_), .Y(_3360_) );
NAND2X1 NAND2X1_618 ( .A(entrada_hash1_contadores_11_), .B(_3359_), .Y(_3361_) );
NAND2X1 NAND2X1_619 ( .A(reset_bF_buf2), .B(_3361_), .Y(_3362_) );
NOR2X1 NOR2X1_392 ( .A(_3360_), .B(_3362_), .Y(_3297__11_) );
NOR2X1 NOR2X1_393 ( .A(_3306_), .B(_3361_), .Y(_3363_) );
AOI21X1 AOI21X1_331 ( .A(entrada_hash1_contadores_11_), .B(_3359_), .C(entrada_hash1_contadores_12_), .Y(_3364_) );
NOR3X1 NOR3X1_87 ( .A(_3299__bF_buf0), .B(_3364_), .C(_3363_), .Y(_3297__12_) );
INVX1 INVX1_488 ( .A(_3358_), .Y(_3365_) );
NAND3X1 NAND3X1_492 ( .A(entrada_hash1_contadores_11_), .B(entrada_hash1_contadores_12_), .C(_3365_), .Y(_3366_) );
NOR2X1 NOR2X1_394 ( .A(_3366_), .B(_3350_), .Y(_3367_) );
NOR2X1 NOR2X1_395 ( .A(entrada_hash1_contadores_13_), .B(_3367_), .Y(_3368_) );
NAND2X1 NAND2X1_620 ( .A(entrada_hash1_contadores_13_), .B(_3367_), .Y(_3369_) );
NAND2X1 NAND2X1_621 ( .A(reset_bF_buf4), .B(_3369_), .Y(_3370_) );
NOR2X1 NOR2X1_396 ( .A(_3368_), .B(_3370_), .Y(_3297__13_) );
NOR2X1 NOR2X1_397 ( .A(_3307_), .B(_3369_), .Y(_3371_) );
AOI21X1 AOI21X1_332 ( .A(entrada_hash1_contadores_13_), .B(_3367_), .C(entrada_hash1_contadores_14_), .Y(_3372_) );
NOR3X1 NOR3X1_88 ( .A(_3299__bF_buf0), .B(_3372_), .C(_3371_), .Y(_3297__14_) );
NAND3X1 NAND3X1_493 ( .A(entrada_hash1_contadores_10_), .B(entrada_hash1_contadores_11_), .C(entrada_hash1_contadores_12_), .Y(_3373_) );
INVX1 INVX1_489 ( .A(_3373_), .Y(_3374_) );
NAND2X1 NAND2X1_622 ( .A(entrada_hash1_contadores_13_), .B(entrada_hash1_contadores_14_), .Y(_3375_) );
NOR2X1 NOR2X1_398 ( .A(_3354_), .B(_3375_), .Y(_3376_) );
NAND2X1 NAND2X1_623 ( .A(_3374_), .B(_3376_), .Y(_3377_) );
NOR2X1 NOR2X1_399 ( .A(_3377_), .B(_3350_), .Y(_3378_) );
OAI21X1 OAI21X1_576 ( .A(_3378_), .B(entrada_hash1_contadores_15_), .C(reset_bF_buf1), .Y(_3379_) );
AOI21X1 AOI21X1_333 ( .A(entrada_hash1_contadores_15_), .B(_3378_), .C(_3379_), .Y(_3297__15_) );
INVX2 INVX2_83 ( .A(_3378_), .Y(_3380_) );
OAI21X1 OAI21X1_577 ( .A(_3380_), .B(_3308_), .C(_3309_), .Y(_3381_) );
NOR2X1 NOR2X1_400 ( .A(_3308_), .B(_3309_), .Y(_3382_) );
AOI21X1 AOI21X1_334 ( .A(_3382_), .B(_3378_), .C(_3299__bF_buf1), .Y(_3383_) );
AND2X2 AND2X2_170 ( .A(_3381_), .B(_3383_), .Y(_3297__16_) );
AOI21X1 AOI21X1_335 ( .A(_3382_), .B(_3378_), .C(entrada_hash1_contadores_17_), .Y(_3384_) );
NAND3X1 NAND3X1_494 ( .A(entrada_hash1_contadores_15_), .B(entrada_hash1_contadores_16_), .C(entrada_hash1_contadores_17_), .Y(_3385_) );
OAI21X1 OAI21X1_578 ( .A(_3380_), .B(_3385_), .C(reset_bF_buf5), .Y(_3386_) );
NOR2X1 NOR2X1_401 ( .A(_3384_), .B(_3386_), .Y(_3297__17_) );
INVX1 INVX1_490 ( .A(_3385_), .Y(_3387_) );
AND2X2 AND2X2_171 ( .A(_3378_), .B(_3387_), .Y(_3388_) );
OAI21X1 OAI21X1_579 ( .A(_3388_), .B(entrada_hash1_contadores_18_), .C(reset_bF_buf4), .Y(_3389_) );
AOI21X1 AOI21X1_336 ( .A(entrada_hash1_contadores_18_), .B(_3388_), .C(_3389_), .Y(_3297__18_) );
NAND2X1 NAND2X1_624 ( .A(entrada_hash1_contadores_18_), .B(_3388_), .Y(_3390_) );
NAND2X1 NAND2X1_625 ( .A(entrada_hash1_contadores_18_), .B(entrada_hash1_contadores_19_), .Y(_3391_) );
NOR2X1 NOR2X1_402 ( .A(_3391_), .B(_3385_), .Y(_3392_) );
NAND2X1 NAND2X1_626 ( .A(_3392_), .B(_3378_), .Y(_3393_) );
NAND2X1 NAND2X1_627 ( .A(reset_bF_buf4), .B(_3393_), .Y(_3394_) );
AOI21X1 AOI21X1_337 ( .A(_3310_), .B(_3390_), .C(_3394_), .Y(_3297__19_) );
AND2X2 AND2X2_172 ( .A(_3378_), .B(_3392_), .Y(_3395_) );
OAI21X1 OAI21X1_580 ( .A(_3395_), .B(entrada_hash1_contadores_20_), .C(reset_bF_buf5), .Y(_3396_) );
AOI21X1 AOI21X1_338 ( .A(entrada_hash1_contadores_20_), .B(_3395_), .C(_3396_), .Y(_3297__20_) );
NAND2X1 NAND2X1_628 ( .A(entrada_hash1_contadores_20_), .B(_3395_), .Y(_3397_) );
NOR2X1 NOR2X1_403 ( .A(_3311_), .B(_3312_), .Y(_3398_) );
NAND2X1 NAND2X1_629 ( .A(_3398_), .B(_3392_), .Y(_3399_) );
OAI21X1 OAI21X1_581 ( .A(_3380_), .B(_3399_), .C(reset_bF_buf2), .Y(_3400_) );
AOI21X1 AOI21X1_339 ( .A(_3312_), .B(_3397_), .C(_3400_), .Y(_3297__21_) );
INVX2 INVX2_84 ( .A(_3399_), .Y(_3401_) );
AND2X2 AND2X2_173 ( .A(_3378_), .B(_3401_), .Y(_3402_) );
OAI21X1 OAI21X1_582 ( .A(_3402_), .B(entrada_hash1_contadores_22_), .C(reset_bF_buf5), .Y(_3403_) );
AOI21X1 AOI21X1_340 ( .A(entrada_hash1_contadores_22_), .B(_3402_), .C(_3403_), .Y(_3297__22_) );
NAND2X1 NAND2X1_630 ( .A(_3401_), .B(_3378_), .Y(_3404_) );
OAI21X1 OAI21X1_583 ( .A(_3404_), .B(_3313_), .C(entrada_hash1_contadores_23_), .Y(_3405_) );
NAND3X1 NAND3X1_495 ( .A(entrada_hash1_contadores_22_), .B(_3314_), .C(_3402_), .Y(_3406_) );
AOI21X1 AOI21X1_341 ( .A(_3405_), .B(_3406_), .C(_3299__bF_buf4), .Y(_3297__23_) );
NAND2X1 NAND2X1_631 ( .A(entrada_hash1_contadores_22_), .B(entrada_hash1_contadores_23_), .Y(_3407_) );
NOR3X1 NOR3X1_89 ( .A(_3325_), .B(_127__bF_buf0), .C(_3407_), .Y(_3408_) );
NAND3X1 NAND3X1_496 ( .A(_3347_), .B(_3349_), .C(_3408_), .Y(_3409_) );
NOR3X1 NOR3X1_90 ( .A(_3399_), .B(_3377_), .C(_3409_), .Y(_3410_) );
OAI21X1 OAI21X1_584 ( .A(_3410_), .B(entrada_hash1_contadores_24_), .C(reset_bF_buf3), .Y(_3411_) );
AOI21X1 AOI21X1_342 ( .A(entrada_hash1_contadores_24_), .B(_3410_), .C(_3411_), .Y(_3297__24_) );
INVX1 INVX1_491 ( .A(_3377_), .Y(_3412_) );
OR2X2 OR2X2_129 ( .A(_3328_), .B(_3346_), .Y(_3413_) );
NAND2X1 NAND2X1_632 ( .A(_3334_), .B(_3344_), .Y(_3414_) );
AND2X2 AND2X2_174 ( .A(entrada_hash1_contadores_22_), .B(entrada_hash1_contadores_23_), .Y(_3415_) );
NAND3X1 NAND3X1_497 ( .A(inicio), .B(_3322_), .C(_3415_), .Y(_3416_) );
NOR3X1 NOR3X1_91 ( .A(_3413_), .B(_3414_), .C(_3416_), .Y(_3417_) );
NAND3X1 NAND3X1_498 ( .A(_3412_), .B(_3417_), .C(_3401_), .Y(_3418_) );
OAI21X1 OAI21X1_585 ( .A(_3418_), .B(_3315_), .C(_3316_), .Y(_3419_) );
NOR2X1 NOR2X1_404 ( .A(_3315_), .B(_3316_), .Y(_3420_) );
AOI21X1 AOI21X1_343 ( .A(_3420_), .B(_3410_), .C(_3299__bF_buf3), .Y(_3421_) );
AND2X2 AND2X2_175 ( .A(_3419_), .B(_3421_), .Y(_3297__25_) );
AOI21X1 AOI21X1_344 ( .A(_3420_), .B(_3410_), .C(entrada_hash1_contadores_26_), .Y(_3422_) );
NAND3X1 NAND3X1_499 ( .A(entrada_hash1_contadores_24_), .B(entrada_hash1_contadores_25_), .C(entrada_hash1_contadores_26_), .Y(_3423_) );
OAI21X1 OAI21X1_586 ( .A(_3418_), .B(_3423_), .C(reset_bF_buf3), .Y(_3424_) );
NOR2X1 NOR2X1_405 ( .A(_3422_), .B(_3424_), .Y(_3297__26_) );
NOR3X1 NOR3X1_92 ( .A(_3317_), .B(_3423_), .C(_3418_), .Y(_3425_) );
INVX1 INVX1_492 ( .A(_3423_), .Y(_3426_) );
AOI21X1 AOI21X1_345 ( .A(_3426_), .B(_3410_), .C(entrada_hash1_contadores_27_), .Y(_3427_) );
NOR3X1 NOR3X1_93 ( .A(_3299__bF_buf3), .B(_3427_), .C(_3425_), .Y(_3297__27_) );
NAND3X1 NAND3X1_500 ( .A(entrada_hash1_contadores_27_), .B(_3426_), .C(_3410_), .Y(_3428_) );
NAND2X1 NAND2X1_633 ( .A(_3347_), .B(_3349_), .Y(_3429_) );
NOR3X1 NOR3X1_94 ( .A(_3377_), .B(_3416_), .C(_3429_), .Y(_3430_) );
NAND2X1 NAND2X1_634 ( .A(entrada_hash1_contadores_27_), .B(entrada_hash1_contadores_28_), .Y(_3431_) );
NOR2X1 NOR2X1_406 ( .A(_3431_), .B(_3423_), .Y(_3432_) );
NAND3X1 NAND3X1_501 ( .A(_3401_), .B(_3432_), .C(_3430_), .Y(_3433_) );
NAND2X1 NAND2X1_635 ( .A(reset_bF_buf0), .B(_3433_), .Y(_3434_) );
AOI21X1 AOI21X1_346 ( .A(_3318_), .B(_3428_), .C(_3434_), .Y(_3297__28_) );
OAI21X1 OAI21X1_587 ( .A(_3433_), .B(_3319_), .C(reset_bF_buf0), .Y(_3435_) );
AOI21X1 AOI21X1_347 ( .A(_3319_), .B(_3433_), .C(_3435_), .Y(_3297__29_) );
NAND3X1 NAND3X1_502 ( .A(entrada_hash1_contadores_29_), .B(_3432_), .C(_3410_), .Y(_3436_) );
NAND2X1 NAND2X1_636 ( .A(entrada_hash1_contadores_29_), .B(entrada_hash1_contadores_30_), .Y(_3437_) );
OAI21X1 OAI21X1_588 ( .A(_3433_), .B(_3437_), .C(reset_bF_buf3), .Y(_3438_) );
AOI21X1 AOI21X1_348 ( .A(_3320_), .B(_3436_), .C(_3438_), .Y(_3297__30_) );
NAND2X1 NAND2X1_637 ( .A(entrada_hash1_contadores_29_), .B(_3432_), .Y(_3439_) );
NOR2X1 NOR2X1_407 ( .A(_3320_), .B(_3439_), .Y(_3440_) );
AOI21X1 AOI21X1_349 ( .A(_3440_), .B(_3410_), .C(entrada_hash1_contadores_31_), .Y(_3441_) );
OR2X2 OR2X2_130 ( .A(_3439_), .B(_3320_), .Y(_3442_) );
NOR3X1 NOR3X1_95 ( .A(_3321_), .B(_3442_), .C(_3418_), .Y(_3443_) );
NOR3X1 NOR3X1_96 ( .A(_3299__bF_buf4), .B(_3441_), .C(_3443_), .Y(_3297__31_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf3), .D(_3298__0_), .Q(entrada_hash1_nonce_0_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf7), .D(_3298__1_), .Q(entrada_hash1_nonce_1_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf9), .D(_3298__2_), .Q(entrada_hash1_nonce_2_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf3), .D(_3298__3_), .Q(entrada_hash1_nonce_3_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf5), .D(_3298__4_), .Q(entrada_hash1_nonce_4_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf9), .D(_3298__5_), .Q(entrada_hash1_nonce_5_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf9), .D(_3298__6_), .Q(entrada_hash1_nonce_6_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf5), .D(_3298__7_), .Q(entrada_hash1_nonce_7_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf7), .D(_3298__8_), .Q(entrada_hash1_nonce_8_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf7), .D(_3298__9_), .Q(entrada_hash1_nonce_9_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf7), .D(_3298__10_), .Q(entrada_hash1_nonce_10_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf7), .D(_3298__11_), .Q(entrada_hash1_nonce_11_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf7), .D(_3298__12_), .Q(entrada_hash1_nonce_12_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf7), .D(_3298__13_), .Q(entrada_hash1_nonce_13_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf5), .D(_3298__14_), .Q(entrada_hash1_nonce_14_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf7), .D(_3298__15_), .Q(entrada_hash1_nonce_15_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf1), .D(_3298__16_), .Q(entrada_hash1_nonce_16_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf1), .D(_3298__17_), .Q(entrada_hash1_nonce_17_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf3), .D(_3298__18_), .Q(entrada_hash1_nonce_18_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf7), .D(_3298__19_), .Q(entrada_hash1_nonce_19_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf3), .D(_3298__20_), .Q(entrada_hash1_nonce_20_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf7), .D(_3298__21_), .Q(entrada_hash1_nonce_21_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf5), .D(_3298__22_), .Q(entrada_hash1_nonce_22_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf7), .D(_3298__23_), .Q(entrada_hash1_nonce_23_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf5), .D(_3298__24_), .Q(entrada_hash1_nonce_24_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf5), .D(_3298__25_), .Q(entrada_hash1_nonce_25_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf9), .D(_3298__26_), .Q(entrada_hash1_nonce_26_) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf5), .D(_3298__27_), .Q(entrada_hash1_nonce_27_) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf5), .D(_3298__28_), .Q(entrada_hash1_nonce_28_) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf5), .D(_3298__29_), .Q(entrada_hash1_nonce_29_) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf5), .D(_3298__30_), .Q(entrada_hash1_nonce_30_) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf5), .D(_3298__31_), .Q(entrada_hash1_nonce_31_) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf4), .D(_3297__0_), .Q(entrada_hash1_contadores_0_) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf4), .D(_3297__1_), .Q(entrada_hash1_contadores_1_) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf4), .D(_3297__2_), .Q(entrada_hash1_contadores_2_) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf4), .D(_3297__3_), .Q(entrada_hash1_contadores_3_) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf4), .D(_3297__4_), .Q(entrada_hash1_contadores_4_) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf9), .D(_3297__5_), .Q(entrada_hash1_contadores_5_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf9), .D(_3297__6_), .Q(entrada_hash1_contadores_6_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf4), .D(_3297__7_), .Q(entrada_hash1_contadores_7_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf1), .D(_3297__8_), .Q(entrada_hash1_contadores_8_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf1), .D(_3297__9_), .Q(entrada_hash1_contadores_9_) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf1), .D(_3297__10_), .Q(entrada_hash1_contadores_10_) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf1), .D(_3297__11_), .Q(entrada_hash1_contadores_11_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf7), .D(_3297__12_), .Q(entrada_hash1_contadores_12_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf3), .D(_3297__13_), .Q(entrada_hash1_contadores_13_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf3), .D(_3297__14_), .Q(entrada_hash1_contadores_14_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf1), .D(_3297__15_), .Q(entrada_hash1_contadores_15_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf1), .D(_3297__16_), .Q(entrada_hash1_contadores_16_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf1), .D(_3297__17_), .Q(entrada_hash1_contadores_17_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf3), .D(_3297__18_), .Q(entrada_hash1_contadores_18_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf3), .D(_3297__19_), .Q(entrada_hash1_contadores_19_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf4), .D(_3297__20_), .Q(entrada_hash1_contadores_20_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf1), .D(_3297__21_), .Q(entrada_hash1_contadores_21_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf4), .D(_3297__22_), .Q(entrada_hash1_contadores_22_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf3), .D(_3297__23_), .Q(entrada_hash1_contadores_23_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf9), .D(_3297__24_), .Q(entrada_hash1_contadores_24_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf9), .D(_3297__25_), .Q(entrada_hash1_contadores_25_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf9), .D(_3297__26_), .Q(entrada_hash1_contadores_26_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf9), .D(_3297__27_), .Q(entrada_hash1_contadores_27_) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf9), .D(_3297__28_), .Q(entrada_hash1_contadores_28_) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf3), .D(_3297__29_), .Q(entrada_hash1_contadores_29_) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf9), .D(_3297__30_), .Q(entrada_hash1_contadores_30_) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf3), .D(_3297__31_), .Q(entrada_hash1_contadores_31_) );
INVX1 INVX1_493 ( .A(bloque_bytes[24]), .Y(_3445_) );
AOI21X1 AOI21X1_350 ( .A(bloque_bytes[64]), .B(_3445_), .C(entrada_hash1_nonce_8_), .Y(_3446_) );
OAI21X1 OAI21X1_589 ( .A(bloque_bytes[64]), .B(_3445_), .C(_3446_), .Y(micro_ucr_hash1_W_17__0_) );
INVX1 INVX1_494 ( .A(bloque_bytes[25]), .Y(_3447_) );
AOI21X1 AOI21X1_351 ( .A(bloque_bytes[65]), .B(_3447_), .C(entrada_hash1_nonce_9_), .Y(_3448_) );
OAI21X1 OAI21X1_590 ( .A(bloque_bytes[65]), .B(_3447_), .C(_3448_), .Y(micro_ucr_hash1_W_17__1_) );
INVX1 INVX1_495 ( .A(bloque_bytes[26]), .Y(_3449_) );
AOI21X1 AOI21X1_352 ( .A(bloque_bytes[66]), .B(_3449_), .C(entrada_hash1_nonce_10_), .Y(_3450_) );
OAI21X1 OAI21X1_591 ( .A(bloque_bytes[66]), .B(_3449_), .C(_3450_), .Y(micro_ucr_hash1_W_17__2_) );
INVX1 INVX1_496 ( .A(bloque_bytes[27]), .Y(_3451_) );
AOI21X1 AOI21X1_353 ( .A(bloque_bytes[67]), .B(_3451_), .C(entrada_hash1_nonce_11_), .Y(_3452_) );
OAI21X1 OAI21X1_592 ( .A(bloque_bytes[67]), .B(_3451_), .C(_3452_), .Y(micro_ucr_hash1_W_17__3_) );
INVX1 INVX1_497 ( .A(bloque_bytes[28]), .Y(_3453_) );
AOI21X1 AOI21X1_354 ( .A(bloque_bytes[68]), .B(_3453_), .C(entrada_hash1_nonce_12_), .Y(_3454_) );
OAI21X1 OAI21X1_593 ( .A(bloque_bytes[68]), .B(_3453_), .C(_3454_), .Y(micro_ucr_hash1_W_17__4_) );
INVX1 INVX1_498 ( .A(bloque_bytes[29]), .Y(_3455_) );
AOI21X1 AOI21X1_355 ( .A(bloque_bytes[69]), .B(_3455_), .C(entrada_hash1_nonce_13_), .Y(_3456_) );
OAI21X1 OAI21X1_594 ( .A(bloque_bytes[69]), .B(_3455_), .C(_3456_), .Y(micro_ucr_hash1_W_17__5_) );
INVX1 INVX1_499 ( .A(bloque_bytes[30]), .Y(_3457_) );
AOI21X1 AOI21X1_356 ( .A(bloque_bytes[70]), .B(_3457_), .C(entrada_hash1_nonce_14_), .Y(_3458_) );
OAI21X1 OAI21X1_595 ( .A(bloque_bytes[70]), .B(_3457_), .C(_3458_), .Y(micro_ucr_hash1_W_17__6_) );
INVX1 INVX1_500 ( .A(bloque_bytes[31]), .Y(_3459_) );
AOI21X1 AOI21X1_357 ( .A(bloque_bytes[71]), .B(_3459_), .C(entrada_hash1_nonce_15_), .Y(_3460_) );
OAI21X1 OAI21X1_596 ( .A(bloque_bytes[71]), .B(_3459_), .C(_3460_), .Y(micro_ucr_hash1_W_17__7_) );
INVX1 INVX1_501 ( .A(entrada_hash1_nonce_16_), .Y(_3461_) );
OR2X2 OR2X2_131 ( .A(bloque_bytes[72]), .B(bloque_bytes[32]), .Y(_3462_) );
NAND2X1 NAND2X1_638 ( .A(bloque_bytes[72]), .B(bloque_bytes[32]), .Y(_3463_) );
NAND2X1 NAND2X1_639 ( .A(_3463_), .B(_3462_), .Y(_3464_) );
NAND2X1 NAND2X1_640 ( .A(_3461_), .B(_3464_), .Y(micro_ucr_hash1_W_16__0_) );
INVX1 INVX1_502 ( .A(entrada_hash1_nonce_17_), .Y(_3465_) );
OR2X2 OR2X2_132 ( .A(bloque_bytes[73]), .B(bloque_bytes[33]), .Y(_3466_) );
NAND2X1 NAND2X1_641 ( .A(bloque_bytes[73]), .B(bloque_bytes[33]), .Y(_3467_) );
NAND2X1 NAND2X1_642 ( .A(_3467_), .B(_3466_), .Y(_3468_) );
NAND2X1 NAND2X1_643 ( .A(_3465_), .B(_3468_), .Y(micro_ucr_hash1_W_16__1_) );
INVX2 INVX2_85 ( .A(bloque_bytes[34]), .Y(_3469_) );
AOI21X1 AOI21X1_358 ( .A(bloque_bytes[74]), .B(_3469_), .C(entrada_hash1_nonce_18_), .Y(_3470_) );
OAI21X1 OAI21X1_597 ( .A(bloque_bytes[74]), .B(_3469_), .C(_3470_), .Y(micro_ucr_hash1_W_16__2_) );
INVX1 INVX1_503 ( .A(entrada_hash1_nonce_19_), .Y(_3471_) );
OR2X2 OR2X2_133 ( .A(bloque_bytes[75]), .B(bloque_bytes[35]), .Y(_3472_) );
NAND2X1 NAND2X1_644 ( .A(bloque_bytes[75]), .B(bloque_bytes[35]), .Y(_3473_) );
NAND2X1 NAND2X1_645 ( .A(_3473_), .B(_3472_), .Y(_3474_) );
NAND2X1 NAND2X1_646 ( .A(_3471_), .B(_3474_), .Y(micro_ucr_hash1_W_16__3_) );
INVX1 INVX1_504 ( .A(entrada_hash1_nonce_20_), .Y(_3475_) );
OR2X2 OR2X2_134 ( .A(bloque_bytes[76]), .B(bloque_bytes[36]), .Y(_3476_) );
NAND2X1 NAND2X1_647 ( .A(bloque_bytes[76]), .B(bloque_bytes[36]), .Y(_3477_) );
NAND2X1 NAND2X1_648 ( .A(_3477_), .B(_3476_), .Y(_3478_) );
NAND2X1 NAND2X1_649 ( .A(_3475_), .B(_3478_), .Y(micro_ucr_hash1_W_16__4_) );
INVX2 INVX2_86 ( .A(bloque_bytes[37]), .Y(_3479_) );
AOI21X1 AOI21X1_359 ( .A(bloque_bytes[77]), .B(_3479_), .C(entrada_hash1_nonce_21_), .Y(_3480_) );
OAI21X1 OAI21X1_598 ( .A(bloque_bytes[77]), .B(_3479_), .C(_3480_), .Y(micro_ucr_hash1_W_16__5_) );
INVX2 INVX2_87 ( .A(bloque_bytes[38]), .Y(_3481_) );
AOI21X1 AOI21X1_360 ( .A(bloque_bytes[78]), .B(_3481_), .C(entrada_hash1_nonce_22_), .Y(_3482_) );
OAI21X1 OAI21X1_599 ( .A(bloque_bytes[78]), .B(_3481_), .C(_3482_), .Y(micro_ucr_hash1_W_16__6_) );
INVX1 INVX1_505 ( .A(bloque_bytes[39]), .Y(_3483_) );
AOI21X1 AOI21X1_361 ( .A(bloque_bytes[79]), .B(_3483_), .C(entrada_hash1_nonce_23_), .Y(_3484_) );
OAI21X1 OAI21X1_600 ( .A(bloque_bytes[79]), .B(_3483_), .C(_3484_), .Y(micro_ucr_hash1_W_16__7_) );
INVX1 INVX1_506 ( .A(bloque_bytes[56]), .Y(_3485_) );
INVX1 INVX1_507 ( .A(entrada_hash1_nonce_0_), .Y(_3486_) );
OAI21X1 OAI21X1_601 ( .A(_3485_), .B(bloque_bytes[16]), .C(_3486_), .Y(_3487_) );
AOI21X1 AOI21X1_362 ( .A(_3485_), .B(bloque_bytes[16]), .C(_3487_), .Y(_3488_) );
INVX1 INVX1_508 ( .A(_3488_), .Y(micro_ucr_hash1_W_18__0_) );
INVX1 INVX1_509 ( .A(bloque_bytes[57]), .Y(_3489_) );
INVX1 INVX1_510 ( .A(entrada_hash1_nonce_1_), .Y(_3490_) );
OAI21X1 OAI21X1_602 ( .A(_3489_), .B(bloque_bytes[17]), .C(_3490_), .Y(_3491_) );
AOI21X1 AOI21X1_363 ( .A(_3489_), .B(bloque_bytes[17]), .C(_3491_), .Y(_3492_) );
INVX1 INVX1_511 ( .A(_3492_), .Y(micro_ucr_hash1_W_18__1_) );
INVX1 INVX1_512 ( .A(bloque_bytes[58]), .Y(_3493_) );
INVX1 INVX1_513 ( .A(entrada_hash1_nonce_2_), .Y(_3494_) );
OAI21X1 OAI21X1_603 ( .A(_3493_), .B(bloque_bytes[18]), .C(_3494_), .Y(_3495_) );
AOI21X1 AOI21X1_364 ( .A(_3493_), .B(bloque_bytes[18]), .C(_3495_), .Y(_3496_) );
INVX1 INVX1_514 ( .A(_3496_), .Y(micro_ucr_hash1_W_18__2_) );
INVX1 INVX1_515 ( .A(bloque_bytes[59]), .Y(_3497_) );
INVX1 INVX1_516 ( .A(entrada_hash1_nonce_3_), .Y(_3498_) );
OAI21X1 OAI21X1_604 ( .A(_3497_), .B(bloque_bytes[19]), .C(_3498_), .Y(_3499_) );
AOI21X1 AOI21X1_365 ( .A(_3497_), .B(bloque_bytes[19]), .C(_3499_), .Y(_3500_) );
INVX1 INVX1_517 ( .A(_3500_), .Y(micro_ucr_hash1_W_18__3_) );
INVX1 INVX1_518 ( .A(bloque_bytes[60]), .Y(_3501_) );
INVX1 INVX1_519 ( .A(entrada_hash1_nonce_4_), .Y(_3502_) );
OAI21X1 OAI21X1_605 ( .A(_3501_), .B(bloque_bytes[20]), .C(_3502_), .Y(_3503_) );
AOI21X1 AOI21X1_366 ( .A(_3501_), .B(bloque_bytes[20]), .C(_3503_), .Y(_3504_) );
INVX1 INVX1_520 ( .A(_3504_), .Y(micro_ucr_hash1_W_18__4_) );
INVX1 INVX1_521 ( .A(bloque_bytes[61]), .Y(_3505_) );
INVX1 INVX1_522 ( .A(entrada_hash1_nonce_5_), .Y(_3506_) );
OAI21X1 OAI21X1_606 ( .A(_3505_), .B(bloque_bytes[21]), .C(_3506_), .Y(_3507_) );
AOI21X1 AOI21X1_367 ( .A(_3505_), .B(bloque_bytes[21]), .C(_3507_), .Y(_3508_) );
INVX1 INVX1_523 ( .A(_3508_), .Y(micro_ucr_hash1_W_18__5_) );
INVX1 INVX1_524 ( .A(bloque_bytes[62]), .Y(_3509_) );
INVX1 INVX1_525 ( .A(entrada_hash1_nonce_6_), .Y(_3510_) );
OAI21X1 OAI21X1_607 ( .A(_3509_), .B(bloque_bytes[22]), .C(_3510_), .Y(_3511_) );
AOI21X1 AOI21X1_368 ( .A(_3509_), .B(bloque_bytes[22]), .C(_3511_), .Y(_3512_) );
INVX1 INVX1_526 ( .A(_3512_), .Y(micro_ucr_hash1_W_18__6_) );
INVX1 INVX1_527 ( .A(bloque_bytes[63]), .Y(_3513_) );
INVX1 INVX1_528 ( .A(entrada_hash1_nonce_7_), .Y(_3514_) );
OAI21X1 OAI21X1_608 ( .A(_3513_), .B(bloque_bytes[23]), .C(_3514_), .Y(_3515_) );
AOI21X1 AOI21X1_369 ( .A(_3513_), .B(bloque_bytes[23]), .C(_3515_), .Y(_3516_) );
INVX1 INVX1_529 ( .A(_3516_), .Y(micro_ucr_hash1_W_18__7_) );
AOI21X1 AOI21X1_370 ( .A(_3463_), .B(_3462_), .C(entrada_hash1_nonce_16_), .Y(_3517_) );
XNOR2X1 XNOR2X1_208 ( .A(bloque_bytes[48]), .B(bloque_bytes[8]), .Y(_3518_) );
NAND2X1 NAND2X1_650 ( .A(_3518_), .B(_3517_), .Y(micro_ucr_hash1_W_19__0_) );
AOI21X1 AOI21X1_371 ( .A(_3467_), .B(_3466_), .C(entrada_hash1_nonce_17_), .Y(_3519_) );
XNOR2X1 XNOR2X1_209 ( .A(bloque_bytes[49]), .B(bloque_bytes[9]), .Y(_3520_) );
NAND2X1 NAND2X1_651 ( .A(_3520_), .B(_3519_), .Y(micro_ucr_hash1_W_19__1_) );
INVX1 INVX1_530 ( .A(bloque_bytes[74]), .Y(_3521_) );
INVX1 INVX1_531 ( .A(entrada_hash1_nonce_18_), .Y(_3522_) );
OAI21X1 OAI21X1_609 ( .A(_3521_), .B(bloque_bytes[34]), .C(_3522_), .Y(_3523_) );
AOI21X1 AOI21X1_372 ( .A(_3521_), .B(bloque_bytes[34]), .C(_3523_), .Y(_3524_) );
XNOR2X1 XNOR2X1_210 ( .A(bloque_bytes[50]), .B(bloque_bytes[10]), .Y(_3525_) );
NAND2X1 NAND2X1_652 ( .A(_3525_), .B(_3524_), .Y(micro_ucr_hash1_W_19__2_) );
AOI21X1 AOI21X1_373 ( .A(_3473_), .B(_3472_), .C(entrada_hash1_nonce_19_), .Y(_3526_) );
XNOR2X1 XNOR2X1_211 ( .A(bloque_bytes[51]), .B(bloque_bytes[11]), .Y(_3527_) );
NAND2X1 NAND2X1_653 ( .A(_3527_), .B(_3526_), .Y(micro_ucr_hash1_W_19__3_) );
AOI21X1 AOI21X1_374 ( .A(_3477_), .B(_3476_), .C(entrada_hash1_nonce_20_), .Y(_3528_) );
XNOR2X1 XNOR2X1_212 ( .A(bloque_bytes[52]), .B(bloque_bytes[12]), .Y(_3529_) );
NAND2X1 NAND2X1_654 ( .A(_3529_), .B(_3528_), .Y(micro_ucr_hash1_W_19__4_) );
INVX1 INVX1_532 ( .A(bloque_bytes[77]), .Y(_3530_) );
INVX1 INVX1_533 ( .A(entrada_hash1_nonce_21_), .Y(_3531_) );
OAI21X1 OAI21X1_610 ( .A(_3530_), .B(bloque_bytes[37]), .C(_3531_), .Y(_3532_) );
AOI21X1 AOI21X1_375 ( .A(_3530_), .B(bloque_bytes[37]), .C(_3532_), .Y(_3533_) );
AND2X2 AND2X2_176 ( .A(bloque_bytes[53]), .B(bloque_bytes[13]), .Y(_3534_) );
NOR2X1 NOR2X1_408 ( .A(bloque_bytes[53]), .B(bloque_bytes[13]), .Y(_3535_) );
OAI21X1 OAI21X1_611 ( .A(_3534_), .B(_3535_), .C(_3533_), .Y(micro_ucr_hash1_W_19__5_) );
XOR2X1 XOR2X1_297 ( .A(bloque_bytes[54]), .B(bloque_bytes[14]), .Y(_3536_) );
NOR2X1 NOR2X1_409 ( .A(_3536_), .B(micro_ucr_hash1_W_16__6_), .Y(_3537_) );
INVX1 INVX1_534 ( .A(_3537_), .Y(micro_ucr_hash1_W_19__6_) );
INVX1 INVX1_535 ( .A(bloque_bytes[79]), .Y(_3538_) );
NAND2X1 NAND2X1_655 ( .A(bloque_bytes[39]), .B(_3538_), .Y(_3539_) );
AND2X2 AND2X2_177 ( .A(_3484_), .B(_3539_), .Y(_3540_) );
XNOR2X1 XNOR2X1_213 ( .A(bloque_bytes[55]), .B(bloque_bytes[15]), .Y(_3541_) );
NAND2X1 NAND2X1_656 ( .A(_3541_), .B(_3540_), .Y(micro_ucr_hash1_W_19__7_) );
XOR2X1 XOR2X1_298 ( .A(bloque_bytes[64]), .B(bloque_bytes[24]), .Y(_3542_) );
NOR2X1 NOR2X1_410 ( .A(entrada_hash1_nonce_8_), .B(_3542_), .Y(_3543_) );
XNOR2X1 XNOR2X1_214 ( .A(bloque_bytes[40]), .B(bloque_bytes[0]), .Y(_3544_) );
NAND2X1 NAND2X1_657 ( .A(_3544_), .B(_3543_), .Y(micro_ucr_hash1_W_20__0_) );
XOR2X1 XOR2X1_299 ( .A(bloque_bytes[65]), .B(bloque_bytes[25]), .Y(_3545_) );
NOR2X1 NOR2X1_411 ( .A(entrada_hash1_nonce_9_), .B(_3545_), .Y(_3546_) );
XNOR2X1 XNOR2X1_215 ( .A(bloque_bytes[41]), .B(bloque_bytes[1]), .Y(_3547_) );
NAND2X1 NAND2X1_658 ( .A(_3547_), .B(_3546_), .Y(micro_ucr_hash1_W_20__1_) );
INVX1 INVX1_536 ( .A(bloque_bytes[66]), .Y(_3548_) );
INVX1 INVX1_537 ( .A(entrada_hash1_nonce_10_), .Y(_3549_) );
OAI21X1 OAI21X1_612 ( .A(_3548_), .B(bloque_bytes[26]), .C(_3549_), .Y(_3550_) );
AOI21X1 AOI21X1_376 ( .A(_3548_), .B(bloque_bytes[26]), .C(_3550_), .Y(_3551_) );
XNOR2X1 XNOR2X1_216 ( .A(bloque_bytes[42]), .B(bloque_bytes[2]), .Y(_3552_) );
NAND2X1 NAND2X1_659 ( .A(_3552_), .B(_3551_), .Y(micro_ucr_hash1_W_20__2_) );
XOR2X1 XOR2X1_300 ( .A(bloque_bytes[43]), .B(bloque_bytes[3]), .Y(_3553_) );
NOR2X1 NOR2X1_412 ( .A(_3553_), .B(micro_ucr_hash1_W_17__3_), .Y(_3554_) );
INVX1 INVX1_538 ( .A(_3554_), .Y(micro_ucr_hash1_W_20__3_) );
XOR2X1 XOR2X1_301 ( .A(bloque_bytes[44]), .B(bloque_bytes[4]), .Y(_3555_) );
NOR2X1 NOR2X1_413 ( .A(_3555_), .B(micro_ucr_hash1_W_17__4_), .Y(_3556_) );
INVX1 INVX1_539 ( .A(_3556_), .Y(micro_ucr_hash1_W_20__4_) );
XOR2X1 XOR2X1_302 ( .A(bloque_bytes[45]), .B(bloque_bytes[5]), .Y(_3557_) );
NOR2X1 NOR2X1_414 ( .A(_3557_), .B(micro_ucr_hash1_W_17__5_), .Y(_3558_) );
INVX1 INVX1_540 ( .A(_3558_), .Y(micro_ucr_hash1_W_20__5_) );
XOR2X1 XOR2X1_303 ( .A(bloque_bytes[46]), .B(bloque_bytes[6]), .Y(_3559_) );
NOR2X1 NOR2X1_415 ( .A(_3559_), .B(micro_ucr_hash1_W_17__6_), .Y(_3560_) );
INVX1 INVX1_541 ( .A(_3560_), .Y(micro_ucr_hash1_W_20__6_) );
INVX1 INVX1_542 ( .A(bloque_bytes[71]), .Y(_3561_) );
INVX1 INVX1_543 ( .A(entrada_hash1_nonce_15_), .Y(_3562_) );
OAI21X1 OAI21X1_613 ( .A(_3561_), .B(bloque_bytes[31]), .C(_3562_), .Y(_3563_) );
AOI21X1 AOI21X1_377 ( .A(_3561_), .B(bloque_bytes[31]), .C(_3563_), .Y(_3564_) );
XNOR2X1 XNOR2X1_217 ( .A(bloque_bytes[47]), .B(bloque_bytes[7]), .Y(_3565_) );
NAND2X1 NAND2X1_660 ( .A(_3565_), .B(_3564_), .Y(micro_ucr_hash1_W_20__7_) );
AND2X2 AND2X2_178 ( .A(bloque_bytes[32]), .B(entrada_hash1_nonce_24_), .Y(_3566_) );
NOR2X1 NOR2X1_416 ( .A(bloque_bytes[32]), .B(entrada_hash1_nonce_24_), .Y(_3567_) );
OAI21X1 OAI21X1_614 ( .A(_3566_), .B(_3567_), .C(_3488_), .Y(micro_ucr_hash1_W_21__0_) );
AND2X2 AND2X2_179 ( .A(bloque_bytes[33]), .B(entrada_hash1_nonce_25_), .Y(_3568_) );
NOR2X1 NOR2X1_417 ( .A(bloque_bytes[33]), .B(entrada_hash1_nonce_25_), .Y(_3569_) );
OAI21X1 OAI21X1_615 ( .A(_3568_), .B(_3569_), .C(_3492_), .Y(micro_ucr_hash1_W_21__1_) );
INVX1 INVX1_544 ( .A(entrada_hash1_nonce_26_), .Y(_3570_) );
NOR2X1 NOR2X1_418 ( .A(_3469_), .B(_3570_), .Y(_3571_) );
NOR2X1 NOR2X1_419 ( .A(bloque_bytes[34]), .B(entrada_hash1_nonce_26_), .Y(_3572_) );
OAI21X1 OAI21X1_616 ( .A(_3571_), .B(_3572_), .C(_3496_), .Y(micro_ucr_hash1_W_21__2_) );
AND2X2 AND2X2_180 ( .A(bloque_bytes[35]), .B(entrada_hash1_nonce_27_), .Y(_3573_) );
NOR2X1 NOR2X1_420 ( .A(bloque_bytes[35]), .B(entrada_hash1_nonce_27_), .Y(_3574_) );
OAI21X1 OAI21X1_617 ( .A(_3573_), .B(_3574_), .C(_3500_), .Y(micro_ucr_hash1_W_21__3_) );
AND2X2 AND2X2_181 ( .A(bloque_bytes[36]), .B(entrada_hash1_nonce_28_), .Y(_3575_) );
NOR2X1 NOR2X1_421 ( .A(bloque_bytes[36]), .B(entrada_hash1_nonce_28_), .Y(_3576_) );
OAI21X1 OAI21X1_618 ( .A(_3575_), .B(_3576_), .C(_3504_), .Y(micro_ucr_hash1_W_21__4_) );
INVX2 INVX2_88 ( .A(entrada_hash1_nonce_29_), .Y(_3577_) );
NOR2X1 NOR2X1_422 ( .A(_3479_), .B(_3577_), .Y(_3578_) );
NOR2X1 NOR2X1_423 ( .A(bloque_bytes[37]), .B(entrada_hash1_nonce_29_), .Y(_3579_) );
OAI21X1 OAI21X1_619 ( .A(_3578_), .B(_3579_), .C(_3508_), .Y(micro_ucr_hash1_W_21__5_) );
INVX2 INVX2_89 ( .A(entrada_hash1_nonce_30_), .Y(_3580_) );
NOR2X1 NOR2X1_424 ( .A(_3481_), .B(_3580_), .Y(_3581_) );
NOR2X1 NOR2X1_425 ( .A(bloque_bytes[38]), .B(entrada_hash1_nonce_30_), .Y(_3582_) );
OAI21X1 OAI21X1_620 ( .A(_3581_), .B(_3582_), .C(_3512_), .Y(micro_ucr_hash1_W_21__6_) );
XNOR2X1 XNOR2X1_218 ( .A(bloque_bytes[39]), .B(entrada_hash1_nonce_31_), .Y(_3583_) );
AND2X2 AND2X2_182 ( .A(_3516_), .B(_3583_), .Y(_3584_) );
INVX1 INVX1_545 ( .A(_3584_), .Y(micro_ucr_hash1_W_21__7_) );
XNOR2X1 XNOR2X1_219 ( .A(bloque_bytes[24]), .B(entrada_hash1_nonce_16_), .Y(_3585_) );
NAND3X1 NAND3X1_503 ( .A(_3518_), .B(_3585_), .C(_3517_), .Y(micro_ucr_hash1_W_22__0_) );
XNOR2X1 XNOR2X1_220 ( .A(bloque_bytes[25]), .B(entrada_hash1_nonce_17_), .Y(_3586_) );
NAND3X1 NAND3X1_504 ( .A(_3520_), .B(_3586_), .C(_3519_), .Y(micro_ucr_hash1_W_22__1_) );
XNOR2X1 XNOR2X1_221 ( .A(bloque_bytes[26]), .B(entrada_hash1_nonce_18_), .Y(_3587_) );
NAND3X1 NAND3X1_505 ( .A(_3525_), .B(_3587_), .C(_3524_), .Y(micro_ucr_hash1_W_22__2_) );
XNOR2X1 XNOR2X1_222 ( .A(bloque_bytes[27]), .B(entrada_hash1_nonce_19_), .Y(_3588_) );
NAND3X1 NAND3X1_506 ( .A(_3527_), .B(_3588_), .C(_3526_), .Y(micro_ucr_hash1_W_22__3_) );
XNOR2X1 XNOR2X1_223 ( .A(bloque_bytes[28]), .B(entrada_hash1_nonce_20_), .Y(_3589_) );
NAND3X1 NAND3X1_507 ( .A(_3529_), .B(_3589_), .C(_3528_), .Y(micro_ucr_hash1_W_22__4_) );
XOR2X1 XOR2X1_304 ( .A(bloque_bytes[29]), .B(entrada_hash1_nonce_21_), .Y(_3590_) );
NOR2X1 NOR2X1_426 ( .A(_3590_), .B(micro_ucr_hash1_W_19__5_), .Y(_3591_) );
INVX1 INVX1_546 ( .A(_3591_), .Y(micro_ucr_hash1_W_22__5_) );
INVX1 INVX1_547 ( .A(bloque_bytes[78]), .Y(_3592_) );
INVX1 INVX1_548 ( .A(entrada_hash1_nonce_22_), .Y(_3593_) );
OAI21X1 OAI21X1_621 ( .A(_3592_), .B(bloque_bytes[38]), .C(_3593_), .Y(_3594_) );
AOI21X1 AOI21X1_378 ( .A(_3592_), .B(bloque_bytes[38]), .C(_3594_), .Y(_3595_) );
INVX1 INVX1_549 ( .A(_3536_), .Y(_3596_) );
XNOR2X1 XNOR2X1_224 ( .A(bloque_bytes[30]), .B(entrada_hash1_nonce_22_), .Y(_3597_) );
NAND3X1 NAND3X1_508 ( .A(_3596_), .B(_3597_), .C(_3595_), .Y(micro_ucr_hash1_W_22__6_) );
XNOR2X1 XNOR2X1_225 ( .A(bloque_bytes[31]), .B(entrada_hash1_nonce_23_), .Y(_3598_) );
NAND3X1 NAND3X1_509 ( .A(_3541_), .B(_3598_), .C(_3540_), .Y(micro_ucr_hash1_W_22__7_) );
XNOR2X1 XNOR2X1_226 ( .A(entrada_hash1_nonce_8_), .B(bloque_bytes[16]), .Y(_3599_) );
NAND3X1 NAND3X1_510 ( .A(_3544_), .B(_3599_), .C(_3543_), .Y(micro_ucr_hash1_W_23__0_) );
XNOR2X1 XNOR2X1_227 ( .A(entrada_hash1_nonce_9_), .B(bloque_bytes[17]), .Y(_3600_) );
NAND3X1 NAND3X1_511 ( .A(_3547_), .B(_3600_), .C(_3546_), .Y(micro_ucr_hash1_W_23__1_) );
XNOR2X1 XNOR2X1_228 ( .A(entrada_hash1_nonce_10_), .B(bloque_bytes[18]), .Y(_3601_) );
NAND3X1 NAND3X1_512 ( .A(_3552_), .B(_3601_), .C(_3551_), .Y(micro_ucr_hash1_W_23__2_) );
XNOR2X1 XNOR2X1_229 ( .A(entrada_hash1_nonce_11_), .B(bloque_bytes[19]), .Y(_3602_) );
AND2X2 AND2X2_183 ( .A(_3554_), .B(_3602_), .Y(_3603_) );
INVX1 INVX1_550 ( .A(_3603_), .Y(micro_ucr_hash1_W_23__3_) );
XNOR2X1 XNOR2X1_230 ( .A(entrada_hash1_nonce_12_), .B(bloque_bytes[20]), .Y(_3604_) );
AND2X2 AND2X2_184 ( .A(_3556_), .B(_3604_), .Y(_3605_) );
INVX1 INVX1_551 ( .A(_3605_), .Y(micro_ucr_hash1_W_23__4_) );
XNOR2X1 XNOR2X1_231 ( .A(entrada_hash1_nonce_13_), .B(bloque_bytes[21]), .Y(_3606_) );
AND2X2 AND2X2_185 ( .A(_3558_), .B(_3606_), .Y(_3607_) );
INVX1 INVX1_552 ( .A(_3607_), .Y(micro_ucr_hash1_W_23__5_) );
XNOR2X1 XNOR2X1_232 ( .A(entrada_hash1_nonce_14_), .B(bloque_bytes[22]), .Y(_3608_) );
AND2X2 AND2X2_186 ( .A(_3560_), .B(_3608_), .Y(_3609_) );
INVX1 INVX1_553 ( .A(_3609_), .Y(micro_ucr_hash1_W_23__6_) );
XNOR2X1 XNOR2X1_233 ( .A(entrada_hash1_nonce_15_), .B(bloque_bytes[23]), .Y(_3610_) );
NAND3X1 NAND3X1_513 ( .A(_3565_), .B(_3610_), .C(_3564_), .Y(micro_ucr_hash1_W_23__7_) );
OR2X2 OR2X2_135 ( .A(micro_ucr_hash1_W_21__0_), .B(bloque_bytes[8]), .Y(micro_ucr_hash1_W_24__0_) );
OR2X2 OR2X2_136 ( .A(micro_ucr_hash1_W_21__1_), .B(bloque_bytes[9]), .Y(micro_ucr_hash1_W_24__1_) );
NOR2X1 NOR2X1_427 ( .A(bloque_bytes[10]), .B(micro_ucr_hash1_W_21__2_), .Y(_3611_) );
INVX1 INVX1_554 ( .A(_3611_), .Y(micro_ucr_hash1_W_24__2_) );
OR2X2 OR2X2_137 ( .A(micro_ucr_hash1_W_21__3_), .B(bloque_bytes[11]), .Y(micro_ucr_hash1_W_24__3_) );
OR2X2 OR2X2_138 ( .A(micro_ucr_hash1_W_21__4_), .B(bloque_bytes[12]), .Y(micro_ucr_hash1_W_24__4_) );
NOR2X1 NOR2X1_428 ( .A(bloque_bytes[13]), .B(micro_ucr_hash1_W_21__5_), .Y(_3612_) );
INVX1 INVX1_555 ( .A(_3612_), .Y(micro_ucr_hash1_W_24__5_) );
NOR2X1 NOR2X1_429 ( .A(bloque_bytes[14]), .B(micro_ucr_hash1_W_21__6_), .Y(_3613_) );
INVX1 INVX1_556 ( .A(_3613_), .Y(micro_ucr_hash1_W_24__6_) );
AND2X2 AND2X2_187 ( .A(entrada_hash1_nonce_7_), .B(bloque_bytes[15]), .Y(_3614_) );
NOR2X1 NOR2X1_430 ( .A(entrada_hash1_nonce_7_), .B(bloque_bytes[15]), .Y(_3615_) );
OAI21X1 OAI21X1_622 ( .A(_3614_), .B(_3615_), .C(_3584_), .Y(micro_ucr_hash1_W_24__7_) );
NAND2X1 NAND2X1_661 ( .A(bloque_bytes[0]), .B(micro_ucr_hash1_W_16__0_), .Y(_3616_) );
INVX1 INVX1_557 ( .A(bloque_bytes[0]), .Y(_3617_) );
NAND2X1 NAND2X1_662 ( .A(_3617_), .B(_3517_), .Y(_3618_) );
AOI21X1 AOI21X1_379 ( .A(_3618_), .B(_3616_), .C(micro_ucr_hash1_W_22__0_), .Y(_3619_) );
INVX1 INVX1_558 ( .A(_3619_), .Y(micro_ucr_hash1_W_25__0_) );
NAND2X1 NAND2X1_663 ( .A(bloque_bytes[1]), .B(micro_ucr_hash1_W_16__1_), .Y(_3620_) );
INVX1 INVX1_559 ( .A(bloque_bytes[1]), .Y(_3621_) );
NAND2X1 NAND2X1_664 ( .A(_3621_), .B(_3519_), .Y(_3622_) );
AOI21X1 AOI21X1_380 ( .A(_3622_), .B(_3620_), .C(micro_ucr_hash1_W_22__1_), .Y(_3623_) );
INVX1 INVX1_560 ( .A(_3623_), .Y(micro_ucr_hash1_W_25__1_) );
NAND2X1 NAND2X1_665 ( .A(bloque_bytes[2]), .B(micro_ucr_hash1_W_16__2_), .Y(_3624_) );
OR2X2 OR2X2_139 ( .A(micro_ucr_hash1_W_16__2_), .B(bloque_bytes[2]), .Y(_3625_) );
AOI21X1 AOI21X1_381 ( .A(_3624_), .B(_3625_), .C(micro_ucr_hash1_W_22__2_), .Y(_3626_) );
INVX1 INVX1_561 ( .A(_3626_), .Y(micro_ucr_hash1_W_25__2_) );
NAND2X1 NAND2X1_666 ( .A(bloque_bytes[3]), .B(micro_ucr_hash1_W_16__3_), .Y(_3627_) );
INVX1 INVX1_562 ( .A(bloque_bytes[3]), .Y(_3628_) );
NAND2X1 NAND2X1_667 ( .A(_3628_), .B(_3526_), .Y(_3629_) );
AOI21X1 AOI21X1_382 ( .A(_3629_), .B(_3627_), .C(micro_ucr_hash1_W_22__3_), .Y(_3630_) );
INVX1 INVX1_563 ( .A(_3630_), .Y(micro_ucr_hash1_W_25__3_) );
NAND2X1 NAND2X1_668 ( .A(bloque_bytes[4]), .B(micro_ucr_hash1_W_16__4_), .Y(_3631_) );
INVX1 INVX1_564 ( .A(bloque_bytes[4]), .Y(_3632_) );
NAND2X1 NAND2X1_669 ( .A(_3632_), .B(_3528_), .Y(_3633_) );
AOI21X1 AOI21X1_383 ( .A(_3633_), .B(_3631_), .C(micro_ucr_hash1_W_22__4_), .Y(_3634_) );
INVX1 INVX1_565 ( .A(_3634_), .Y(micro_ucr_hash1_W_25__4_) );
XNOR2X1 XNOR2X1_234 ( .A(micro_ucr_hash1_W_16__5_), .B(bloque_bytes[5]), .Y(_3635_) );
NAND2X1 NAND2X1_670 ( .A(_3635_), .B(_3591_), .Y(micro_ucr_hash1_W_25__5_) );
NAND2X1 NAND2X1_671 ( .A(bloque_bytes[6]), .B(micro_ucr_hash1_W_16__6_), .Y(_3636_) );
OR2X2 OR2X2_140 ( .A(micro_ucr_hash1_W_16__6_), .B(bloque_bytes[6]), .Y(_3637_) );
AOI21X1 AOI21X1_384 ( .A(_3636_), .B(_3637_), .C(micro_ucr_hash1_W_22__6_), .Y(_3638_) );
INVX1 INVX1_566 ( .A(_3638_), .Y(micro_ucr_hash1_W_25__6_) );
NAND2X1 NAND2X1_672 ( .A(bloque_bytes[7]), .B(micro_ucr_hash1_W_16__7_), .Y(_3639_) );
OR2X2 OR2X2_141 ( .A(micro_ucr_hash1_W_16__7_), .B(bloque_bytes[7]), .Y(_3640_) );
AOI21X1 AOI21X1_385 ( .A(_3639_), .B(_3640_), .C(micro_ucr_hash1_W_22__7_), .Y(_3641_) );
INVX1 INVX1_567 ( .A(_3641_), .Y(micro_ucr_hash1_W_25__7_) );
OAI21X1 OAI21X1_623 ( .A(_3542_), .B(entrada_hash1_nonce_8_), .C(entrada_hash1_nonce_24_), .Y(_3642_) );
OR2X2 OR2X2_142 ( .A(micro_ucr_hash1_W_17__0_), .B(entrada_hash1_nonce_24_), .Y(_3643_) );
AOI21X1 AOI21X1_386 ( .A(_3642_), .B(_3643_), .C(micro_ucr_hash1_W_23__0_), .Y(_3644_) );
INVX1 INVX1_568 ( .A(_3644_), .Y(micro_ucr_hash1_W_26__0_) );
OAI21X1 OAI21X1_624 ( .A(_3545_), .B(entrada_hash1_nonce_9_), .C(entrada_hash1_nonce_25_), .Y(_3645_) );
OR2X2 OR2X2_143 ( .A(micro_ucr_hash1_W_17__1_), .B(entrada_hash1_nonce_25_), .Y(_3646_) );
AOI21X1 AOI21X1_387 ( .A(_3645_), .B(_3646_), .C(micro_ucr_hash1_W_23__1_), .Y(_3647_) );
INVX1 INVX1_569 ( .A(_3647_), .Y(micro_ucr_hash1_W_26__1_) );
NAND2X1 NAND2X1_673 ( .A(entrada_hash1_nonce_26_), .B(micro_ucr_hash1_W_17__2_), .Y(_3648_) );
NAND2X1 NAND2X1_674 ( .A(_3570_), .B(_3551_), .Y(_3649_) );
AOI21X1 AOI21X1_388 ( .A(_3648_), .B(_3649_), .C(micro_ucr_hash1_W_23__2_), .Y(_3650_) );
INVX1 INVX1_570 ( .A(_3650_), .Y(micro_ucr_hash1_W_26__2_) );
INVX1 INVX1_571 ( .A(entrada_hash1_nonce_27_), .Y(_3651_) );
NAND2X1 NAND2X1_675 ( .A(_3651_), .B(_3603_), .Y(micro_ucr_hash1_W_26__3_) );
INVX1 INVX1_572 ( .A(entrada_hash1_nonce_28_), .Y(_3652_) );
NAND2X1 NAND2X1_676 ( .A(_3652_), .B(_3605_), .Y(micro_ucr_hash1_W_26__4_) );
NAND2X1 NAND2X1_677 ( .A(_3577_), .B(_3607_), .Y(micro_ucr_hash1_W_26__5_) );
NAND2X1 NAND2X1_678 ( .A(_3580_), .B(_3609_), .Y(micro_ucr_hash1_W_26__6_) );
NAND2X1 NAND2X1_679 ( .A(entrada_hash1_nonce_31_), .B(micro_ucr_hash1_W_17__7_), .Y(_3653_) );
OR2X2 OR2X2_144 ( .A(micro_ucr_hash1_W_17__7_), .B(entrada_hash1_nonce_31_), .Y(_3654_) );
AOI21X1 AOI21X1_389 ( .A(_3653_), .B(_3654_), .C(micro_ucr_hash1_W_23__7_), .Y(_3655_) );
INVX1 INVX1_573 ( .A(_3655_), .Y(micro_ucr_hash1_W_26__7_) );
OR2X2 OR2X2_145 ( .A(micro_ucr_hash1_W_24__0_), .B(entrada_hash1_nonce_16_), .Y(micro_ucr_hash1_W_27__0_) );
OR2X2 OR2X2_146 ( .A(micro_ucr_hash1_W_24__1_), .B(entrada_hash1_nonce_17_), .Y(micro_ucr_hash1_W_27__1_) );
NAND2X1 NAND2X1_680 ( .A(_3522_), .B(_3611_), .Y(micro_ucr_hash1_W_27__2_) );
OR2X2 OR2X2_147 ( .A(micro_ucr_hash1_W_24__3_), .B(entrada_hash1_nonce_19_), .Y(micro_ucr_hash1_W_27__3_) );
OR2X2 OR2X2_148 ( .A(micro_ucr_hash1_W_24__4_), .B(entrada_hash1_nonce_20_), .Y(micro_ucr_hash1_W_27__4_) );
NAND2X1 NAND2X1_681 ( .A(_3531_), .B(_3612_), .Y(micro_ucr_hash1_W_27__5_) );
NAND2X1 NAND2X1_682 ( .A(_3593_), .B(_3613_), .Y(micro_ucr_hash1_W_27__6_) );
OR2X2 OR2X2_149 ( .A(micro_ucr_hash1_W_24__7_), .B(entrada_hash1_nonce_23_), .Y(micro_ucr_hash1_W_27__7_) );
XNOR2X1 XNOR2X1_235 ( .A(micro_ucr_hash1_W_19__0_), .B(entrada_hash1_nonce_8_), .Y(_3656_) );
NAND2X1 NAND2X1_683 ( .A(_3619_), .B(_3656_), .Y(micro_ucr_hash1_W_28__0_) );
XNOR2X1 XNOR2X1_236 ( .A(micro_ucr_hash1_W_19__1_), .B(entrada_hash1_nonce_9_), .Y(_3657_) );
NAND2X1 NAND2X1_684 ( .A(_3623_), .B(_3657_), .Y(micro_ucr_hash1_W_28__1_) );
NAND2X1 NAND2X1_685 ( .A(_3549_), .B(_3626_), .Y(micro_ucr_hash1_W_28__2_) );
XNOR2X1 XNOR2X1_237 ( .A(micro_ucr_hash1_W_19__3_), .B(entrada_hash1_nonce_11_), .Y(_3658_) );
NAND2X1 NAND2X1_686 ( .A(_3630_), .B(_3658_), .Y(micro_ucr_hash1_W_28__3_) );
XNOR2X1 XNOR2X1_238 ( .A(micro_ucr_hash1_W_19__4_), .B(entrada_hash1_nonce_12_), .Y(_3659_) );
NAND2X1 NAND2X1_687 ( .A(_3634_), .B(_3659_), .Y(micro_ucr_hash1_W_28__4_) );
INVX1 INVX1_574 ( .A(entrada_hash1_nonce_13_), .Y(_3660_) );
NAND3X1 NAND3X1_514 ( .A(_3660_), .B(_3635_), .C(_3591_), .Y(micro_ucr_hash1_W_28__5_) );
OAI21X1 OAI21X1_625 ( .A(micro_ucr_hash1_W_16__6_), .B(_3536_), .C(entrada_hash1_nonce_14_), .Y(_3661_) );
INVX1 INVX1_575 ( .A(entrada_hash1_nonce_14_), .Y(_3662_) );
NAND3X1 NAND3X1_515 ( .A(_3662_), .B(_3596_), .C(_3595_), .Y(_3663_) );
NAND2X1 NAND2X1_688 ( .A(_3661_), .B(_3663_), .Y(_3664_) );
NAND2X1 NAND2X1_689 ( .A(_3664_), .B(_3638_), .Y(micro_ucr_hash1_W_28__6_) );
NAND2X1 NAND2X1_690 ( .A(_3562_), .B(_3641_), .Y(micro_ucr_hash1_W_28__7_) );
AOI21X1 AOI21X1_390 ( .A(_3544_), .B(_3543_), .C(_3486_), .Y(_3665_) );
NOR2X1 NOR2X1_431 ( .A(entrada_hash1_nonce_0_), .B(micro_ucr_hash1_W_20__0_), .Y(_3666_) );
OAI21X1 OAI21X1_626 ( .A(_3666_), .B(_3665_), .C(_3644_), .Y(micro_ucr_hash1_W_29__0_) );
AOI21X1 AOI21X1_391 ( .A(_3547_), .B(_3546_), .C(_3490_), .Y(_3667_) );
NOR2X1 NOR2X1_432 ( .A(entrada_hash1_nonce_1_), .B(micro_ucr_hash1_W_20__1_), .Y(_3668_) );
OAI21X1 OAI21X1_627 ( .A(_3668_), .B(_3667_), .C(_3647_), .Y(micro_ucr_hash1_W_29__1_) );
AOI21X1 AOI21X1_392 ( .A(_3552_), .B(_3551_), .C(_3494_), .Y(_3669_) );
NOR2X1 NOR2X1_433 ( .A(entrada_hash1_nonce_2_), .B(micro_ucr_hash1_W_20__2_), .Y(_3670_) );
OAI21X1 OAI21X1_628 ( .A(_3670_), .B(_3669_), .C(_3650_), .Y(micro_ucr_hash1_W_29__2_) );
NAND3X1 NAND3X1_516 ( .A(_3498_), .B(_3651_), .C(_3603_), .Y(micro_ucr_hash1_W_29__3_) );
NAND3X1 NAND3X1_517 ( .A(_3502_), .B(_3652_), .C(_3605_), .Y(micro_ucr_hash1_W_29__4_) );
NAND3X1 NAND3X1_518 ( .A(_3506_), .B(_3577_), .C(_3607_), .Y(micro_ucr_hash1_W_29__5_) );
NAND3X1 NAND3X1_519 ( .A(_3510_), .B(_3580_), .C(_3609_), .Y(micro_ucr_hash1_W_29__6_) );
AOI21X1 AOI21X1_393 ( .A(_3565_), .B(_3564_), .C(_3514_), .Y(_3671_) );
NOR2X1 NOR2X1_434 ( .A(entrada_hash1_nonce_7_), .B(micro_ucr_hash1_W_20__7_), .Y(_3672_) );
OAI21X1 OAI21X1_629 ( .A(_3671_), .B(_3672_), .C(_3655_), .Y(micro_ucr_hash1_W_29__7_) );
OR2X2 OR2X2_150 ( .A(micro_ucr_hash1_W_24__0_), .B(micro_ucr_hash1_W_16__0_), .Y(micro_ucr_hash1_W_30__0_) );
OR2X2 OR2X2_151 ( .A(micro_ucr_hash1_W_24__1_), .B(micro_ucr_hash1_W_16__1_), .Y(micro_ucr_hash1_W_30__1_) );
NAND2X1 NAND2X1_691 ( .A(_3524_), .B(_3611_), .Y(micro_ucr_hash1_W_30__2_) );
OR2X2 OR2X2_152 ( .A(micro_ucr_hash1_W_24__3_), .B(micro_ucr_hash1_W_16__3_), .Y(micro_ucr_hash1_W_30__3_) );
OR2X2 OR2X2_153 ( .A(micro_ucr_hash1_W_24__4_), .B(micro_ucr_hash1_W_16__4_), .Y(micro_ucr_hash1_W_30__4_) );
NAND2X1 NAND2X1_692 ( .A(_3533_), .B(_3612_), .Y(micro_ucr_hash1_W_30__5_) );
NAND2X1 NAND2X1_693 ( .A(_3595_), .B(_3613_), .Y(micro_ucr_hash1_W_30__6_) );
OR2X2 OR2X2_154 ( .A(micro_ucr_hash1_W_24__7_), .B(micro_ucr_hash1_W_16__7_), .Y(micro_ucr_hash1_W_30__7_) );
XNOR2X1 XNOR2X1_239 ( .A(micro_ucr_hash1_W_22__0_), .B(micro_ucr_hash1_W_17__0_), .Y(_3673_) );
NAND3X1 NAND3X1_520 ( .A(_3619_), .B(_3656_), .C(_3673_), .Y(micro_ucr_hash1_W_31__0_) );
XNOR2X1 XNOR2X1_240 ( .A(micro_ucr_hash1_W_22__1_), .B(micro_ucr_hash1_W_17__1_), .Y(_3674_) );
NAND3X1 NAND3X1_521 ( .A(_3623_), .B(_3657_), .C(_3674_), .Y(micro_ucr_hash1_W_31__1_) );
NAND3X1 NAND3X1_522 ( .A(_3549_), .B(_3551_), .C(_3626_), .Y(micro_ucr_hash1_W_31__2_) );
XNOR2X1 XNOR2X1_241 ( .A(micro_ucr_hash1_W_22__3_), .B(micro_ucr_hash1_W_17__3_), .Y(_3675_) );
NAND3X1 NAND3X1_523 ( .A(_3630_), .B(_3658_), .C(_3675_), .Y(micro_ucr_hash1_W_31__3_) );
XNOR2X1 XNOR2X1_242 ( .A(micro_ucr_hash1_W_22__4_), .B(micro_ucr_hash1_W_17__4_), .Y(_3676_) );
NAND3X1 NAND3X1_524 ( .A(_3634_), .B(_3659_), .C(_3676_), .Y(micro_ucr_hash1_W_31__4_) );
INVX1 INVX1_576 ( .A(micro_ucr_hash1_W_17__5_), .Y(_3677_) );
NAND3X1 NAND3X1_525 ( .A(_3677_), .B(_3635_), .C(_3591_), .Y(micro_ucr_hash1_W_31__5_) );
INVX1 INVX1_577 ( .A(micro_ucr_hash1_W_17__6_), .Y(_3678_) );
NAND3X1 NAND3X1_526 ( .A(_3678_), .B(_3664_), .C(_3638_), .Y(micro_ucr_hash1_W_31__6_) );
NAND3X1 NAND3X1_527 ( .A(_3562_), .B(_3564_), .C(_3641_), .Y(micro_ucr_hash1_W_31__7_) );
INVX1 INVX1_578 ( .A(gnd), .Y(_3444__8_) );
NAND2X1 NAND2X1_694 ( .A(gnd), .B(gnd), .Y(_3679_) );
INVX1 INVX1_579 ( .A(_3679_), .Y(_3680_) );
NOR2X1 NOR2X1_435 ( .A(gnd), .B(gnd), .Y(_3681_) );
NOR2X1 NOR2X1_436 ( .A(_3681_), .B(_3680_), .Y(_3444__9_) );
XNOR2X1 XNOR2X1_243 ( .A(_3679_), .B(gnd), .Y(_3444__10_) );
INVX2 INVX2_90 ( .A(gnd), .Y(_3682_) );
NAND2X1 NAND2X1_695 ( .A(gnd), .B(_3680_), .Y(_3683_) );
XNOR2X1 XNOR2X1_244 ( .A(_3683_), .B(_3682_), .Y(_3444__11_) );
INVX1 INVX1_580 ( .A(gnd), .Y(_3684_) );
OAI21X1 OAI21X1_630 ( .A(_3679_), .B(_3684_), .C(_3682_), .Y(_3685_) );
XOR2X1 XOR2X1_305 ( .A(_3685_), .B(micro_ucr_hash1_b_31__4_), .Y(_3444__12_) );
AND2X2 AND2X2_188 ( .A(_3685_), .B(micro_ucr_hash1_b_31__4_), .Y(_3686_) );
AND2X2 AND2X2_189 ( .A(_3686_), .B(micro_ucr_hash1_b_31__5_), .Y(_3687_) );
NOR2X1 NOR2X1_437 ( .A(micro_ucr_hash1_b_31__5_), .B(_3686_), .Y(_3688_) );
NOR2X1 NOR2X1_438 ( .A(_3688_), .B(_3687_), .Y(_3444__13_) );
XOR2X1 XOR2X1_306 ( .A(_3687_), .B(micro_ucr_hash1_b_31__6_), .Y(_3444__14_) );
NAND3X1 NAND3X1_528 ( .A(micro_ucr_hash1_b_31__5_), .B(micro_ucr_hash1_b_31__6_), .C(_3686_), .Y(_3689_) );
XOR2X1 XOR2X1_307 ( .A(_3689_), .B(micro_ucr_hash1_b_31__7_), .Y(_3444__15_) );
AND2X2 AND2X2_190 ( .A(micro_ucr_hash1_a_31__0_), .B(micro_ucr_hash1_a_31__1_), .Y(_3690_) );
NOR2X1 NOR2X1_439 ( .A(micro_ucr_hash1_a_31__0_), .B(micro_ucr_hash1_a_31__1_), .Y(_3691_) );
NOR2X1 NOR2X1_440 ( .A(_3691_), .B(_3690_), .Y(_3444__17_) );
INVX2 INVX2_91 ( .A(micro_ucr_hash1_a_31__2_), .Y(_3692_) );
XNOR2X1 XNOR2X1_245 ( .A(_3690_), .B(_3692_), .Y(_3444__18_) );
NAND2X1 NAND2X1_696 ( .A(micro_ucr_hash1_a_31__2_), .B(_3690_), .Y(_3693_) );
XNOR2X1 XNOR2X1_246 ( .A(_3693_), .B(micro_ucr_hash1_a_31__3_), .Y(_3444__19_) );
INVX1 INVX1_581 ( .A(micro_ucr_hash1_a_31__3_), .Y(_3694_) );
NOR2X1 NOR2X1_441 ( .A(_3692_), .B(_3694_), .Y(_3695_) );
NAND3X1 NAND3X1_529 ( .A(micro_ucr_hash1_a_31__4_), .B(_3690_), .C(_3695_), .Y(_3696_) );
INVX1 INVX1_582 ( .A(micro_ucr_hash1_a_31__4_), .Y(_3697_) );
OAI21X1 OAI21X1_631 ( .A(_3693_), .B(_3694_), .C(_3697_), .Y(_3698_) );
AND2X2 AND2X2_191 ( .A(_3698_), .B(_3696_), .Y(_3444__20_) );
XNOR2X1 XNOR2X1_247 ( .A(_3696_), .B(micro_ucr_hash1_a_31__5_), .Y(_3444__21_) );
AND2X2 AND2X2_192 ( .A(micro_ucr_hash1_a_31__4_), .B(micro_ucr_hash1_a_31__5_), .Y(_3699_) );
NAND3X1 NAND3X1_530 ( .A(_3690_), .B(_3699_), .C(_3695_), .Y(_3700_) );
XNOR2X1 XNOR2X1_248 ( .A(_3700_), .B(micro_ucr_hash1_a_31__6_), .Y(_3444__22_) );
INVX1 INVX1_583 ( .A(micro_ucr_hash1_a_31__6_), .Y(_3701_) );
NOR2X1 NOR2X1_442 ( .A(_3701_), .B(_3700_), .Y(_3702_) );
XOR2X1 XOR2X1_308 ( .A(_3702_), .B(micro_ucr_hash1_a_31__7_), .Y(_3444__23_) );
INVX1 INVX1_584 ( .A(micro_ucr_hash1_a_31__0_), .Y(_3444__16_) );
INVX1 INVX1_585 ( .A(micro_ucr_hash1_c_31__1_), .Y(_3444__1_) );
NOR2X1 NOR2X1_443 ( .A(micro_ucr_hash1_c_31__1_), .B(micro_ucr_hash1_c_31__2_), .Y(_3703_) );
INVX1 INVX1_586 ( .A(_3703_), .Y(_3704_) );
NAND2X1 NAND2X1_697 ( .A(micro_ucr_hash1_c_31__1_), .B(micro_ucr_hash1_c_31__2_), .Y(_3705_) );
NAND2X1 NAND2X1_698 ( .A(_3705_), .B(_3704_), .Y(_3444__2_) );
OAI21X1 OAI21X1_632 ( .A(micro_ucr_hash1_c_31__1_), .B(micro_ucr_hash1_c_31__2_), .C(micro_ucr_hash1_c_31__3_), .Y(_3706_) );
INVX1 INVX1_587 ( .A(micro_ucr_hash1_c_31__3_), .Y(_3707_) );
NAND2X1 NAND2X1_699 ( .A(_3707_), .B(_3703_), .Y(_3708_) );
NAND2X1 NAND2X1_700 ( .A(_3706_), .B(_3708_), .Y(_3444__3_) );
INVX1 INVX1_588 ( .A(micro_ucr_hash1_c_31__4_), .Y(_3709_) );
NAND3X1 NAND3X1_531 ( .A(_3707_), .B(_3709_), .C(_3703_), .Y(_3710_) );
OAI21X1 OAI21X1_633 ( .A(_3704_), .B(micro_ucr_hash1_c_31__3_), .C(micro_ucr_hash1_c_31__4_), .Y(_3711_) );
NAND2X1 NAND2X1_701 ( .A(_3710_), .B(_3711_), .Y(_3444__4_) );
XNOR2X1 XNOR2X1_249 ( .A(_3710_), .B(micro_ucr_hash1_c_31__5_), .Y(_3444__5_) );
INVX1 INVX1_589 ( .A(micro_ucr_hash1_c_31__6_), .Y(_3712_) );
NOR2X1 NOR2X1_444 ( .A(micro_ucr_hash1_c_31__5_), .B(_3710_), .Y(_3713_) );
NAND2X1 NAND2X1_702 ( .A(_3712_), .B(_3713_), .Y(_3714_) );
OAI21X1 OAI21X1_634 ( .A(_3710_), .B(micro_ucr_hash1_c_31__5_), .C(micro_ucr_hash1_c_31__6_), .Y(_3715_) );
NAND2X1 NAND2X1_703 ( .A(_3715_), .B(_3714_), .Y(_3444__6_) );
XNOR2X1 XNOR2X1_250 ( .A(_3714_), .B(micro_ucr_hash1_c_31__7_), .Y(_3444__7_) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf8), .D(micro_ucr_hash1_c_31__0_), .Q(micro_ucr_hash1_hash_0_) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf8), .D(_3444__1_), .Q(micro_ucr_hash1_hash_1_) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf8), .D(_3444__2_), .Q(micro_ucr_hash1_hash_2_) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf8), .D(_3444__3_), .Q(micro_ucr_hash1_hash_3_) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf8), .D(_3444__4_), .Q(micro_ucr_hash1_hash_4_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf8), .D(_3444__5_), .Q(micro_ucr_hash1_hash_5_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf8), .D(_3444__6_), .Q(micro_ucr_hash1_hash_6_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf8), .D(_3444__7_), .Q(micro_ucr_hash1_hash_7_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf2), .D(_3444__8_), .Q(micro_ucr_hash1_hash_8_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf2), .D(_3444__9_), .Q(micro_ucr_hash1_hash_9_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf2), .D(_3444__10_), .Q(micro_ucr_hash1_hash_10_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf4), .D(_3444__11_), .Q(micro_ucr_hash1_hash_11_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf1), .D(_3444__12_), .Q(micro_ucr_hash1_hash_12_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf0), .D(_3444__13_), .Q(micro_ucr_hash1_hash_13_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf2), .D(_3444__14_), .Q(micro_ucr_hash1_hash_14_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf0), .D(_3444__15_), .Q(micro_ucr_hash1_hash_15_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf4), .D(_3444__16_), .Q(micro_ucr_hash1_hash_16_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf0), .D(_3444__17_), .Q(micro_ucr_hash1_hash_17_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf6), .D(_3444__18_), .Q(micro_ucr_hash1_hash_18_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf6), .D(_3444__19_), .Q(micro_ucr_hash1_hash_19_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf6), .D(_3444__20_), .Q(micro_ucr_hash1_hash_20_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf6), .D(_3444__21_), .Q(micro_ucr_hash1_hash_21_) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf6), .D(_3444__22_), .Q(micro_ucr_hash1_hash_22_) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf6), .D(_3444__23_), .Q(micro_ucr_hash1_hash_23_) );
XOR2X1 XOR2X1_309 ( .A(gnd), .B(vdd), .Y(micro_ucr_hash1_a_0__0_) );
XOR2X1 XOR2X1_310 ( .A(vdd), .B(gnd), .Y(micro_ucr_hash1_a_0__1_) );
XOR2X1 XOR2X1_311 ( .A(vdd), .B(gnd), .Y(micro_ucr_hash1_a_0__2_) );
XOR2X1 XOR2X1_312 ( .A(vdd), .B(vdd), .Y(micro_ucr_hash1_a_0__3_) );
XOR2X1 XOR2X1_313 ( .A(vdd), .B(gnd), .Y(micro_ucr_hash1_a_0__4_) );
XOR2X1 XOR2X1_314 ( .A(vdd), .B(gnd), .Y(micro_ucr_hash1_a_0__5_) );
XOR2X1 XOR2X1_315 ( .A(vdd), .B(gnd), .Y(micro_ucr_hash1_a_0__6_) );
XOR2X1 XOR2X1_316 ( .A(vdd), .B(vdd), .Y(micro_ucr_hash1_a_0__7_) );
INVX2 INVX2_92 ( .A(bloque_bytes[88]), .Y(_3785_) );
XNOR2X1 XNOR2X1_251 ( .A(vdd), .B(vdd), .Y(_3786_) );
XNOR2X1 XNOR2X1_252 ( .A(_3786_), .B(_3785_), .Y(micro_ucr_hash1_b_1__4_) );
NAND2X1 NAND2X1_704 ( .A(_3785_), .B(_3786_), .Y(_3787_) );
OR2X2 OR2X2_155 ( .A(gnd), .B(gnd), .Y(_3788_) );
NAND2X1 NAND2X1_705 ( .A(gnd), .B(gnd), .Y(_3789_) );
NAND3X1 NAND3X1_532 ( .A(bloque_bytes[89]), .B(_3789_), .C(_3788_), .Y(_3790_) );
INVX1 INVX1_590 ( .A(bloque_bytes[89]), .Y(_3791_) );
NOR2X1 NOR2X1_445 ( .A(gnd), .B(gnd), .Y(_3792_) );
AND2X2 AND2X2_193 ( .A(gnd), .B(gnd), .Y(_3793_) );
OAI21X1 OAI21X1_635 ( .A(_3793_), .B(_3792_), .C(_3791_), .Y(_3794_) );
NAND2X1 NAND2X1_706 ( .A(_3794_), .B(_3790_), .Y(_3795_) );
XNOR2X1 XNOR2X1_253 ( .A(_3795_), .B(_3787_), .Y(micro_ucr_hash1_b_1__5_) );
NAND3X1 NAND3X1_533 ( .A(_3790_), .B(_3794_), .C(_3787_), .Y(_3796_) );
NOR3X1 NOR3X1_97 ( .A(_3791_), .B(_3792_), .C(_3793_), .Y(_3797_) );
INVX1 INVX1_591 ( .A(bloque_bytes[90]), .Y(_3798_) );
NOR2X1 NOR2X1_446 ( .A(gnd), .B(gnd), .Y(_3799_) );
AND2X2 AND2X2_194 ( .A(gnd), .B(gnd), .Y(_3800_) );
NOR3X1 NOR3X1_98 ( .A(_3798_), .B(_3799_), .C(_3800_), .Y(_3801_) );
OR2X2 OR2X2_156 ( .A(gnd), .B(gnd), .Y(_3802_) );
NAND2X1 NAND2X1_707 ( .A(gnd), .B(gnd), .Y(_3803_) );
AOI21X1 AOI21X1_394 ( .A(_3803_), .B(_3802_), .C(bloque_bytes[90]), .Y(_3804_) );
OAI21X1 OAI21X1_636 ( .A(_3801_), .B(_3804_), .C(_3797_), .Y(_3805_) );
NAND3X1 NAND3X1_534 ( .A(bloque_bytes[90]), .B(_3803_), .C(_3802_), .Y(_3806_) );
OAI21X1 OAI21X1_637 ( .A(_3800_), .B(_3799_), .C(_3798_), .Y(_3807_) );
NAND3X1 NAND3X1_535 ( .A(_3807_), .B(_3790_), .C(_3806_), .Y(_3808_) );
NAND2X1 NAND2X1_708 ( .A(_3808_), .B(_3805_), .Y(_3809_) );
XNOR2X1 XNOR2X1_254 ( .A(_3809_), .B(_3796_), .Y(micro_ucr_hash1_b_1__6_) );
NAND3X1 NAND3X1_536 ( .A(_3806_), .B(_3807_), .C(_3797_), .Y(_3810_) );
OAI21X1 OAI21X1_638 ( .A(_3801_), .B(_3804_), .C(_3790_), .Y(_3811_) );
NAND2X1 NAND2X1_709 ( .A(_3810_), .B(_3811_), .Y(_3812_) );
OAI21X1 OAI21X1_639 ( .A(_3812_), .B(_3796_), .C(_3810_), .Y(_3813_) );
INVX1 INVX1_592 ( .A(bloque_bytes[91]), .Y(_3814_) );
NOR2X1 NOR2X1_447 ( .A(vdd), .B(gnd), .Y(_3815_) );
AND2X2 AND2X2_195 ( .A(vdd), .B(gnd), .Y(_3816_) );
OAI21X1 OAI21X1_640 ( .A(_3816_), .B(_3815_), .C(_3814_), .Y(_3817_) );
OR2X2 OR2X2_157 ( .A(vdd), .B(gnd), .Y(_3818_) );
NAND2X1 NAND2X1_710 ( .A(vdd), .B(gnd), .Y(_3819_) );
NAND3X1 NAND3X1_537 ( .A(bloque_bytes[91]), .B(_3819_), .C(_3818_), .Y(_3820_) );
AOI21X1 AOI21X1_395 ( .A(_3817_), .B(_3820_), .C(_3806_), .Y(_3821_) );
NAND3X1 NAND3X1_538 ( .A(_3814_), .B(_3819_), .C(_3818_), .Y(_3822_) );
OAI21X1 OAI21X1_641 ( .A(_3816_), .B(_3815_), .C(bloque_bytes[91]), .Y(_3823_) );
AOI21X1 AOI21X1_396 ( .A(_3823_), .B(_3822_), .C(_3801_), .Y(_3824_) );
NOR2X1 NOR2X1_448 ( .A(_3821_), .B(_3824_), .Y(_3716_) );
XOR2X1 XOR2X1_317 ( .A(_3813_), .B(_3716_), .Y(micro_ucr_hash1_b_1__7_) );
INVX1 INVX1_593 ( .A(bloque_bytes[92]), .Y(_3717_) );
OR2X2 OR2X2_158 ( .A(gnd), .B(gnd), .Y(_3718_) );
NAND2X1 NAND2X1_711 ( .A(gnd), .B(gnd), .Y(_3719_) );
NAND3X1 NAND3X1_539 ( .A(_3717_), .B(_3719_), .C(_3718_), .Y(_3720_) );
NOR2X1 NOR2X1_449 ( .A(gnd), .B(gnd), .Y(_3721_) );
AND2X2 AND2X2_196 ( .A(gnd), .B(gnd), .Y(_3722_) );
OAI21X1 OAI21X1_642 ( .A(_3722_), .B(_3721_), .C(bloque_bytes[92]), .Y(_3723_) );
NAND3X1 NAND3X1_540 ( .A(_3817_), .B(_3720_), .C(_3723_), .Y(_3724_) );
AOI21X1 AOI21X1_397 ( .A(_3819_), .B(_3818_), .C(bloque_bytes[91]), .Y(_3725_) );
OAI21X1 OAI21X1_643 ( .A(_3722_), .B(_3721_), .C(_3717_), .Y(_3726_) );
NAND3X1 NAND3X1_541 ( .A(bloque_bytes[92]), .B(_3719_), .C(_3718_), .Y(_3727_) );
NAND3X1 NAND3X1_542 ( .A(_3726_), .B(_3727_), .C(_3725_), .Y(_3728_) );
AND2X2 AND2X2_197 ( .A(_3728_), .B(_3724_), .Y(_3729_) );
INVX2 INVX2_93 ( .A(_3824_), .Y(_3730_) );
NOR2X1 NOR2X1_450 ( .A(_3804_), .B(_3801_), .Y(_3731_) );
AOI21X1 AOI21X1_398 ( .A(_3797_), .B(_3731_), .C(_3821_), .Y(_3732_) );
OAI21X1 OAI21X1_644 ( .A(_3812_), .B(_3796_), .C(_3732_), .Y(_3733_) );
NAND2X1 NAND2X1_712 ( .A(_3730_), .B(_3733_), .Y(_3734_) );
XNOR2X1 XNOR2X1_255 ( .A(_3734_), .B(_3729_), .Y(micro_ucr_hash1_c_0__4_) );
NAND2X1 NAND2X1_713 ( .A(_3724_), .B(_3728_), .Y(_3735_) );
OAI21X1 OAI21X1_645 ( .A(_3734_), .B(_3735_), .C(_3724_), .Y(_3736_) );
INVX1 INVX1_594 ( .A(bloque_bytes[93]), .Y(_3737_) );
OR2X2 OR2X2_159 ( .A(gnd), .B(gnd), .Y(_3738_) );
NAND2X1 NAND2X1_714 ( .A(gnd), .B(gnd), .Y(_3739_) );
NAND3X1 NAND3X1_543 ( .A(_3737_), .B(_3739_), .C(_3738_), .Y(_3740_) );
NOR2X1 NOR2X1_451 ( .A(gnd), .B(gnd), .Y(_3741_) );
AND2X2 AND2X2_198 ( .A(gnd), .B(gnd), .Y(_3742_) );
OAI21X1 OAI21X1_646 ( .A(_3742_), .B(_3741_), .C(bloque_bytes[93]), .Y(_3743_) );
NAND3X1 NAND3X1_544 ( .A(_3726_), .B(_3743_), .C(_3740_), .Y(_3744_) );
AOI21X1 AOI21X1_399 ( .A(_3719_), .B(_3718_), .C(bloque_bytes[92]), .Y(_3745_) );
NAND3X1 NAND3X1_545 ( .A(bloque_bytes[93]), .B(_3739_), .C(_3738_), .Y(_3746_) );
OAI21X1 OAI21X1_647 ( .A(_3742_), .B(_3741_), .C(_3737_), .Y(_3747_) );
NAND3X1 NAND3X1_546 ( .A(_3747_), .B(_3746_), .C(_3745_), .Y(_3748_) );
NAND2X1 NAND2X1_715 ( .A(_3744_), .B(_3748_), .Y(_3749_) );
INVX2 INVX2_94 ( .A(_3749_), .Y(_3750_) );
XNOR2X1 XNOR2X1_256 ( .A(_3736_), .B(_3750_), .Y(micro_ucr_hash1_c_0__5_) );
AOI21X1 AOI21X1_400 ( .A(_3744_), .B(_3748_), .C(_3735_), .Y(_3751_) );
NAND3X1 NAND3X1_547 ( .A(_3730_), .B(_3751_), .C(_3733_), .Y(_3752_) );
NAND2X1 NAND2X1_716 ( .A(_3747_), .B(_3746_), .Y(_3753_) );
OR2X2 OR2X2_160 ( .A(_3753_), .B(_3745_), .Y(_3754_) );
INVX1 INVX1_595 ( .A(_3754_), .Y(_3755_) );
AOI21X1 AOI21X1_401 ( .A(_3745_), .B(_3753_), .C(_3724_), .Y(_3756_) );
NOR2X1 NOR2X1_452 ( .A(_3756_), .B(_3755_), .Y(_3757_) );
INVX1 INVX1_596 ( .A(bloque_bytes[94]), .Y(_3758_) );
XNOR2X1 XNOR2X1_257 ( .A(gnd), .B(gnd), .Y(_3759_) );
OR2X2 OR2X2_161 ( .A(_3759_), .B(_3758_), .Y(_3760_) );
NAND2X1 NAND2X1_717 ( .A(_3758_), .B(_3759_), .Y(_3761_) );
NAND2X1 NAND2X1_718 ( .A(_3761_), .B(_3760_), .Y(_3762_) );
OR2X2 OR2X2_162 ( .A(_3762_), .B(_3746_), .Y(_3763_) );
NAND2X1 NAND2X1_719 ( .A(_3746_), .B(_3762_), .Y(_3764_) );
NAND2X1 NAND2X1_720 ( .A(_3764_), .B(_3763_), .Y(_3765_) );
AOI21X1 AOI21X1_402 ( .A(_3757_), .B(_3752_), .C(_3765_), .Y(_3766_) );
NAND2X1 NAND2X1_721 ( .A(_3749_), .B(_3729_), .Y(_3767_) );
OAI21X1 OAI21X1_648 ( .A(_3734_), .B(_3767_), .C(_3757_), .Y(_3768_) );
INVX1 INVX1_597 ( .A(_3765_), .Y(_3769_) );
NOR2X1 NOR2X1_453 ( .A(_3769_), .B(_3768_), .Y(_3770_) );
NOR2X1 NOR2X1_454 ( .A(_3766_), .B(_3770_), .Y(micro_ucr_hash1_c_0__6_) );
INVX1 INVX1_598 ( .A(_3810_), .Y(_3771_) );
AOI21X1 AOI21X1_403 ( .A(_3730_), .B(_3771_), .C(_3821_), .Y(_3772_) );
AOI21X1 AOI21X1_404 ( .A(_3785_), .B(_3786_), .C(_3795_), .Y(_3773_) );
NAND3X1 NAND3X1_548 ( .A(_3773_), .B(_3809_), .C(_3716_), .Y(_3774_) );
AOI21X1 AOI21X1_405 ( .A(_3772_), .B(_3774_), .C(_3767_), .Y(_3775_) );
OAI21X1 OAI21X1_649 ( .A(_3750_), .B(_3724_), .C(_3754_), .Y(_3776_) );
OAI21X1 OAI21X1_650 ( .A(_3775_), .B(_3776_), .C(_3769_), .Y(_3777_) );
XOR2X1 XOR2X1_318 ( .A(vdd), .B(bloque_bytes[95]), .Y(_3778_) );
XNOR2X1 XNOR2X1_258 ( .A(_3778_), .B(gnd), .Y(_3779_) );
XNOR2X1 XNOR2X1_259 ( .A(_3779_), .B(_3760_), .Y(_3780_) );
NAND3X1 NAND3X1_549 ( .A(_3763_), .B(_3780_), .C(_3777_), .Y(_3781_) );
INVX1 INVX1_599 ( .A(_3763_), .Y(_3782_) );
INVX1 INVX1_600 ( .A(_3780_), .Y(_3783_) );
OAI21X1 OAI21X1_651 ( .A(_3766_), .B(_3782_), .C(_3783_), .Y(_3784_) );
NAND2X1 NAND2X1_722 ( .A(_3781_), .B(_3784_), .Y(micro_ucr_hash1_c_0__7_) );
BUFX2 BUFX2_26 ( .A(micro_ucr_hash1_c_31__0_), .Y(_3444__0_) );
BUFX2 BUFX2_27 ( .A(gnd), .Y(micro_ucr_hash1_b_10__0_) );
BUFX2 BUFX2_28 ( .A(gnd), .Y(micro_ucr_hash1_b_10__1_) );
BUFX2 BUFX2_29 ( .A(gnd), .Y(micro_ucr_hash1_b_10__2_) );
BUFX2 BUFX2_30 ( .A(gnd), .Y(micro_ucr_hash1_b_10__3_) );
BUFX2 BUFX2_31 ( .A(gnd), .Y(micro_ucr_hash1_b_11__0_) );
BUFX2 BUFX2_32 ( .A(gnd), .Y(micro_ucr_hash1_b_11__1_) );
BUFX2 BUFX2_33 ( .A(gnd), .Y(micro_ucr_hash1_b_11__2_) );
BUFX2 BUFX2_34 ( .A(gnd), .Y(micro_ucr_hash1_b_11__3_) );
BUFX2 BUFX2_35 ( .A(gnd), .Y(micro_ucr_hash1_b_12__0_) );
BUFX2 BUFX2_36 ( .A(gnd), .Y(micro_ucr_hash1_b_12__1_) );
BUFX2 BUFX2_37 ( .A(gnd), .Y(micro_ucr_hash1_b_12__2_) );
BUFX2 BUFX2_38 ( .A(gnd), .Y(micro_ucr_hash1_b_12__3_) );
BUFX2 BUFX2_39 ( .A(gnd), .Y(micro_ucr_hash1_b_13__0_) );
BUFX2 BUFX2_40 ( .A(gnd), .Y(micro_ucr_hash1_b_13__1_) );
BUFX2 BUFX2_41 ( .A(gnd), .Y(micro_ucr_hash1_b_13__2_) );
BUFX2 BUFX2_42 ( .A(gnd), .Y(micro_ucr_hash1_b_13__3_) );
BUFX2 BUFX2_43 ( .A(gnd), .Y(micro_ucr_hash1_b_14__0_) );
BUFX2 BUFX2_44 ( .A(gnd), .Y(micro_ucr_hash1_b_14__1_) );
BUFX2 BUFX2_45 ( .A(gnd), .Y(micro_ucr_hash1_b_14__2_) );
BUFX2 BUFX2_46 ( .A(gnd), .Y(micro_ucr_hash1_b_14__3_) );
BUFX2 BUFX2_47 ( .A(gnd), .Y(micro_ucr_hash1_b_15__0_) );
BUFX2 BUFX2_48 ( .A(gnd), .Y(micro_ucr_hash1_b_15__1_) );
BUFX2 BUFX2_49 ( .A(gnd), .Y(micro_ucr_hash1_b_15__2_) );
BUFX2 BUFX2_50 ( .A(gnd), .Y(micro_ucr_hash1_b_15__3_) );
BUFX2 BUFX2_51 ( .A(gnd), .Y(micro_ucr_hash1_b_16__0_) );
BUFX2 BUFX2_52 ( .A(gnd), .Y(micro_ucr_hash1_b_16__1_) );
BUFX2 BUFX2_53 ( .A(gnd), .Y(micro_ucr_hash1_b_16__2_) );
BUFX2 BUFX2_54 ( .A(gnd), .Y(micro_ucr_hash1_b_16__3_) );
BUFX2 BUFX2_55 ( .A(gnd), .Y(micro_ucr_hash1_b_17__0_) );
BUFX2 BUFX2_56 ( .A(gnd), .Y(micro_ucr_hash1_b_17__1_) );
BUFX2 BUFX2_57 ( .A(gnd), .Y(micro_ucr_hash1_b_17__2_) );
BUFX2 BUFX2_58 ( .A(gnd), .Y(micro_ucr_hash1_b_17__3_) );
BUFX2 BUFX2_59 ( .A(gnd), .Y(micro_ucr_hash1_b_18__0_) );
BUFX2 BUFX2_60 ( .A(gnd), .Y(micro_ucr_hash1_b_18__1_) );
BUFX2 BUFX2_61 ( .A(gnd), .Y(micro_ucr_hash1_b_18__2_) );
BUFX2 BUFX2_62 ( .A(gnd), .Y(micro_ucr_hash1_b_18__3_) );
BUFX2 BUFX2_63 ( .A(gnd), .Y(micro_ucr_hash1_b_19__0_) );
BUFX2 BUFX2_64 ( .A(gnd), .Y(micro_ucr_hash1_b_19__1_) );
BUFX2 BUFX2_65 ( .A(gnd), .Y(micro_ucr_hash1_b_19__2_) );
BUFX2 BUFX2_66 ( .A(gnd), .Y(micro_ucr_hash1_b_19__3_) );
BUFX2 BUFX2_67 ( .A(gnd), .Y(micro_ucr_hash1_b_1__0_) );
BUFX2 BUFX2_68 ( .A(gnd), .Y(micro_ucr_hash1_b_1__1_) );
BUFX2 BUFX2_69 ( .A(gnd), .Y(micro_ucr_hash1_b_1__2_) );
BUFX2 BUFX2_70 ( .A(gnd), .Y(micro_ucr_hash1_b_1__3_) );
BUFX2 BUFX2_71 ( .A(gnd), .Y(micro_ucr_hash1_b_20__0_) );
BUFX2 BUFX2_72 ( .A(gnd), .Y(micro_ucr_hash1_b_20__1_) );
BUFX2 BUFX2_73 ( .A(gnd), .Y(micro_ucr_hash1_b_20__2_) );
BUFX2 BUFX2_74 ( .A(gnd), .Y(micro_ucr_hash1_b_20__3_) );
BUFX2 BUFX2_75 ( .A(gnd), .Y(micro_ucr_hash1_b_21__0_) );
BUFX2 BUFX2_76 ( .A(gnd), .Y(micro_ucr_hash1_b_21__1_) );
BUFX2 BUFX2_77 ( .A(gnd), .Y(micro_ucr_hash1_b_21__2_) );
BUFX2 BUFX2_78 ( .A(gnd), .Y(micro_ucr_hash1_b_21__3_) );
BUFX2 BUFX2_79 ( .A(gnd), .Y(micro_ucr_hash1_b_22__0_) );
BUFX2 BUFX2_80 ( .A(gnd), .Y(micro_ucr_hash1_b_22__1_) );
BUFX2 BUFX2_81 ( .A(gnd), .Y(micro_ucr_hash1_b_22__2_) );
BUFX2 BUFX2_82 ( .A(gnd), .Y(micro_ucr_hash1_b_22__3_) );
BUFX2 BUFX2_83 ( .A(gnd), .Y(micro_ucr_hash1_b_23__0_) );
BUFX2 BUFX2_84 ( .A(gnd), .Y(micro_ucr_hash1_b_23__1_) );
BUFX2 BUFX2_85 ( .A(gnd), .Y(micro_ucr_hash1_b_23__2_) );
BUFX2 BUFX2_86 ( .A(gnd), .Y(micro_ucr_hash1_b_23__3_) );
BUFX2 BUFX2_87 ( .A(gnd), .Y(micro_ucr_hash1_b_24__0_) );
BUFX2 BUFX2_88 ( .A(gnd), .Y(micro_ucr_hash1_b_24__1_) );
BUFX2 BUFX2_89 ( .A(gnd), .Y(micro_ucr_hash1_b_24__2_) );
BUFX2 BUFX2_90 ( .A(gnd), .Y(micro_ucr_hash1_b_24__3_) );
BUFX2 BUFX2_91 ( .A(gnd), .Y(micro_ucr_hash1_b_25__0_) );
BUFX2 BUFX2_92 ( .A(gnd), .Y(micro_ucr_hash1_b_25__1_) );
BUFX2 BUFX2_93 ( .A(gnd), .Y(micro_ucr_hash1_b_25__2_) );
BUFX2 BUFX2_94 ( .A(gnd), .Y(micro_ucr_hash1_b_25__3_) );
BUFX2 BUFX2_95 ( .A(gnd), .Y(micro_ucr_hash1_b_26__0_) );
BUFX2 BUFX2_96 ( .A(gnd), .Y(micro_ucr_hash1_b_26__1_) );
BUFX2 BUFX2_97 ( .A(gnd), .Y(micro_ucr_hash1_b_26__2_) );
BUFX2 BUFX2_98 ( .A(gnd), .Y(micro_ucr_hash1_b_26__3_) );
BUFX2 BUFX2_99 ( .A(gnd), .Y(micro_ucr_hash1_b_27__0_) );
BUFX2 BUFX2_100 ( .A(gnd), .Y(micro_ucr_hash1_b_27__1_) );
BUFX2 BUFX2_101 ( .A(gnd), .Y(micro_ucr_hash1_b_27__2_) );
BUFX2 BUFX2_102 ( .A(gnd), .Y(micro_ucr_hash1_b_27__3_) );
BUFX2 BUFX2_103 ( .A(gnd), .Y(micro_ucr_hash1_b_28__0_) );
BUFX2 BUFX2_104 ( .A(gnd), .Y(micro_ucr_hash1_b_28__1_) );
BUFX2 BUFX2_105 ( .A(gnd), .Y(micro_ucr_hash1_b_28__2_) );
BUFX2 BUFX2_106 ( .A(gnd), .Y(micro_ucr_hash1_b_28__3_) );
BUFX2 BUFX2_107 ( .A(gnd), .Y(micro_ucr_hash1_b_29__0_) );
BUFX2 BUFX2_108 ( .A(gnd), .Y(micro_ucr_hash1_b_29__1_) );
BUFX2 BUFX2_109 ( .A(gnd), .Y(micro_ucr_hash1_b_29__2_) );
BUFX2 BUFX2_110 ( .A(gnd), .Y(micro_ucr_hash1_b_29__3_) );
BUFX2 BUFX2_111 ( .A(gnd), .Y(micro_ucr_hash1_b_2__0_) );
BUFX2 BUFX2_112 ( .A(gnd), .Y(micro_ucr_hash1_b_2__1_) );
BUFX2 BUFX2_113 ( .A(gnd), .Y(micro_ucr_hash1_b_2__2_) );
BUFX2 BUFX2_114 ( .A(gnd), .Y(micro_ucr_hash1_b_2__3_) );
BUFX2 BUFX2_115 ( .A(gnd), .Y(micro_ucr_hash1_b_30__0_) );
BUFX2 BUFX2_116 ( .A(gnd), .Y(micro_ucr_hash1_b_30__1_) );
BUFX2 BUFX2_117 ( .A(gnd), .Y(micro_ucr_hash1_b_30__2_) );
BUFX2 BUFX2_118 ( .A(gnd), .Y(micro_ucr_hash1_b_30__3_) );
BUFX2 BUFX2_119 ( .A(gnd), .Y(micro_ucr_hash1_b_31__0_) );
BUFX2 BUFX2_120 ( .A(gnd), .Y(micro_ucr_hash1_b_31__1_) );
BUFX2 BUFX2_121 ( .A(gnd), .Y(micro_ucr_hash1_b_31__2_) );
BUFX2 BUFX2_122 ( .A(gnd), .Y(micro_ucr_hash1_b_31__3_) );
BUFX2 BUFX2_123 ( .A(gnd), .Y(micro_ucr_hash1_b_3__0_) );
BUFX2 BUFX2_124 ( .A(gnd), .Y(micro_ucr_hash1_b_3__1_) );
BUFX2 BUFX2_125 ( .A(gnd), .Y(micro_ucr_hash1_b_3__2_) );
BUFX2 BUFX2_126 ( .A(gnd), .Y(micro_ucr_hash1_b_3__3_) );
BUFX2 BUFX2_127 ( .A(gnd), .Y(micro_ucr_hash1_b_4__0_) );
BUFX2 BUFX2_128 ( .A(gnd), .Y(micro_ucr_hash1_b_4__1_) );
BUFX2 BUFX2_129 ( .A(gnd), .Y(micro_ucr_hash1_b_4__2_) );
BUFX2 BUFX2_130 ( .A(gnd), .Y(micro_ucr_hash1_b_4__3_) );
BUFX2 BUFX2_131 ( .A(gnd), .Y(micro_ucr_hash1_b_5__0_) );
BUFX2 BUFX2_132 ( .A(gnd), .Y(micro_ucr_hash1_b_5__1_) );
BUFX2 BUFX2_133 ( .A(gnd), .Y(micro_ucr_hash1_b_5__2_) );
BUFX2 BUFX2_134 ( .A(gnd), .Y(micro_ucr_hash1_b_5__3_) );
BUFX2 BUFX2_135 ( .A(gnd), .Y(micro_ucr_hash1_b_6__0_) );
BUFX2 BUFX2_136 ( .A(gnd), .Y(micro_ucr_hash1_b_6__1_) );
BUFX2 BUFX2_137 ( .A(gnd), .Y(micro_ucr_hash1_b_6__2_) );
BUFX2 BUFX2_138 ( .A(gnd), .Y(micro_ucr_hash1_b_6__3_) );
BUFX2 BUFX2_139 ( .A(gnd), .Y(micro_ucr_hash1_b_7__0_) );
BUFX2 BUFX2_140 ( .A(gnd), .Y(micro_ucr_hash1_b_7__1_) );
BUFX2 BUFX2_141 ( .A(gnd), .Y(micro_ucr_hash1_b_7__2_) );
BUFX2 BUFX2_142 ( .A(gnd), .Y(micro_ucr_hash1_b_7__3_) );
BUFX2 BUFX2_143 ( .A(gnd), .Y(micro_ucr_hash1_b_8__0_) );
BUFX2 BUFX2_144 ( .A(gnd), .Y(micro_ucr_hash1_b_8__1_) );
BUFX2 BUFX2_145 ( .A(gnd), .Y(micro_ucr_hash1_b_8__2_) );
BUFX2 BUFX2_146 ( .A(gnd), .Y(micro_ucr_hash1_b_8__3_) );
BUFX2 BUFX2_147 ( .A(gnd), .Y(micro_ucr_hash1_b_9__0_) );
BUFX2 BUFX2_148 ( .A(gnd), .Y(micro_ucr_hash1_b_9__1_) );
BUFX2 BUFX2_149 ( .A(gnd), .Y(micro_ucr_hash1_b_9__2_) );
BUFX2 BUFX2_150 ( .A(gnd), .Y(micro_ucr_hash1_b_9__3_) );
BUFX2 BUFX2_151 ( .A(micro_ucr_hash1_b_1__4_), .Y(micro_ucr_hash1_c_0__0_) );
BUFX2 BUFX2_152 ( .A(micro_ucr_hash1_b_1__5_), .Y(micro_ucr_hash1_c_0__1_) );
BUFX2 BUFX2_153 ( .A(micro_ucr_hash1_b_1__6_), .Y(micro_ucr_hash1_c_0__2_) );
BUFX2 BUFX2_154 ( .A(micro_ucr_hash1_b_1__7_), .Y(micro_ucr_hash1_c_0__3_) );
BUFX2 BUFX2_155 ( .A(micro_ucr_hash1_b_11__4_), .Y(micro_ucr_hash1_c_10__0_) );
BUFX2 BUFX2_156 ( .A(micro_ucr_hash1_b_11__5_), .Y(micro_ucr_hash1_c_10__1_) );
BUFX2 BUFX2_157 ( .A(micro_ucr_hash1_b_11__6_), .Y(micro_ucr_hash1_c_10__2_) );
BUFX2 BUFX2_158 ( .A(micro_ucr_hash1_b_11__7_), .Y(micro_ucr_hash1_c_10__3_) );
BUFX2 BUFX2_159 ( .A(micro_ucr_hash1_b_12__4_), .Y(micro_ucr_hash1_c_11__0_) );
BUFX2 BUFX2_160 ( .A(micro_ucr_hash1_b_12__5_), .Y(micro_ucr_hash1_c_11__1_) );
BUFX2 BUFX2_161 ( .A(micro_ucr_hash1_b_12__6_), .Y(micro_ucr_hash1_c_11__2_) );
BUFX2 BUFX2_162 ( .A(micro_ucr_hash1_b_12__7_), .Y(micro_ucr_hash1_c_11__3_) );
BUFX2 BUFX2_163 ( .A(micro_ucr_hash1_b_13__4_), .Y(micro_ucr_hash1_c_12__0_) );
BUFX2 BUFX2_164 ( .A(micro_ucr_hash1_b_13__5_), .Y(micro_ucr_hash1_c_12__1_) );
BUFX2 BUFX2_165 ( .A(micro_ucr_hash1_b_13__6_), .Y(micro_ucr_hash1_c_12__2_) );
BUFX2 BUFX2_166 ( .A(micro_ucr_hash1_b_13__7_), .Y(micro_ucr_hash1_c_12__3_) );
BUFX2 BUFX2_167 ( .A(micro_ucr_hash1_b_14__4_), .Y(micro_ucr_hash1_c_13__0_) );
BUFX2 BUFX2_168 ( .A(micro_ucr_hash1_b_14__5_), .Y(micro_ucr_hash1_c_13__1_) );
BUFX2 BUFX2_169 ( .A(micro_ucr_hash1_b_14__6_), .Y(micro_ucr_hash1_c_13__2_) );
BUFX2 BUFX2_170 ( .A(micro_ucr_hash1_b_14__7_), .Y(micro_ucr_hash1_c_13__3_) );
BUFX2 BUFX2_171 ( .A(micro_ucr_hash1_b_15__4_), .Y(micro_ucr_hash1_c_14__0_) );
BUFX2 BUFX2_172 ( .A(micro_ucr_hash1_b_15__5_), .Y(micro_ucr_hash1_c_14__1_) );
BUFX2 BUFX2_173 ( .A(micro_ucr_hash1_b_15__6_), .Y(micro_ucr_hash1_c_14__2_) );
BUFX2 BUFX2_174 ( .A(micro_ucr_hash1_b_15__7_), .Y(micro_ucr_hash1_c_14__3_) );
BUFX2 BUFX2_175 ( .A(micro_ucr_hash1_b_16__4_), .Y(micro_ucr_hash1_c_15__0_) );
BUFX2 BUFX2_176 ( .A(micro_ucr_hash1_b_16__5_), .Y(micro_ucr_hash1_c_15__1_) );
BUFX2 BUFX2_177 ( .A(micro_ucr_hash1_b_16__6_), .Y(micro_ucr_hash1_c_15__2_) );
BUFX2 BUFX2_178 ( .A(micro_ucr_hash1_b_16__7_), .Y(micro_ucr_hash1_c_15__3_) );
BUFX2 BUFX2_179 ( .A(micro_ucr_hash1_b_17__4_), .Y(micro_ucr_hash1_c_16__0_) );
BUFX2 BUFX2_180 ( .A(micro_ucr_hash1_b_17__5_), .Y(micro_ucr_hash1_c_16__1_) );
BUFX2 BUFX2_181 ( .A(micro_ucr_hash1_b_17__6_), .Y(micro_ucr_hash1_c_16__2_) );
BUFX2 BUFX2_182 ( .A(micro_ucr_hash1_b_17__7_), .Y(micro_ucr_hash1_c_16__3_) );
BUFX2 BUFX2_183 ( .A(micro_ucr_hash1_b_18__4_), .Y(micro_ucr_hash1_c_17__0_) );
BUFX2 BUFX2_184 ( .A(micro_ucr_hash1_b_18__5_), .Y(micro_ucr_hash1_c_17__1_) );
BUFX2 BUFX2_185 ( .A(micro_ucr_hash1_b_18__6_), .Y(micro_ucr_hash1_c_17__2_) );
BUFX2 BUFX2_186 ( .A(micro_ucr_hash1_b_18__7_), .Y(micro_ucr_hash1_c_17__3_) );
BUFX2 BUFX2_187 ( .A(micro_ucr_hash1_b_19__4_), .Y(micro_ucr_hash1_c_18__0_) );
BUFX2 BUFX2_188 ( .A(micro_ucr_hash1_b_19__5_), .Y(micro_ucr_hash1_c_18__1_) );
BUFX2 BUFX2_189 ( .A(micro_ucr_hash1_b_19__6_), .Y(micro_ucr_hash1_c_18__2_) );
BUFX2 BUFX2_190 ( .A(micro_ucr_hash1_b_19__7_), .Y(micro_ucr_hash1_c_18__3_) );
BUFX2 BUFX2_191 ( .A(micro_ucr_hash1_b_20__4_), .Y(micro_ucr_hash1_c_19__0_) );
BUFX2 BUFX2_192 ( .A(micro_ucr_hash1_b_20__5_), .Y(micro_ucr_hash1_c_19__1_) );
BUFX2 BUFX2_193 ( .A(micro_ucr_hash1_b_20__6_), .Y(micro_ucr_hash1_c_19__2_) );
BUFX2 BUFX2_194 ( .A(micro_ucr_hash1_b_20__7_), .Y(micro_ucr_hash1_c_19__3_) );
BUFX2 BUFX2_195 ( .A(micro_ucr_hash1_b_2__4_), .Y(micro_ucr_hash1_c_1__0_) );
BUFX2 BUFX2_196 ( .A(micro_ucr_hash1_b_2__5_), .Y(micro_ucr_hash1_c_1__1_) );
BUFX2 BUFX2_197 ( .A(micro_ucr_hash1_b_2__6_), .Y(micro_ucr_hash1_c_1__2_) );
BUFX2 BUFX2_198 ( .A(micro_ucr_hash1_b_2__7_), .Y(micro_ucr_hash1_c_1__3_) );
BUFX2 BUFX2_199 ( .A(micro_ucr_hash1_b_21__4_), .Y(micro_ucr_hash1_c_20__0_) );
BUFX2 BUFX2_200 ( .A(micro_ucr_hash1_b_21__5_), .Y(micro_ucr_hash1_c_20__1_) );
BUFX2 BUFX2_201 ( .A(micro_ucr_hash1_b_21__6_), .Y(micro_ucr_hash1_c_20__2_) );
BUFX2 BUFX2_202 ( .A(micro_ucr_hash1_b_21__7_), .Y(micro_ucr_hash1_c_20__3_) );
BUFX2 BUFX2_203 ( .A(micro_ucr_hash1_b_22__4_), .Y(micro_ucr_hash1_c_21__0_) );
BUFX2 BUFX2_204 ( .A(micro_ucr_hash1_b_22__5_), .Y(micro_ucr_hash1_c_21__1_) );
BUFX2 BUFX2_205 ( .A(micro_ucr_hash1_b_22__6_), .Y(micro_ucr_hash1_c_21__2_) );
BUFX2 BUFX2_206 ( .A(micro_ucr_hash1_b_22__7_), .Y(micro_ucr_hash1_c_21__3_) );
BUFX2 BUFX2_207 ( .A(micro_ucr_hash1_b_23__4_), .Y(micro_ucr_hash1_c_22__0_) );
BUFX2 BUFX2_208 ( .A(micro_ucr_hash1_b_23__5_), .Y(micro_ucr_hash1_c_22__1_) );
BUFX2 BUFX2_209 ( .A(micro_ucr_hash1_b_23__6_), .Y(micro_ucr_hash1_c_22__2_) );
BUFX2 BUFX2_210 ( .A(micro_ucr_hash1_b_23__7_), .Y(micro_ucr_hash1_c_22__3_) );
BUFX2 BUFX2_211 ( .A(micro_ucr_hash1_b_24__4_), .Y(micro_ucr_hash1_c_23__0_) );
BUFX2 BUFX2_212 ( .A(micro_ucr_hash1_b_24__5_), .Y(micro_ucr_hash1_c_23__1_) );
BUFX2 BUFX2_213 ( .A(micro_ucr_hash1_b_24__6_), .Y(micro_ucr_hash1_c_23__2_) );
BUFX2 BUFX2_214 ( .A(micro_ucr_hash1_b_24__7_), .Y(micro_ucr_hash1_c_23__3_) );
BUFX2 BUFX2_215 ( .A(micro_ucr_hash1_b_25__4_), .Y(micro_ucr_hash1_c_24__0_) );
BUFX2 BUFX2_216 ( .A(micro_ucr_hash1_b_25__5_), .Y(micro_ucr_hash1_c_24__1_) );
BUFX2 BUFX2_217 ( .A(micro_ucr_hash1_b_25__6_), .Y(micro_ucr_hash1_c_24__2_) );
BUFX2 BUFX2_218 ( .A(micro_ucr_hash1_b_25__7_), .Y(micro_ucr_hash1_c_24__3_) );
BUFX2 BUFX2_219 ( .A(micro_ucr_hash1_b_26__4_), .Y(micro_ucr_hash1_c_25__0_) );
BUFX2 BUFX2_220 ( .A(micro_ucr_hash1_b_26__5_), .Y(micro_ucr_hash1_c_25__1_) );
BUFX2 BUFX2_221 ( .A(micro_ucr_hash1_b_26__6_), .Y(micro_ucr_hash1_c_25__2_) );
BUFX2 BUFX2_222 ( .A(micro_ucr_hash1_b_26__7_), .Y(micro_ucr_hash1_c_25__3_) );
BUFX2 BUFX2_223 ( .A(micro_ucr_hash1_b_27__4_), .Y(micro_ucr_hash1_c_26__0_) );
BUFX2 BUFX2_224 ( .A(micro_ucr_hash1_b_27__5_), .Y(micro_ucr_hash1_c_26__1_) );
BUFX2 BUFX2_225 ( .A(micro_ucr_hash1_b_27__6_), .Y(micro_ucr_hash1_c_26__2_) );
BUFX2 BUFX2_226 ( .A(micro_ucr_hash1_b_27__7_), .Y(micro_ucr_hash1_c_26__3_) );
BUFX2 BUFX2_227 ( .A(micro_ucr_hash1_b_28__4_), .Y(micro_ucr_hash1_c_27__0_) );
BUFX2 BUFX2_228 ( .A(micro_ucr_hash1_b_28__5_), .Y(micro_ucr_hash1_c_27__1_) );
BUFX2 BUFX2_229 ( .A(micro_ucr_hash1_b_28__6_), .Y(micro_ucr_hash1_c_27__2_) );
BUFX2 BUFX2_230 ( .A(micro_ucr_hash1_b_28__7_), .Y(micro_ucr_hash1_c_27__3_) );
BUFX2 BUFX2_231 ( .A(micro_ucr_hash1_b_29__4_), .Y(micro_ucr_hash1_c_28__0_) );
BUFX2 BUFX2_232 ( .A(micro_ucr_hash1_b_29__5_), .Y(micro_ucr_hash1_c_28__1_) );
BUFX2 BUFX2_233 ( .A(micro_ucr_hash1_b_29__6_), .Y(micro_ucr_hash1_c_28__2_) );
BUFX2 BUFX2_234 ( .A(micro_ucr_hash1_b_29__7_), .Y(micro_ucr_hash1_c_28__3_) );
BUFX2 BUFX2_235 ( .A(micro_ucr_hash1_b_30__4_), .Y(micro_ucr_hash1_c_29__0_) );
BUFX2 BUFX2_236 ( .A(micro_ucr_hash1_b_30__5_), .Y(micro_ucr_hash1_c_29__1_) );
BUFX2 BUFX2_237 ( .A(micro_ucr_hash1_b_30__6_), .Y(micro_ucr_hash1_c_29__2_) );
BUFX2 BUFX2_238 ( .A(micro_ucr_hash1_b_30__7_), .Y(micro_ucr_hash1_c_29__3_) );
BUFX2 BUFX2_239 ( .A(micro_ucr_hash1_b_3__4_), .Y(micro_ucr_hash1_c_2__0_) );
BUFX2 BUFX2_240 ( .A(micro_ucr_hash1_b_3__5_), .Y(micro_ucr_hash1_c_2__1_) );
BUFX2 BUFX2_241 ( .A(micro_ucr_hash1_b_3__6_), .Y(micro_ucr_hash1_c_2__2_) );
BUFX2 BUFX2_242 ( .A(micro_ucr_hash1_b_3__7_), .Y(micro_ucr_hash1_c_2__3_) );
BUFX2 BUFX2_243 ( .A(micro_ucr_hash1_b_31__4_), .Y(micro_ucr_hash1_c_30__0_) );
BUFX2 BUFX2_244 ( .A(micro_ucr_hash1_b_31__5_), .Y(micro_ucr_hash1_c_30__1_) );
BUFX2 BUFX2_245 ( .A(micro_ucr_hash1_b_31__6_), .Y(micro_ucr_hash1_c_30__2_) );
BUFX2 BUFX2_246 ( .A(micro_ucr_hash1_b_31__7_), .Y(micro_ucr_hash1_c_30__3_) );
BUFX2 BUFX2_247 ( .A(micro_ucr_hash1_b_4__4_), .Y(micro_ucr_hash1_c_3__0_) );
BUFX2 BUFX2_248 ( .A(micro_ucr_hash1_b_4__5_), .Y(micro_ucr_hash1_c_3__1_) );
BUFX2 BUFX2_249 ( .A(micro_ucr_hash1_b_4__6_), .Y(micro_ucr_hash1_c_3__2_) );
BUFX2 BUFX2_250 ( .A(micro_ucr_hash1_b_4__7_), .Y(micro_ucr_hash1_c_3__3_) );
BUFX2 BUFX2_251 ( .A(micro_ucr_hash1_b_5__4_), .Y(micro_ucr_hash1_c_4__0_) );
BUFX2 BUFX2_252 ( .A(micro_ucr_hash1_b_5__5_), .Y(micro_ucr_hash1_c_4__1_) );
BUFX2 BUFX2_253 ( .A(micro_ucr_hash1_b_5__6_), .Y(micro_ucr_hash1_c_4__2_) );
BUFX2 BUFX2_254 ( .A(micro_ucr_hash1_b_5__7_), .Y(micro_ucr_hash1_c_4__3_) );
BUFX2 BUFX2_255 ( .A(micro_ucr_hash1_b_6__4_), .Y(micro_ucr_hash1_c_5__0_) );
BUFX2 BUFX2_256 ( .A(micro_ucr_hash1_b_6__5_), .Y(micro_ucr_hash1_c_5__1_) );
BUFX2 BUFX2_257 ( .A(micro_ucr_hash1_b_6__6_), .Y(micro_ucr_hash1_c_5__2_) );
BUFX2 BUFX2_258 ( .A(micro_ucr_hash1_b_6__7_), .Y(micro_ucr_hash1_c_5__3_) );
BUFX2 BUFX2_259 ( .A(micro_ucr_hash1_b_7__4_), .Y(micro_ucr_hash1_c_6__0_) );
BUFX2 BUFX2_260 ( .A(micro_ucr_hash1_b_7__5_), .Y(micro_ucr_hash1_c_6__1_) );
BUFX2 BUFX2_261 ( .A(micro_ucr_hash1_b_7__6_), .Y(micro_ucr_hash1_c_6__2_) );
BUFX2 BUFX2_262 ( .A(micro_ucr_hash1_b_7__7_), .Y(micro_ucr_hash1_c_6__3_) );
BUFX2 BUFX2_263 ( .A(micro_ucr_hash1_b_8__4_), .Y(micro_ucr_hash1_c_7__0_) );
BUFX2 BUFX2_264 ( .A(micro_ucr_hash1_b_8__5_), .Y(micro_ucr_hash1_c_7__1_) );
BUFX2 BUFX2_265 ( .A(micro_ucr_hash1_b_8__6_), .Y(micro_ucr_hash1_c_7__2_) );
BUFX2 BUFX2_266 ( .A(micro_ucr_hash1_b_8__7_), .Y(micro_ucr_hash1_c_7__3_) );
BUFX2 BUFX2_267 ( .A(micro_ucr_hash1_b_9__4_), .Y(micro_ucr_hash1_c_8__0_) );
BUFX2 BUFX2_268 ( .A(micro_ucr_hash1_b_9__5_), .Y(micro_ucr_hash1_c_8__1_) );
BUFX2 BUFX2_269 ( .A(micro_ucr_hash1_b_9__6_), .Y(micro_ucr_hash1_c_8__2_) );
BUFX2 BUFX2_270 ( .A(micro_ucr_hash1_b_9__7_), .Y(micro_ucr_hash1_c_8__3_) );
BUFX2 BUFX2_271 ( .A(micro_ucr_hash1_b_10__4_), .Y(micro_ucr_hash1_c_9__0_) );
BUFX2 BUFX2_272 ( .A(micro_ucr_hash1_b_10__5_), .Y(micro_ucr_hash1_c_9__1_) );
BUFX2 BUFX2_273 ( .A(micro_ucr_hash1_b_10__6_), .Y(micro_ucr_hash1_c_9__2_) );
BUFX2 BUFX2_274 ( .A(micro_ucr_hash1_b_10__7_), .Y(micro_ucr_hash1_c_9__3_) );
endmodule
