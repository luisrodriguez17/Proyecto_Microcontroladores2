`timescale 	1ns	/ 100ps
`include "cmos_cells.v"

module BancoPruebas;

				  



endmodule
