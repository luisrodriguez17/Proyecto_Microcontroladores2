* NGSPICE file created from modulo_rendimiento.ext - technology: scmos

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

.subckt modulo_rendimiento vdd gnd inicio bloque_bytes[0] bloque_bytes[1] bloque_bytes[2]
+ bloque_bytes[3] bloque_bytes[4] bloque_bytes[5] bloque_bytes[6] bloque_bytes[7]
+ bloque_bytes[8] bloque_bytes[9] bloque_bytes[10] bloque_bytes[11] bloque_bytes[12]
+ bloque_bytes[13] bloque_bytes[14] bloque_bytes[15] bloque_bytes[16] bloque_bytes[17]
+ bloque_bytes[18] bloque_bytes[19] bloque_bytes[20] bloque_bytes[21] bloque_bytes[22]
+ bloque_bytes[23] bloque_bytes[24] bloque_bytes[25] bloque_bytes[26] bloque_bytes[27]
+ bloque_bytes[28] bloque_bytes[29] bloque_bytes[30] bloque_bytes[31] bloque_bytes[32]
+ bloque_bytes[33] bloque_bytes[34] bloque_bytes[35] bloque_bytes[36] bloque_bytes[37]
+ bloque_bytes[38] bloque_bytes[39] bloque_bytes[40] bloque_bytes[41] bloque_bytes[42]
+ bloque_bytes[43] bloque_bytes[44] bloque_bytes[45] bloque_bytes[46] bloque_bytes[47]
+ bloque_bytes[48] bloque_bytes[49] bloque_bytes[50] bloque_bytes[51] bloque_bytes[52]
+ bloque_bytes[53] bloque_bytes[54] bloque_bytes[55] bloque_bytes[56] bloque_bytes[57]
+ bloque_bytes[58] bloque_bytes[59] bloque_bytes[60] bloque_bytes[61] bloque_bytes[62]
+ bloque_bytes[63] bloque_bytes[64] bloque_bytes[65] bloque_bytes[66] bloque_bytes[67]
+ bloque_bytes[68] bloque_bytes[69] bloque_bytes[70] bloque_bytes[71] bloque_bytes[72]
+ bloque_bytes[73] bloque_bytes[74] bloque_bytes[75] bloque_bytes[76] bloque_bytes[77]
+ bloque_bytes[78] bloque_bytes[79] bloque_bytes[80] bloque_bytes[81] bloque_bytes[82]
+ bloque_bytes[83] bloque_bytes[84] bloque_bytes[85] bloque_bytes[86] bloque_bytes[87]
+ bloque_bytes[88] bloque_bytes[89] bloque_bytes[90] bloque_bytes[91] bloque_bytes[92]
+ bloque_bytes[93] bloque_bytes[94] bloque_bytes[95] clk reset target[0] target[1]
+ target[2] target[3] target[4] target[5] target[6] target[7] terminado hash[0] hash[1]
+ hash[2] hash[3] hash[4] hash[5] hash[6] hash[7] hash[8] hash[9] hash[10] hash[11]
+ hash[12] hash[13] hash[14] hash[15] hash[16] hash[17] hash[18] hash[19] hash[20]
+ hash[21] hash[22] hash[23]
XNAND2X1_376 NAND2X1_376/A NAND2X1_375/Y gnd NOR2X1_212/B vdd NAND2X1
XNAND3X1_208 INVX1_134/A NAND3X1_208/B OR2X2_91/Y gnd AOI21X1_144/B vdd NAND3X1
XBUFX2_209 BUFX2_209/A gnd BUFX2_209/Y vdd BUFX2
XNOR2X1_62 OR2X2_36/A OR2X2_36/B gnd NOR2X1_62/Y vdd NOR2X1
XOAI21X1_226 INVX2_49/Y AND2X2_78/B INVX1_148/A gnd OAI21X1_227/B vdd OAI21X1
XXNOR2X1_247 AND2X2_191/B AND2X2_192/B gnd XNOR2X1_247/Y vdd XNOR2X1
XNAND2X1_340 NAND2X1_340/A INVX1_202/Y gnd INVX1_203/A vdd NAND2X1
XINVX2_47 INVX2_47/A gnd INVX2_47/Y vdd INVX2
XNOR2X1_259 BUFX2_205/A XOR2X1_213/Y gnd NOR2X1_259/Y vdd NOR2X1
XCLKBUF1_50 BUFX4_7/Y gnd CLKBUF1_50/Y vdd CLKBUF1
XXNOR2X1_211 bloque_bytes[51] bloque_bytes[11] gnd XNOR2X1_211/Y vdd XNOR2X1
XBUFX2_173 BUFX2_173/A gnd BUFX2_173/Y vdd BUFX2
XINVX1_588 INVX1_588/A gnd INVX1_588/Y vdd INVX1
XNAND3X1_172 INVX1_112/A NAND3X1_173/B OR2X2_75/Y gnd AOI21X1_120/B vdd NAND3X1
XNOR2X1_26 INVX1_18/Y NOR2X1_26/B gnd NOR2X1_27/B vdd NOR2X1
XOAI21X1_190 AND2X2_67/Y NOR2X1_124/Y INVX1_125/Y gnd NAND2X1_222/A vdd OAI21X1
XINVX2_11 INVX2_11/A gnd INVX2_11/Y vdd INVX2
XFILL_12_2_1 gnd vdd FILL
XNAND2X1_304 NAND2X1_304/A OAI21X1_262/Y gnd XOR2X1_159/A vdd NAND2X1
XFILL_14_0_0 gnd vdd FILL
XNOR2X1_223 BUFX2_189/A NOR2X1_223/B gnd NOR2X1_223/Y vdd NOR2X1
XCLKBUF1_14 BUFX4_3/Y gnd CLKBUF1_14/Y vdd CLKBUF1
XNAND3X1_136 INVX1_90/A AOI21X1_98/A OR2X2_59/Y gnd AOI21X1_96/B vdd NAND3X1
XINVX1_552 INVX1_552/A gnd INVX1_552/Y vdd INVX1
XBUFX2_137 gnd gnd BUFX2_137/Y vdd BUFX2
XXNOR2X1_175 XNOR2X1_174/Y OAI21X1_409/Y gnd INVX1_319/A vdd XNOR2X1
XOAI21X1_154 XNOR2X1_80/A AOI21X1_113/C AND2X2_54/B gnd XNOR2X1_81/A vdd OAI21X1
XXNOR2X1_97 XNOR2X1_97/A XNOR2X1_97/B gnd BUFX2_161/A vdd XNOR2X1
XNOR2X1_187 BUFX2_177/A NOR2X1_187/B gnd NOR2X1_187/Y vdd NOR2X1
XNAND2X1_268 gnd OR2X2_105/B gnd NAND3X1_239/B vdd NAND2X1
XNOR3X1_67 NOR3X1_67/A NOR3X1_67/B NOR3X1_67/C gnd NOR3X1_67/Y vdd NOR3X1
XFILL_35_9_1 gnd vdd FILL
XBUFX2_101 gnd gnd BUFX2_101/Y vdd BUFX2
XNAND3X1_100 INVX1_68/A AOI21X1_74/A OR2X2_43/Y gnd AOI21X1_72/B vdd NAND3X1
XINVX1_516 INVX1_516/A gnd INVX1_516/Y vdd INVX1
XDFFPOSX1_334 INVX1_386/A CLKBUF1_45/Y OR2X2_148/Y gnd vdd DFFPOSX1
XOAI21X1_118 AND2X2_41/Y NOR2X1_82/Y INVX1_80/Y gnd NAND3X1_123/A vdd OAI21X1
XXNOR2X1_61 XNOR2X1_61/A XNOR2X1_61/B gnd XOR2X1_74/A vdd XNOR2X1
XXNOR2X1_139 gnd XOR2X1_142/Y gnd XNOR2X1_140/A vdd XNOR2X1
XNAND2X1_232 gnd OR2X2_90/B gnd NAND2X1_232/Y vdd NAND2X1
XNOR2X1_151 NOR2X1_151/A INVX2_51/A gnd XOR2X1_140/B vdd NOR2X1
XNOR3X1_31 INVX1_44/Y NOR3X1_31/B NOR3X1_31/C gnd NOR3X1_31/Y vdd NOR3X1
XDFFPOSX1_298 INVX1_301/A CLKBUF1_17/Y AOI21X1_386/C gnd vdd DFFPOSX1
XFILL_11_5_0 gnd vdd FILL
XINVX1_480 INVX1_480/A gnd INVX1_480/Y vdd INVX1
XXNOR2X1_103 gnd XOR2X1_102/Y gnd XNOR2X1_104/A vdd XNOR2X1
XXOR2X1_295 XOR2X1_295/A BUFX2_238/A gnd XOR2X1_295/Y vdd XOR2X1
XXNOR2X1_25 XNOR2X1_25/A OAI21X1_46/B gnd BUFX2_249/A vdd XNOR2X1
XNOR2X1_115 NOR2X1_115/A INVX1_115/Y gnd NOR2X1_115/Y vdd NOR2X1
XNAND2X1_196 INVX1_118/A NAND2X1_196/B gnd OAI21X1_165/A vdd NAND2X1
XAOI21X1_94 AOI21X1_92/Y AOI21X1_94/B AOI21X1_94/C gnd AOI21X1_94/Y vdd AOI21X1
XDFFPOSX1_262 INVX1_215/A CLKBUF1_31/Y INVX1_520/Y gnd vdd DFFPOSX1
XOAI21X1_623 NOR2X1_410/B NOR2X1_410/A OR2X2_142/B gnd AOI21X1_386/A vdd OAI21X1
XFILL_21_0_0 gnd vdd FILL
XOR2X2_83 gnd OR2X2_83/B gnd OR2X2_83/Y vdd OR2X2
XINVX1_444 INVX1_444/A gnd INVX1_444/Y vdd INVX1
XFILL_1_1_0 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XBUFX2_97 gnd gnd BUFX2_97/Y vdd BUFX2
XXOR2X1_259 XOR2X1_259/A BUFX2_222/A gnd XOR2X1_259/Y vdd XOR2X1
XAOI21X1_396 AOI21X1_396/A AOI21X1_396/B NOR3X1_98/Y gnd INVX2_93/A vdd AOI21X1
XNAND2X1_160 OR2X2_60/A OR2X2_60/B gnd AOI21X1_100/A vdd NAND2X1
XDFFPOSX1_226 INVX2_50/A CLKBUF1_18/Y NOR2X1_410/A gnd vdd DFFPOSX1
XAOI21X1_58 AOI21X1_58/A AOI21X1_58/B NAND2X1_94/Y gnd OAI21X1_74/A vdd AOI21X1
XOR2X2_47 OR2X2_47/A INVX1_72/Y gnd OR2X2_47/Y vdd OR2X2
XOAI21X1_587 NAND3X1_501/Y INVX2_80/Y BUFX4_30/Y gnd AOI21X1_347/C vdd OAI21X1
XINVX1_408 INVX1_408/A gnd INVX1_408/Y vdd INVX1
XNAND2X1_701 NOR2X1_444/B OAI21X1_633/Y gnd NAND2X1_701/Y vdd NAND2X1
XXOR2X1_223 XOR2X1_223/A BUFX2_206/A gnd XOR2X1_223/Y vdd XOR2X1
XBUFX2_61 gnd gnd BUFX2_61/Y vdd BUFX2
XNAND3X1_533 NAND3X1_533/A NAND3X1_533/B NAND2X1_704/Y gnd XNOR2X1_254/B vdd NAND3X1
XNAND2X1_124 AND2X2_36/B AND2X2_36/A gnd AOI21X1_77/C vdd NAND2X1
XAOI21X1_360 bloque_bytes[78] INVX2_87/Y INVX1_548/A gnd OAI21X1_599/C vdd AOI21X1
XAOI21X1_22 AOI21X1_22/A AOI21X1_22/B OAI21X1_21/B gnd OAI21X1_23/A vdd AOI21X1
XFILL_9_1 gnd vdd FILL
XDFFPOSX1_190 INVX1_102/A CLKBUF1_49/Y bloque_bytes[20] gnd vdd DFFPOSX1
XDFFPOSX1_2 BUFX2_1/A CLKBUF1_4/Y NOR3X1_1/Y gnd vdd DFFPOSX1
XOR2X2_11 gnd OR2X2_11/B gnd OR2X2_11/Y vdd OR2X2
XXOR2X1_187 XOR2X1_187/A BUFX2_186/A gnd XOR2X1_187/Y vdd XOR2X1
XINVX1_372 INVX1_372/A gnd INVX1_372/Y vdd INVX1
XOAI21X1_551 NOR3X1_86/A NOR3X1_86/C INVX2_73/A gnd NOR2X1_349/A vdd OAI21X1
XNAND2X1_665 bloque_bytes[2] OR2X2_139/A gnd AOI21X1_381/A vdd NAND2X1
XBUFX2_25 BUFX4_8/Y gnd terminado vdd BUFX2
XOAI21X1_70 AND2X2_25/Y NOR2X1_54/Y INVX1_48/A gnd NAND3X1_71/B vdd OAI21X1
XNAND2X1_85 INVX2_21/Y NAND3X1_74/C gnd OAI21X1_69/A vdd NAND2X1
XNAND3X1_497 inicio INVX1_486/Y AND2X2_174/Y gnd NOR3X1_91/C vdd NAND3X1
XDFFPOSX1_88 INVX2_81/A CLKBUF1_6/Y AOI21X1_348/Y gnd vdd DFFPOSX1
XAOI21X1_324 INVX2_74/Y NAND2X1_611/Y OAI21X1_568/Y gnd AOI21X1_324/Y vdd AOI21X1
XFILL_16_7_1 gnd vdd FILL
XFILL_18_5_0 gnd vdd FILL
XDFFPOSX1_154 INVX2_23/A CLKBUF1_44/Y bloque_bytes[48] gnd vdd DFFPOSX1
XINVX1_336 INVX1_336/A gnd INVX1_336/Y vdd INVX1
XOAI21X1_515 gnd NOR2X1_327/B INVX1_419/A gnd INVX1_421/A vdd OAI21X1
XNAND2X1_629 NOR2X1_403/Y AND2X2_172/B gnd INVX2_84/A vdd NAND2X1
XXOR2X1_151 BUFX2_170/A XOR2X1_151/B gnd XOR2X1_151/Y vdd XOR2X1
XBUFX2_3 BUFX2_3/A gnd hash[2] vdd BUFX2
XFILL_26_2_1 gnd vdd FILL
XAOI21X1_288 AOI21X1_288/A AOI21X1_288/B AOI21X1_288/C gnd OAI21X1_486/A vdd AOI21X1
XFILL_28_0_0 gnd vdd FILL
XNAND2X1_49 XOR2X1_3/A OR2X2_13/B gnd NAND3X1_34/B vdd NAND2X1
XOAI21X1_34 OAI21X1_29/A XNOR2X1_16/B OAI21X1_34/C gnd OAI21X1_34/Y vdd OAI21X1
XDFFPOSX1_118 INVX1_593/A CLKBUF1_25/Y bloque_bytes[92] gnd vdd DFFPOSX1
XFILL_6_3_1 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XDFFPOSX1_52 INVX1_544/A CLKBUF1_36/Y AND2X2_167/Y gnd vdd DFFPOSX1
XNAND3X1_461 INVX1_430/Y INVX1_433/Y AND2X2_149/A gnd NAND3X1_461/Y vdd NAND3X1
XXOR2X1_95 XOR2X1_90/Y gnd gnd OR2X2_83/B vdd XOR2X1
XXOR2X1_115 BUFX2_162/A gnd gnd OR2X2_99/B vdd XOR2X1
XINVX1_300 INVX1_300/A gnd INVX1_300/Y vdd INVX1
XOAI21X1_479 BUFX2_219/A INVX1_385/A INVX1_386/Y gnd OAI21X1_479/Y vdd OAI21X1
XNAND2X1_593 INVX1_455/Y NOR2X1_348/Y gnd NAND3X1_476/B vdd NAND2X1
XNAND2X1_13 INVX1_7/A INVX4_1/Y gnd NAND3X1_3/A vdd NAND2X1
XNAND3X1_425 INVX1_382/A NAND3X1_425/B NAND3X1_425/C gnd AOI21X1_287/A vdd NAND3X1
XAOI21X1_252 OAI21X1_403/Y AOI21X1_252/B INVX1_307/A gnd NOR2X1_256/A vdd AOI21X1
XINVX1_264 INVX1_264/A gnd INVX1_264/Y vdd INVX1
XDFFPOSX1_16 BUFX2_15/A CLKBUF1_28/Y NOR3X1_15/Y gnd vdd DFFPOSX1
XNAND3X1_90 INVX1_59/A NAND3X1_88/B OR2X2_37/Y gnd OR2X2_40/B vdd NAND3X1
XAND2X2_195 vdd gnd gnd AND2X2_195/Y vdd AND2X2
XXOR2X1_59 XOR2X1_59/A XOR2X1_61/A gnd XOR2X1_59/Y vdd XOR2X1
XOAI21X1_443 NOR2X1_281/Y NOR2X1_280/B AOI22X1_16/C gnd XOR2X1_242/A vdd OAI21X1
XNAND2X1_557 INVX1_419/A NOR2X1_327/Y gnd NAND3X1_451/C vdd NAND2X1
XOR2X2_142 OR2X2_142/A OR2X2_142/B gnd OR2X2_142/Y vdd OR2X2
XAOI21X1_216 AOI21X1_216/A AOI21X1_216/B NAND2X1_355/Y gnd OAI21X1_315/A vdd AOI21X1
XNAND3X1_389 INVX1_329/A INVX1_327/Y INVX1_328/Y gnd NAND3X1_389/Y vdd NAND3X1
XAND2X2_159 BUFX4_33/Y AND2X2_159/B gnd AND2X2_159/Y vdd AND2X2
XINVX1_228 NOR3X1_61/B gnd INVX1_228/Y vdd INVX1
XFILL_25_5_0 gnd vdd FILL
XOAI21X1_407 BUFX2_204/A XOR2X1_212/Y INVX1_311/A gnd AOI22X1_14/B vdd OAI21X1
XNAND3X1_54 INVX1_37/A NAND3X1_52/B OR2X2_21/Y gnd OR2X2_24/B vdd NAND3X1
XXOR2X1_23 OR2X2_29/A gnd gnd OR2X2_25/B vdd XOR2X1
XFILL_5_6_0 gnd vdd FILL
XFILL_23_7_1 gnd vdd FILL
XOR2X2_106 gnd AND2X2_81/B gnd OR2X2_106/Y vdd OR2X2
XNAND2X1_521 AOI21X1_287/A INVX1_389/A gnd NAND2X1_521/Y vdd NAND2X1
XNOR2X1_440 NOR2X1_439/Y NOR2X1_440/B gnd NOR2X1_440/Y vdd NOR2X1
XFILL_3_8_1 gnd vdd FILL
XAOI21X1_180 AOI21X1_180/A AOI21X1_180/B AOI21X1_180/C gnd NOR2X1_161/A vdd AOI21X1
XNAND3X1_353 AOI22X1_12/B INVX1_276/A INVX1_274/Y gnd NAND2X1_410/B vdd NAND3X1
XNAND2X1_2 NAND2X1_2/A NAND2X1_2/B gnd NOR2X1_2/A vdd NAND2X1
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XFILL_35_0_0 gnd vdd FILL
XOAI22X1_1 INVX4_1/Y INVX2_1/A INVX2_3/Y INVX2_2/A gnd NOR2X1_8/A vdd OAI22X1
XNAND3X1_18 INVX1_15/A NAND3X1_16/B OR2X2_5/Y gnd OR2X2_8/B vdd NAND3X1
XINVX1_192 INVX1_192/A gnd INVX1_192/Y vdd INVX1
XNOR2X1_404 INVX2_78/Y INVX2_79/Y gnd NOR2X1_404/Y vdd NOR2X1
XOAI21X1_371 BUFX2_193/A XOR2X1_195/Y INVX1_277/A gnd OAI21X1_371/Y vdd OAI21X1
XAND2X2_123 AND2X2_123/A INVX1_302/Y gnd NOR3X1_70/C vdd AND2X2
XFILL_33_2_1 gnd vdd FILL
XNAND2X1_485 INVX1_349/Y NOR2X1_282/Y gnd INVX1_352/A vdd NAND2X1
XNAND3X1_317 INVX1_223/Y INVX1_222/A AOI21X1_218/B gnd AND2X2_105/B vdd NAND3X1
XAND2X2_96 AND2X2_96/A AND2X2_96/B gnd AND2X2_96/Y vdd AND2X2
XAOI21X1_144 AOI21X1_144/A AOI21X1_144/B NAND3X1_206/C gnd NOR2X1_131/A vdd AOI21X1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XOAI21X1_335 NOR2X1_209/A NOR3X1_61/Y OAI21X1_335/C gnd AOI21X1_226/B vdd OAI21X1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XNOR2X1_368 BUFX4_16/Y INVX1_479/Y gnd NOR2X1_368/Y vdd NOR2X1
XNAND2X1_449 INVX1_303/A NOR2X1_252/Y gnd NAND2X1_449/Y vdd NAND2X1
XAOI21X1_108 NAND3X1_157/A NAND3X1_154/Y AOI21X1_108/C gnd NOR2X1_101/A vdd AOI21X1
XAND2X2_60 AND2X2_60/A AND2X2_60/B gnd AND2X2_60/Y vdd AND2X2
XNAND3X1_281 INVX1_178/Y NAND3X1_281/B OR2X2_123/Y gnd AOI21X1_193/B vdd NAND3X1
XOAI21X1_299 gnd XOR2X1_162/Y INVX1_206/A gnd NAND2X1_344/A vdd OAI21X1
XINVX1_120 INVX1_120/A gnd INVX1_120/Y vdd INVX1
XNOR2X1_332 INVX1_428/Y NOR2X1_332/B gnd INVX1_430/A vdd NOR2X1
XNAND2X1_413 INVX1_277/Y NOR2X1_235/Y gnd NAND2X1_414/B vdd NAND2X1
XAND2X2_24 AND2X2_24/A AND2X2_24/B gnd AND2X2_24/Y vdd AND2X2
XNAND3X1_245 INVX1_156/Y NAND3X1_245/B OR2X2_107/Y gnd AOI21X1_169/B vdd NAND3X1
XFILL_32_5_0 gnd vdd FILL
XFILL_30_7_1 gnd vdd FILL
XBUFX2_246 BUFX2_246/A gnd BUFX2_246/Y vdd BUFX2
XNOR2X1_99 gnd OR2X2_66/B gnd NOR3X1_42/B vdd NOR2X1
XINVX2_84 INVX2_84/A gnd INVX2_84/Y vdd INVX2
XOAI21X1_263 NOR3X1_55/C NOR3X1_55/B NOR3X1_55/A gnd OAI21X1_263/Y vdd OAI21X1
XNOR2X1_296 INVX1_371/Y NOR2X1_296/B gnd INVX1_373/A vdd NOR2X1
XNAND2X1_377 INVX1_238/Y NOR2X1_212/B gnd NAND2X1_378/A vdd NAND2X1
XNAND3X1_209 INVX1_134/Y NAND3X1_208/B OR2X2_91/Y gnd AOI21X1_145/B vdd NAND3X1
XBUFX2_210 BUFX2_210/A gnd BUFX2_210/Y vdd BUFX2
XNOR2X1_63 NOR2X1_63/A NOR2X1_63/B gnd NOR2X1_63/Y vdd NOR2X1
XOAI21X1_227 OAI21X1_227/A OAI21X1_227/B INVX1_150/Y gnd NAND3X1_238/C vdd OAI21X1
XXNOR2X1_248 NOR2X1_442/B INVX1_583/A gnd XNOR2X1_248/Y vdd XNOR2X1
XNAND2X1_341 NAND2X1_341/A AOI22X1_8/C gnd AOI21X1_209/C vdd NAND2X1
XINVX2_48 INVX2_48/A gnd INVX2_48/Y vdd INVX2
XNOR2X1_260 INVX1_314/Y NOR2X1_260/B gnd INVX1_316/A vdd NOR2X1
XNOR2X1_27 NOR2X1_27/A NOR2X1_27/B gnd XOR2X1_18/A vdd NOR2X1
XBUFX2_174 BUFX2_174/A gnd BUFX2_174/Y vdd BUFX2
XXNOR2X1_212 bloque_bytes[52] bloque_bytes[12] gnd NAND2X1_654/A vdd XNOR2X1
XCLKBUF1_51 BUFX4_4/Y gnd CLKBUF1_51/Y vdd CLKBUF1
XINVX1_589 INVX1_589/A gnd INVX1_589/Y vdd INVX1
XNAND3X1_173 INVX1_112/Y NAND3X1_173/B OR2X2_75/Y gnd AOI21X1_121/B vdd NAND3X1
XINVX2_12 INVX2_12/A gnd INVX2_12/Y vdd INVX2
XFILL_14_0_1 gnd vdd FILL
XOAI21X1_191 XNOR2X1_98/A AOI21X1_142/C NOR2X1_125/Y gnd NOR2X1_126/B vdd OAI21X1
XNOR2X1_224 INVX1_257/Y NOR2X1_224/B gnd INVX1_259/A vdd NOR2X1
XNAND2X1_305 INVX2_56/Y XNOR2X1_140/A gnd NAND3X1_276/C vdd NAND2X1
XCLKBUF1_15 BUFX4_7/Y gnd CLKBUF1_15/Y vdd CLKBUF1
XBUFX2_138 gnd gnd BUFX2_138/Y vdd BUFX2
XINVX1_553 INVX1_553/A gnd INVX1_553/Y vdd INVX1
XNAND3X1_137 INVX1_90/Y AOI21X1_98/A OR2X2_59/Y gnd AOI21X1_97/B vdd NAND3X1
XXNOR2X1_98 XNOR2X1_98/A AND2X2_66/Y gnd XNOR2X1_98/Y vdd XNOR2X1
XOAI21X1_155 AND2X2_55/Y NOR2X1_104/Y INVX1_103/A gnd OAI21X1_155/Y vdd OAI21X1
XXNOR2X1_176 NOR2X1_266/A NAND2X1_464/Y gnd BUFX2_218/A vdd XNOR2X1
XNOR2X1_188 INVX1_200/Y NOR2X1_188/B gnd INVX1_202/A vdd NOR2X1
XNAND2X1_269 NAND2X1_269/A NAND2X1_269/B gnd XNOR2X1_123/A vdd NAND2X1
XDFFPOSX1_335 INVX1_387/A CLKBUF1_19/Y NAND2X1_681/Y gnd vdd DFFPOSX1
XNOR3X1_68 NOR3X1_68/A INVX2_64/Y NOR3X1_68/C gnd NOR3X1_68/Y vdd NOR3X1
XNAND3X1_101 INVX1_68/Y AOI21X1_74/A OR2X2_43/Y gnd AOI21X1_73/B vdd NAND3X1
XINVX1_517 INVX1_517/A gnd INVX1_517/Y vdd INVX1
XBUFX2_102 gnd gnd BUFX2_102/Y vdd BUFX2
XOAI21X1_119 OAI21X1_119/A XNOR2X1_61/B AOI21X1_87/Y gnd NAND3X1_128/C vdd OAI21X1
XXNOR2X1_62 XNOR2X1_62/A AND2X2_42/Y gnd XOR2X1_76/A vdd XNOR2X1
XXNOR2X1_140 XNOR2X1_140/A INVX2_56/Y gnd BUFX2_179/A vdd XNOR2X1
XNAND2X1_233 NAND2X1_233/A NAND2X1_233/B gnd XNOR2X1_106/A vdd NAND2X1
XNOR2X1_152 OR2X2_108/A OR2X2_108/B gnd NOR2X1_152/Y vdd NOR2X1
XNOR3X1_32 INVX1_45/Y NOR2X1_49/Y AND2X2_21/Y gnd NOR2X1_53/B vdd NOR3X1
XINVX1_481 INVX1_481/A gnd INVX1_481/Y vdd INVX1
XFILL_13_3_0 gnd vdd FILL
XDFFPOSX1_299 INVX1_302/A CLKBUF1_34/Y AOI21X1_387/C gnd vdd DFFPOSX1
XFILL_11_5_1 gnd vdd FILL
XXNOR2X1_104 XNOR2X1_104/A INVX2_44/Y gnd OR2X2_108/A vdd XNOR2X1
XXOR2X1_296 XOR2X1_296/A XOR2X1_296/B gnd XOR2X1_296/Y vdd XOR2X1
XXNOR2X1_26 OAI21X1_55/A AND2X2_18/Y gnd XOR2X1_36/A vdd XNOR2X1
XNOR2X1_116 INVX1_117/Y NOR2X1_116/B gnd NOR2X1_117/B vdd NOR2X1
XNAND2X1_197 gnd OR2X2_75/B gnd NAND3X1_173/B vdd NAND2X1
XDFFPOSX1_263 INVX1_216/A CLKBUF1_11/Y INVX1_523/Y gnd vdd DFFPOSX1
XOR2X2_84 OR2X2_84/A OR2X2_84/B gnd OR2X2_84/Y vdd OR2X2
XOAI21X1_624 NOR2X1_411/B NOR2X1_411/A OR2X2_143/B gnd OAI21X1_624/Y vdd OAI21X1
XFILL_21_0_1 gnd vdd FILL
XAOI21X1_95 AOI21X1_95/A OR2X2_58/Y INVX1_89/A gnd NOR2X1_93/A vdd AOI21X1
XINVX1_445 INVX1_445/A gnd INVX1_445/Y vdd INVX1
XFILL_1_1_1 gnd vdd FILL
XBUFX2_98 gnd gnd BUFX2_98/Y vdd BUFX2
XXOR2X1_260 XOR2X1_260/A XOR2X1_260/B gnd XOR2X1_266/A vdd XOR2X1
XAOI21X1_397 NAND3X1_537/B OR2X2_157/Y INVX1_592/A gnd NAND3X1_542/C vdd AOI21X1
XNAND2X1_161 INVX2_33/Y NAND3X1_146/C gnd XNOR2X1_71/A vdd NAND2X1
XAOI21X1_59 NAND2X1_99/Y OR2X2_34/Y INVX1_56/A gnd NOR2X1_63/A vdd AOI21X1
XDFFPOSX1_227 INVX1_154/A CLKBUF1_40/Y NOR2X1_411/A gnd vdd DFFPOSX1
XOR2X2_48 OR2X2_48/A OR2X2_48/B gnd OR2X2_48/Y vdd OR2X2
XOAI21X1_588 NAND3X1_501/Y NAND2X1_636/Y BUFX4_30/Y gnd OAI21X1_588/Y vdd OAI21X1
XINVX1_409 INVX1_409/A gnd INVX1_409/Y vdd INVX1
XXOR2X1_224 XOR2X1_224/A XOR2X1_224/B gnd XOR2X1_230/A vdd XOR2X1
XNAND2X1_702 INVX1_589/Y NOR2X1_444/Y gnd NAND2X1_703/B vdd NAND2X1
XBUFX2_62 gnd gnd BUFX2_62/Y vdd BUFX2
XNAND3X1_534 INVX1_591/A AOI21X1_394/A OR2X2_156/Y gnd NAND3X1_535/C vdd NAND3X1
XNAND2X1_125 OR2X2_45/A OR2X2_45/B gnd NAND3X1_106/B vdd NAND2X1
XFILL_9_2 gnd vdd FILL
XFILL_10_8_0 gnd vdd FILL
XAOI21X1_361 bloque_bytes[79] INVX1_505/Y OR2X2_149/B gnd AND2X2_177/A vdd AOI21X1
XOR2X2_12 XOR2X1_2/A OR2X2_12/B gnd OR2X2_12/Y vdd OR2X2
XAOI21X1_23 NAND3X1_25/B OR2X2_10/Y INVX1_23/A gnd NOR2X1_33/A vdd AOI21X1
XDFFPOSX1_191 INVX1_103/A CLKBUF1_16/Y bloque_bytes[21] gnd vdd DFFPOSX1
XOAI21X1_552 gnd XOR2X1_282/Y INVX1_457/Y gnd OAI21X1_552/Y vdd OAI21X1
XDFFPOSX1_3 BUFX2_2/A CLKBUF1_4/Y NOR3X1_2/Y gnd vdd DFFPOSX1
XINVX1_373 INVX1_373/A gnd INVX1_373/Y vdd INVX1
XXOR2X1_188 XOR2X1_188/A XOR2X1_188/B gnd XOR2X1_188/Y vdd XOR2X1
XNAND2X1_666 bloque_bytes[3] OR2X2_152/B gnd AOI21X1_382/B vdd NAND2X1
XAOI21X1_325 INVX1_474/A INVX4_2/Y OAI21X1_570/Y gnd DFFPOSX1_63/D vdd AOI21X1
XFILL_18_5_1 gnd vdd FILL
XFILL_20_3_0 gnd vdd FILL
XBUFX2_26 BUFX2_26/A gnd BUFX2_26/Y vdd BUFX2
XFILL_0_4_0 gnd vdd FILL
XOAI21X1_71 AND2X2_25/Y NOR2X1_54/Y INVX1_48/Y gnd NAND3X1_73/A vdd OAI21X1
XNAND2X1_86 AND2X2_24/B AND2X2_24/A gnd OAI21X1_69/B vdd NAND2X1
XDFFPOSX1_89 INVX1_485/A CLKBUF1_16/Y NOR3X1_96/Y gnd vdd DFFPOSX1
XDFFPOSX1_155 INVX1_55/A CLKBUF1_33/Y bloque_bytes[49] gnd vdd DFFPOSX1
XNAND3X1_498 INVX1_491/Y NOR3X1_91/Y INVX2_84/Y gnd NOR3X1_95/C vdd NAND3X1
XINVX1_337 INVX1_337/A gnd INVX1_337/Y vdd INVX1
XOAI21X1_516 INVX1_422/A INVX1_423/A INVX1_424/A gnd INVX1_426/A vdd OAI21X1
XNAND2X1_630 INVX2_84/Y INVX2_83/A gnd OAI21X1_583/A vdd NAND2X1
XXOR2X1_152 INVX1_194/A gnd gnd NOR2X1_178/B vdd XOR2X1
XBUFX2_4 BUFX2_4/A gnd hash[3] vdd BUFX2
XNAND2X1_50 AOI21X1_29/A AOI21X1_29/B gnd INVX2_16/A vdd NAND2X1
XNAND3X1_462 INVX2_72/A NAND3X1_462/B NAND2X1_573/Y gnd NOR3X1_83/A vdd NAND3X1
XAOI21X1_289 NAND2X1_524/A NAND2X1_524/B AOI21X1_289/C gnd AOI21X1_289/Y vdd AOI21X1
XFILL_28_0_1 gnd vdd FILL
XOAI21X1_35 OAI21X1_35/A OAI21X1_35/B AND2X2_12/B gnd OAI21X1_35/Y vdd OAI21X1
XDFFPOSX1_119 INVX1_594/A CLKBUF1_25/Y bloque_bytes[93] gnd vdd DFFPOSX1
XFILL_8_1_1 gnd vdd FILL
XDFFPOSX1_53 INVX1_571/A CLKBUF1_14/Y NOR2X1_375/Y gnd vdd DFFPOSX1
XXOR2X1_116 XNOR2X1_98/Y OR2X2_92/A gnd AND2X2_77/B vdd XOR2X1
XXOR2X1_96 XOR2X1_96/A OR2X2_76/A gnd OR2X2_84/B vdd XOR2X1
XOAI21X1_480 NOR3X1_77/C OAI21X1_474/C INVX1_389/A gnd NOR2X1_305/A vdd OAI21X1
XINVX1_301 INVX1_301/A gnd INVX1_301/Y vdd INVX1
XNAND2X1_594 INVX1_458/A NAND3X1_476/B gnd INVX1_456/A vdd NAND2X1
XDFFPOSX1_17 BUFX2_16/A CLKBUF1_48/Y NOR3X1_16/Y gnd vdd DFFPOSX1
XNAND2X1_14 INVX1_8/A INVX2_3/Y gnd NAND3X1_3/B vdd NAND2X1
XNAND3X1_426 INVX1_383/A AOI21X1_285/B INVX1_382/Y gnd INVX1_389/A vdd NAND3X1
XAOI21X1_253 INVX1_307/A AOI21X1_253/B INVX1_306/Y gnd NOR3X1_69/C vdd AOI21X1
XAND2X2_196 gnd gnd gnd AND2X2_196/Y vdd AND2X2
XFILL_17_8_0 gnd vdd FILL
XINVX1_265 INVX1_265/A gnd INVX1_265/Y vdd INVX1
XOAI21X1_444 BUFX2_212/A XOR2X1_230/Y INVX1_349/Y gnd OAI21X1_444/Y vdd OAI21X1
XNAND3X1_91 NAND3X1_91/A OR2X2_40/B OR2X2_38/B gnd AOI21X1_65/B vdd NAND3X1
XXOR2X1_60 XOR2X1_60/A NOR2X1_71/Y gnd BUFX2_262/A vdd XOR2X1
XOR2X2_143 OR2X2_143/A OR2X2_143/B gnd OR2X2_143/Y vdd OR2X2
XNAND2X1_558 INVX1_419/Y NOR2X1_327/Y gnd NAND3X1_452/B vdd NAND2X1
XAOI21X1_217 AOI21X1_217/A AOI21X1_217/B NAND2X1_360/Y gnd OAI21X1_316/C vdd AOI21X1
XFILL_27_3_0 gnd vdd FILL
XNAND3X1_390 INVX1_331/A NAND3X1_388/Y INVX1_326/Y gnd AOI22X1_15/C vdd NAND3X1
XXOR2X1_24 BUFX2_241/A gnd gnd OR2X2_26/B vdd XOR2X1
XFILL_7_4_0 gnd vdd FILL
XAND2X2_160 INVX8_2/A AND2X2_169/B gnd AND2X2_160/Y vdd AND2X2
XINVX1_229 INVX1_229/A gnd INVX1_229/Y vdd INVX1
XFILL_25_5_1 gnd vdd FILL
XOAI21X1_408 gnd NOR2X1_252/B INVX1_303/Y gnd OAI21X1_408/Y vdd OAI21X1
XNOR2X1_441 INVX2_91/Y INVX1_581/Y gnd NOR2X1_441/Y vdd NOR2X1
XNAND3X1_55 NAND3X1_55/A OR2X2_24/B OR2X2_22/B gnd AOI21X1_41/B vdd NAND3X1
XFILL_5_6_1 gnd vdd FILL
XOR2X2_107 gnd AND2X2_82/B gnd OR2X2_107/Y vdd OR2X2
XNAND2X1_522 INVX1_387/A NOR2X1_306/Y gnd NAND3X1_430/C vdd NAND2X1
XAOI21X1_181 OAI21X1_252/Y NAND3X1_263/Y NOR3X1_54/Y gnd INVX2_54/A vdd AOI21X1
XNAND3X1_354 INVX1_266/Y NAND3X1_347/Y NOR3X1_66/Y gnd AOI21X1_240/B vdd NAND3X1
XNAND2X1_3 NAND2X1_3/A NAND2X1_3/B gnd OAI21X1_2/A vdd NAND2X1
XINVX1_75 OR2X2_48/Y gnd INVX1_75/Y vdd INVX1
XINVX1_193 INVX1_193/A gnd INVX1_193/Y vdd INVX1
XOAI22X1_2 INVX2_1/Y target[5] target[4] INVX2_2/Y gnd NOR2X1_8/B vdd OAI22X1
XFILL_35_0_1 gnd vdd FILL
XNAND3X1_19 NAND3X1_19/A OR2X2_8/B OR2X2_6/B gnd AOI21X1_17/B vdd NAND3X1
XNOR2X1_405 NOR2X1_405/A NOR2X1_405/B gnd NOR2X1_405/Y vdd NOR2X1
XOAI21X1_372 OAI21X1_372/A INVX1_280/A INVX1_279/Y gnd AND2X2_117/A vdd OAI21X1
XAND2X2_124 AND2X2_124/A NOR3X1_69/A gnd BUFX2_212/A vdd AND2X2
XNAND2X1_486 NAND2X1_486/A NAND2X1_486/B gnd XOR2X1_242/B vdd NAND2X1
XAOI21X1_145 AOI21X1_145/A AOI21X1_145/B NOR3X1_48/Y gnd INVX2_45/A vdd AOI21X1
XINVX1_39 INVX1_39/A gnd OR2X2_23/B vdd INVX1
XNAND3X1_318 INVX1_221/Y INVX1_224/Y AND2X2_105/A gnd NAND2X1_361/B vdd NAND3X1
XAND2X2_97 OR2X2_125/A OR2X2_125/B gnd AND2X2_97/Y vdd AND2X2
XOAI21X1_336 OAI21X1_336/A INVX1_240/A INVX1_243/A gnd NAND2X1_380/A vdd OAI21X1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XNOR2X1_369 BUFX4_16/Y INVX1_480/Y gnd NOR2X1_369/Y vdd NOR2X1
XNAND2X1_450 XOR2X1_224/B NOR2X1_256/Y gnd NAND2X1_450/Y vdd NAND2X1
XAOI21X1_109 AOI21X1_109/A AOI21X1_109/B NOR3X1_42/Y gnd INVX2_36/A vdd AOI21X1
XNAND3X1_282 INVX1_179/Y AOI21X1_196/A OR2X2_124/Y gnd NAND3X1_283/B vdd NAND3X1
XFILL_24_8_0 gnd vdd FILL
XAND2X2_61 OR2X2_77/A OR2X2_77/B gnd AND2X2_61/Y vdd AND2X2
XFILL_4_9_0 gnd vdd FILL
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XOAI21X1_300 gnd NOR2X1_191/B INVX1_207/A gnd INVX2_60/A vdd OAI21X1
XNOR2X1_333 BUFX2_230/A NOR2X1_333/B gnd NOR2X1_333/Y vdd NOR2X1
XNAND2X1_414 OAI21X1_371/Y NAND2X1_414/B gnd NOR2X1_236/B vdd NAND2X1
XFILL_34_3_0 gnd vdd FILL
XAND2X2_25 OR2X2_29/A OR2X2_29/B gnd AND2X2_25/Y vdd AND2X2
XBUFX2_247 OR2X2_36/A gnd BUFX2_247/Y vdd BUFX2
XNAND3X1_246 INVX1_157/Y NAND3X1_248/B OR2X2_108/Y gnd NAND3X1_247/B vdd NAND3X1
XFILL_32_5_1 gnd vdd FILL
XOAI21X1_264 NOR3X1_56/Y NOR2X1_173/A NOR3X1_55/Y gnd NAND2X1_309/B vdd OAI21X1
XBUFX4_10 BUFX4_8/A gnd MUX2X1_9/S vdd BUFX4
XNAND2X1_378 NAND2X1_378/A INVX1_240/Y gnd INVX1_241/A vdd NAND2X1
XINVX2_85 bloque_bytes[34] gnd INVX2_85/Y vdd INVX2
XNOR2X1_297 BUFX2_218/A XOR2X1_241/Y gnd NOR2X1_297/Y vdd NOR2X1
XNOR2X1_64 OR2X2_37/A OR2X2_37/B gnd NOR2X1_64/Y vdd NOR2X1
XNAND3X1_210 INVX1_135/Y AOI21X1_148/A OR2X2_92/Y gnd NAND3X1_211/B vdd NAND3X1
XBUFX2_211 INVX1_346/A gnd BUFX2_211/Y vdd BUFX2
XXNOR2X1_249 NOR2X1_444/B XOR2X1_296/Y gnd XNOR2X1_249/Y vdd XNOR2X1
XOAI21X1_228 NOR2X1_147/A INVX1_152/Y INVX1_153/Y gnd NAND2X1_266/B vdd OAI21X1
XNAND2X1_342 OAI21X1_298/Y NAND2X1_342/B gnd XOR2X1_178/A vdd NAND2X1
XINVX2_49 INVX2_49/A gnd INVX2_49/Y vdd INVX2
XNOR2X1_261 BUFX2_206/A XOR2X1_214/Y gnd NOR2X1_261/Y vdd NOR2X1
XINVX1_590 INVX1_590/A gnd INVX1_590/Y vdd INVX1
XNAND3X1_174 INVX1_113/Y NAND3X1_176/B OR2X2_76/Y gnd NAND3X1_174/Y vdd NAND3X1
XNOR2X1_28 gnd OR2X2_9/B gnd NOR2X1_28/Y vdd NOR2X1
XXNOR2X1_213 bloque_bytes[55] bloque_bytes[15] gnd XNOR2X1_213/Y vdd XNOR2X1
XBUFX2_175 INVX1_194/A gnd BUFX2_175/Y vdd BUFX2
XFILL_31_8_0 gnd vdd FILL
XINVX2_13 INVX2_13/A gnd INVX2_13/Y vdd INVX2
XNOR2X1_225 BUFX2_190/A XOR2X1_187/Y gnd NOR2X1_225/Y vdd NOR2X1
XOAI21X1_192 INVX2_43/Y AND2X2_66/B OR2X2_86/Y gnd OAI21X1_193/B vdd OAI21X1
XNAND2X1_306 gnd AND2X2_92/B gnd NAND2X1_306/Y vdd NAND2X1
XCLKBUF1_16 BUFX4_7/Y gnd CLKBUF1_16/Y vdd CLKBUF1
XNAND3X1_138 INVX1_91/Y AOI21X1_100/A OR2X2_60/Y gnd NAND3X1_138/Y vdd NAND3X1
XBUFX2_139 gnd gnd BUFX2_139/Y vdd BUFX2
XINVX1_554 INVX1_554/A gnd INVX1_554/Y vdd INVX1
XOAI21X1_156 AND2X2_55/Y NOR2X1_104/Y INVX1_103/Y gnd OAI21X1_156/Y vdd OAI21X1
XXNOR2X1_99 XNOR2X1_99/A INVX2_43/Y gnd XOR2X1_117/A vdd XNOR2X1
XXNOR2X1_177 NOR2X1_269/Y NOR2X1_268/Y gnd XOR2X1_238/A vdd XNOR2X1
XNOR2X1_189 BUFX2_178/A NOR2X1_189/B gnd NOR2X1_189/Y vdd NOR2X1
XNAND2X1_270 gnd AND2X2_81/B gnd AOI21X1_167/A vdd NAND2X1
XDFFPOSX1_336 INVX1_391/A CLKBUF1_19/Y NAND2X1_682/Y gnd vdd DFFPOSX1
XNOR3X1_69 NOR3X1_69/A NOR3X1_69/B NOR3X1_69/C gnd NOR3X1_69/Y vdd NOR3X1
XINVX1_518 bloque_bytes[60] gnd INVX1_518/Y vdd INVX1
XNAND3X1_102 INVX1_69/Y AOI21X1_76/A OR2X2_44/Y gnd NAND3X1_102/Y vdd NAND3X1
XXNOR2X1_141 XNOR2X1_141/A NAND3X1_276/C gnd BUFX2_180/A vdd XNOR2X1
XBUFX2_103 gnd gnd BUFX2_103/Y vdd BUFX2
XOAI21X1_120 XNOR2X1_62/A AOI21X1_89/C AND2X2_42/B gnd XNOR2X1_63/A vdd OAI21X1
XXNOR2X1_63 XNOR2X1_63/A INVX2_31/Y gnd XOR2X1_77/A vdd XNOR2X1
XNOR2X1_153 NOR2X1_153/A NOR3X1_52/Y gnd NOR2X1_153/Y vdd NOR2X1
XNOR3X1_33 INVX1_55/Y NOR2X1_58/Y AND2X2_26/Y gnd NOR3X1_33/Y vdd NOR3X1
XFILL_15_1_0 gnd vdd FILL
XNAND2X1_234 INVX1_140/A OAI21X1_198/Y gnd OAI21X1_199/A vdd NAND2X1
XINVX1_482 INVX1_482/A gnd INVX1_482/Y vdd INVX1
XFILL_13_3_1 gnd vdd FILL
XDFFPOSX1_300 INVX1_303/A CLKBUF1_34/Y AOI21X1_388/C gnd vdd DFFPOSX1
XXNOR2X1_27 OAI21X1_52/Y INVX2_19/Y gnd XOR2X1_37/A vdd XNOR2X1
XXOR2X1_297 bloque_bytes[54] bloque_bytes[14] gnd INVX1_549/A vdd XOR2X1
XXNOR2X1_105 AOI21X1_153/C XNOR2X1_105/B gnd BUFX2_164/A vdd XNOR2X1
XNOR2X1_117 NOR2X1_117/A NOR2X1_117/B gnd XOR2X1_108/A vdd NOR2X1
XNAND2X1_198 OR2X2_76/A OR2X2_76/B gnd NAND3X1_176/B vdd NAND2X1
XDFFPOSX1_264 INVX1_220/A CLKBUF1_11/Y INVX1_526/Y gnd vdd DFFPOSX1
XOR2X2_85 OR2X2_85/A OR2X2_85/B gnd OR2X2_85/Y vdd OR2X2
XOAI21X1_625 OR2X2_140/A INVX1_549/A INVX1_575/A gnd NAND2X1_688/A vdd OAI21X1
XAOI21X1_96 AOI21X1_96/A AOI21X1_96/B AOI21X1_96/C gnd NOR2X1_91/A vdd AOI21X1
XINVX1_446 INVX1_446/A gnd INVX1_446/Y vdd INVX1
XXOR2X1_261 INVX1_422/A gnd gnd NOR2X1_322/B vdd XOR2X1
XBUFX2_99 gnd gnd BUFX2_99/Y vdd BUFX2
XAOI21X1_398 NOR3X1_97/Y NOR2X1_450/Y NOR2X1_448/A gnd OAI21X1_644/C vdd AOI21X1
XNAND2X1_162 AND2X2_48/B AND2X2_48/A gnd AOI21X1_101/C vdd NAND2X1
XXOR2X1_1 target[6] XOR2X1_1/B gnd XOR2X1_1/Y vdd XOR2X1
XOR2X2_49 gnd OR2X2_49/B gnd OR2X2_49/Y vdd OR2X2
XAOI21X1_60 NAND3X1_85/A AOI21X1_60/B NAND3X1_79/Y gnd NOR2X1_61/A vdd AOI21X1
XDFFPOSX1_228 INVX1_155/A CLKBUF1_13/Y INVX1_537/A gnd vdd DFFPOSX1
XINVX1_410 INVX1_410/A gnd INVX1_410/Y vdd INVX1
XOAI21X1_589 bloque_bytes[64] INVX1_493/Y OAI21X1_589/C gnd OR2X2_142/A vdd OAI21X1
XNAND2X1_703 NAND2X1_703/A NAND2X1_703/B gnd NAND2X1_703/Y vdd NAND2X1
XXOR2X1_225 INVX1_346/A gnd gnd XOR2X1_225/Y vdd XOR2X1
XFILL_10_8_1 gnd vdd FILL
XFILL_12_6_0 gnd vdd FILL
XBUFX2_63 gnd gnd BUFX2_63/Y vdd BUFX2
XNAND3X1_535 NAND3X1_535/A NAND3X1_533/A NAND3X1_535/C gnd NAND2X1_708/A vdd NAND3X1
XFILL_9_3 gnd vdd FILL
XNAND2X1_126 AOI21X1_77/A AOI21X1_77/B gnd INVX2_28/A vdd NAND2X1
XAOI21X1_362 INVX1_506/Y bloque_bytes[16] AOI21X1_362/C gnd INVX1_508/A vdd AOI21X1
XOR2X2_13 XOR2X1_3/A OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XAOI21X1_24 AOI21X1_24/A AOI21X1_24/B NAND3X1_26/C gnd NOR2X1_31/A vdd AOI21X1
XDFFPOSX1_192 INVX1_105/A CLKBUF1_38/Y bloque_bytes[22] gnd vdd DFFPOSX1
XOAI21X1_553 gnd XOR2X1_282/Y INVX1_457/A gnd INVX1_459/A vdd OAI21X1
XINVX1_374 INVX1_374/A gnd INVX1_374/Y vdd INVX1
XDFFPOSX1_4 BUFX2_3/A CLKBUF1_35/Y NOR3X1_3/Y gnd vdd DFFPOSX1
XNAND2X1_667 INVX1_562/Y NAND2X1_653/B gnd AOI21X1_382/A vdd NAND2X1
XFILL_22_1_0 gnd vdd FILL
XBUFX2_27 gnd gnd BUFX2_27/Y vdd BUFX2
XXOR2X1_189 BUFX2_191/A gnd gnd XOR2X1_189/Y vdd XOR2X1
XNAND2X1_87 OR2X2_29/A OR2X2_29/B gnd NAND3X1_72/B vdd NAND2X1
XFILL_2_2_0 gnd vdd FILL
XAOI21X1_326 INVX1_474/A INVX4_2/Y AND2X2_169/B gnd NOR2X1_386/B vdd AOI21X1
XFILL_20_3_1 gnd vdd FILL
XFILL_0_4_1 gnd vdd FILL
XOAI21X1_72 OAI21X1_69/A NAND2X1_94/Y NOR2X1_55/Y gnd NOR2X1_56/B vdd OAI21X1
XDFFPOSX1_156 INVX1_56/A CLKBUF1_33/Y bloque_bytes[50] gnd vdd DFFPOSX1
XNAND3X1_499 INVX2_78/A INVX2_79/A AND2X2_167/B gnd INVX1_492/A vdd NAND3X1
XDFFPOSX1_90 MUX2X1_1/B CLKBUF1_4/Y BUFX2_26/A gnd vdd DFFPOSX1
XXOR2X1_153 BUFX2_176/A gnd gnd NOR2X1_179/B vdd XOR2X1
XBUFX2_5 BUFX2_5/A gnd hash[4] vdd BUFX2
XINVX1_338 INVX1_338/A gnd INVX1_338/Y vdd INVX1
XOAI21X1_517 INVX1_422/A INVX1_423/A INVX1_424/Y gnd AOI21X1_300/A vdd OAI21X1
XNAND2X1_631 INVX1_481/A INVX1_482/A gnd NOR3X1_89/C vdd NAND2X1
XOAI21X1_36 AND2X2_13/Y NOR2X1_34/Y INVX1_26/A gnd NAND3X1_35/B vdd OAI21X1
XNAND2X1_51 NAND3X1_37/A OR2X2_16/B gnd OR2X2_14/A vdd NAND2X1
XAOI21X1_290 INVX1_394/Y NAND3X1_434/C INVX1_393/A gnd OAI21X1_488/A vdd AOI21X1
XNAND3X1_463 INVX1_439/A NAND2X1_574/Y INVX2_72/Y gnd OAI21X1_537/B vdd NAND3X1
XDFFPOSX1_120 INVX1_596/A CLKBUF1_25/Y bloque_bytes[94] gnd vdd DFFPOSX1
XDFFPOSX1_54 INVX1_572/A CLKBUF1_24/Y NOR2X1_376/Y gnd vdd DFFPOSX1
XOAI21X1_481 NOR2X1_305/Y NOR2X1_304/B AOI22X1_18/C gnd XOR2X1_260/A vdd OAI21X1
XINVX1_302 INVX1_302/A gnd INVX1_302/Y vdd INVX1
XXOR2X1_97 XOR2X1_97/A OR2X2_77/A gnd OR2X2_85/B vdd XOR2X1
XXOR2X1_117 XOR2X1_117/A OR2X2_93/A gnd OR2X2_101/B vdd XOR2X1
XNAND2X1_595 INVX1_457/A NOR2X1_351/Y gnd NAND2X1_595/Y vdd NAND2X1
XAOI21X1_254 OAI21X1_408/Y NAND2X1_449/Y INVX2_65/A gnd AOI21X1_255/B vdd AOI21X1
XFILL_19_6_0 gnd vdd FILL
XNAND3X1_427 INVX1_384/Y INVX1_385/Y INVX1_386/Y gnd NAND3X1_429/B vdd NAND3X1
XNAND2X1_15 AOI22X1_5/Y AOI22X1_6/Y gnd OAI21X1_7/A vdd NAND2X1
XDFFPOSX1_18 BUFX2_17/A CLKBUF1_41/Y NOR3X1_17/Y gnd vdd DFFPOSX1
XAND2X2_197 AND2X2_197/A AND2X2_197/B gnd AND2X2_197/Y vdd AND2X2
XFILL_17_8_1 gnd vdd FILL
XINVX1_266 NOR3X1_65/B gnd INVX1_266/Y vdd INVX1
XOAI21X1_445 BUFX2_212/A XOR2X1_230/Y INVX1_349/A gnd AOI22X1_16/B vdd OAI21X1
XXOR2X1_61 XOR2X1_61/A XOR2X1_61/B gnd XOR2X1_61/Y vdd XOR2X1
XNAND3X1_92 INVX2_24/Y NAND3X1_92/B OAI21X1_85/Y gnd AOI21X1_67/B vdd NAND3X1
XFILL_13_1 gnd vdd FILL
XOR2X2_144 OR2X2_144/A OR2X2_144/B gnd OR2X2_144/Y vdd OR2X2
XNAND2X1_559 AOI21X1_303/A INVX1_427/A gnd NAND2X1_559/Y vdd NAND2X1
XAOI21X1_218 INVX1_223/Y AOI21X1_218/B INVX1_222/A gnd OAI21X1_317/A vdd AOI21X1
XNAND3X1_391 INVX1_331/A NAND3X1_391/B NAND3X1_391/C gnd NAND3X1_391/Y vdd NAND3X1
XFILL_27_3_1 gnd vdd FILL
XFILL_29_1_0 gnd vdd FILL
XNAND3X1_56 INVX2_18/Y NAND3X1_56/B OAI21X1_51/Y gnd NAND3X1_56/Y vdd NAND3X1
XXOR2X1_25 XOR2X1_39/B gnd gnd OR2X2_27/B vdd XOR2X1
XFILL_7_4_1 gnd vdd FILL
XFILL_9_2_0 gnd vdd FILL
XINVX1_230 INVX1_230/A gnd INVX1_230/Y vdd INVX1
XAND2X2_161 BUFX4_31/Y AND2X2_161/B gnd AND2X2_161/Y vdd AND2X2
XNOR2X1_442 INVX1_583/Y NOR2X1_442/B gnd XOR2X1_308/A vdd NOR2X1
XOAI21X1_409 BUFX2_205/A XOR2X1_213/Y INVX1_315/A gnd OAI21X1_409/Y vdd OAI21X1
XOR2X2_108 OR2X2_108/A OR2X2_108/B gnd OR2X2_108/Y vdd OR2X2
XNAND2X1_523 INVX1_387/Y NOR2X1_306/Y gnd INVX1_390/A vdd NAND2X1
XAOI21X1_182 NAND3X1_262/B OR2X2_115/Y INVX1_167/A gnd AOI21X1_182/Y vdd AOI21X1
XNAND3X1_355 INVX1_269/A AOI21X1_236/A AOI21X1_236/B gnd NAND3X1_355/Y vdd NAND3X1
XNAND2X1_4 INVX1_4/A INVX2_5/Y gnd AOI21X1_1/A vdd NAND2X1
XOAI22X1_3 INVX1_3/Y target[1] target[0] INVX1_4/Y gnd NOR2X1_9/A vdd OAI22X1
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_194 INVX1_194/A gnd INVX1_194/Y vdd INVX1
XOAI21X1_373 NOR2X1_233/A NOR3X1_65/Y OAI21X1_373/C gnd NAND3X1_356/C vdd OAI21X1
XFILL_35_1 gnd vdd FILL
XAND2X2_125 AND2X2_125/A AND2X2_125/B gnd AND2X2_125/Y vdd AND2X2
XNAND3X1_20 INVX2_12/Y NAND3X1_20/B NAND2X1_28/B gnd AOI21X1_19/B vdd NAND3X1
XNOR2X1_406 NOR2X1_406/A INVX1_492/A gnd NOR2X1_406/Y vdd NOR2X1
XNAND2X1_487 INVX1_341/A NOR2X1_276/Y gnd NAND2X1_487/Y vdd NAND2X1
XAND2X2_98 AND2X2_98/A AND2X2_98/B gnd NOR3X1_58/A vdd AND2X2
XAOI21X1_146 NAND3X1_208/B OR2X2_91/Y INVX1_134/A gnd AOI21X1_146/Y vdd AOI21X1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XNAND3X1_319 INVX2_61/A NAND3X1_319/B NAND3X1_319/C gnd NOR3X1_61/A vdd NAND3X1
XNOR2X1_370 BUFX4_14/Y INVX2_77/Y gnd NOR2X1_370/Y vdd NOR2X1
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XOAI21X1_337 gnd NOR2X1_214/B INVX1_244/A gnd OAI21X1_337/Y vdd OAI21X1
XFILL_26_6_0 gnd vdd FILL
XNAND2X1_451 INVX1_315/Y NOR2X1_259/Y gnd NAND2X1_452/B vdd NAND2X1
XFILL_4_9_1 gnd vdd FILL
XFILL_6_7_0 gnd vdd FILL
XAOI21X1_110 AOI21X1_110/A OR2X2_67/Y INVX1_101/A gnd NAND3X1_159/C vdd AOI21X1
XAND2X2_62 gnd OR2X2_81/B gnd AND2X2_62/Y vdd AND2X2
XNAND3X1_283 AOI21X1_192/A NAND3X1_283/B NAND3X1_283/C gnd AND2X2_96/B vdd NAND3X1
XFILL_24_8_1 gnd vdd FILL
XINVX1_122 INVX1_122/A gnd NOR3X1_46/A vdd INVX1
XOAI21X1_301 NOR3X1_60/C INVX2_60/Y NOR3X1_60/A gnd AND2X2_104/A vdd OAI21X1
XNAND2X1_415 INVX1_276/Y NOR2X1_236/B gnd NAND2X1_416/A vdd NAND2X1
XNOR2X1_334 gnd XOR2X1_270/Y gnd NOR2X1_334/Y vdd NOR2X1
XFILL_36_1_0 gnd vdd FILL
XFILL_34_3_1 gnd vdd FILL
XBUFX2_248 OR2X2_37/A gnd BUFX2_248/Y vdd BUFX2
XAND2X2_26 gnd OR2X2_33/B gnd AND2X2_26/Y vdd AND2X2
XNAND3X1_247 AOI21X1_168/A NAND3X1_247/B NAND3X1_247/C gnd AND2X2_84/B vdd NAND3X1
XOAI21X1_265 AND2X2_93/Y NOR3X1_56/B NOR3X1_56/A gnd NAND3X1_279/B vdd OAI21X1
XBUFX4_11 BUFX4_8/A gnd MUX2X1_3/S vdd BUFX4
XNAND2X1_379 NAND3X1_329/Y AOI22X1_10/C gnd AOI21X1_225/C vdd NAND2X1
XINVX2_86 bloque_bytes[37] gnd INVX2_86/Y vdd INVX2
XNOR2X1_298 gnd XOR2X1_243/Y gnd NOR2X1_298/Y vdd NOR2X1
XNAND3X1_211 AOI21X1_144/A NAND3X1_211/B NAND3X1_211/C gnd AND2X2_72/B vdd NAND3X1
XNOR2X1_65 NOR2X1_65/A INVX1_60/Y gnd NOR2X1_65/Y vdd NOR2X1
XXNOR2X1_250 NAND2X1_703/B NAND2X1_608/Y gnd DFFPOSX1_97/D vdd XNOR2X1
XBUFX2_212 BUFX2_212/A gnd BUFX2_212/Y vdd BUFX2
XINVX2_50 INVX2_50/A gnd INVX2_50/Y vdd INVX2
XOAI21X1_229 NOR3X1_51/C NOR3X1_51/B INVX1_154/Y gnd NAND2X1_269/A vdd OAI21X1
XNOR2X1_262 gnd NOR2X1_262/B gnd AND2X2_126/A vdd NOR2X1
XNAND2X1_343 INVX1_206/Y AND2X2_102/A gnd NAND3X1_306/B vdd NAND2X1
XINVX1_591 INVX1_591/A gnd NOR3X1_98/A vdd INVX1
XBUFX2_176 BUFX2_176/A gnd BUFX2_176/Y vdd BUFX2
XNAND3X1_175 NAND3X1_175/A NAND3X1_174/Y NAND3X1_175/C gnd AND2X2_60/B vdd NAND3X1
XNOR2X1_29 gnd AND2X2_9/B gnd NOR3X1_28/B vdd NOR2X1
XOAI21X1_193 AOI21X1_142/Y OAI21X1_193/B INVX1_128/Y gnd NAND3X1_202/C vdd OAI21X1
XXNOR2X1_214 bloque_bytes[40] bloque_bytes[0] gnd NAND2X1_657/A vdd XNOR2X1
XFILL_33_6_0 gnd vdd FILL
XFILL_31_8_1 gnd vdd FILL
XINVX2_14 INVX2_14/A gnd INVX2_14/Y vdd INVX2
XNAND2X1_307 OAI21X1_263/Y NAND3X1_276/A gnd XNOR2X1_141/A vdd NAND2X1
XNOR2X1_226 gnd XOR2X1_189/Y gnd AND2X2_114/A vdd NOR2X1
XBUFX2_140 gnd gnd BUFX2_140/Y vdd BUFX2
XCLKBUF1_17 BUFX4_1/Y gnd CLKBUF1_17/Y vdd CLKBUF1
XNAND3X1_139 AOI21X1_96/A NAND3X1_138/Y OAI21X1_134/Y gnd AND2X2_48/B vdd NAND3X1
XINVX1_555 INVX1_555/A gnd INVX1_555/Y vdd INVX1
XXNOR2X1_178 NOR2X1_273/Y XNOR2X1_178/B gnd XNOR2X1_178/Y vdd XNOR2X1
XOAI21X1_157 XNOR2X1_80/A NAND2X1_189/Y NOR2X1_105/Y gnd NOR2X1_106/B vdd OAI21X1
XNOR2X1_190 gnd XOR2X1_162/Y gnd AND2X2_102/A vdd NOR2X1
XNAND2X1_271 NAND2X1_271/A OAI21X1_230/Y gnd XNOR2X1_124/A vdd NAND2X1
XNAND3X1_103 OAI21X1_98/Y NAND3X1_102/Y OAI21X1_100/Y gnd AND2X2_36/B vdd NAND3X1
XINVX1_519 INVX1_519/A gnd INVX1_519/Y vdd INVX1
XDFFPOSX1_337 XNOR2X1_190/B CLKBUF1_22/Y OR2X2_149/Y gnd vdd DFFPOSX1
XNOR3X1_70 NOR3X1_70/A INVX2_65/Y NOR3X1_70/C gnd NOR3X1_70/Y vdd NOR3X1
XBUFX2_104 gnd gnd BUFX2_104/Y vdd BUFX2
XXNOR2X1_142 XNOR2X1_142/A XNOR2X1_142/B gnd BUFX2_181/A vdd XNOR2X1
XOAI21X1_121 AND2X2_43/Y NOR2X1_84/Y INVX1_81/A gnd OAI21X1_121/Y vdd OAI21X1
XXNOR2X1_64 XOR2X1_54/A XOR2X1_58/Y gnd OR2X2_55/A vdd XNOR2X1
XNOR2X1_154 BUFX2_164/A OR2X2_109/B gnd NOR2X1_154/Y vdd NOR2X1
XNOR3X1_34 INVX1_56/Y NOR3X1_34/B NOR3X1_34/C gnd NOR2X1_63/B vdd NOR3X1
XFILL_15_1_1 gnd vdd FILL
XNAND2X1_235 gnd OR2X2_91/B gnd NAND3X1_208/B vdd NAND2X1
XINVX1_483 INVX1_483/A gnd NOR3X1_92/A vdd INVX1
XDFFPOSX1_301 INVX1_305/A CLKBUF1_34/Y INVX1_550/Y gnd vdd DFFPOSX1
XXNOR2X1_28 XOR2X1_28/B XOR2X1_18/Y gnd OR2X2_23/A vdd XNOR2X1
XXOR2X1_298 bloque_bytes[64] bloque_bytes[24] gnd NOR2X1_410/B vdd XOR2X1
XXNOR2X1_106 XNOR2X1_106/A XNOR2X1_106/B gnd BUFX2_165/A vdd XNOR2X1
XNOR2X1_118 gnd OR2X2_81/B gnd NOR3X1_45/B vdd NOR2X1
XNAND2X1_199 INVX2_39/Y OAI21X1_170/Y gnd XNOR2X1_89/A vdd NAND2X1
XDFFPOSX1_265 XNOR2X1_154/B CLKBUF1_11/Y INVX1_529/Y gnd vdd DFFPOSX1
XAOI21X1_97 AOI21X1_97/A AOI21X1_97/B NOR3X1_40/Y gnd INVX2_33/A vdd AOI21X1
XOR2X2_86 OR2X2_86/A OR2X2_86/B gnd OR2X2_86/Y vdd OR2X2
XOAI21X1_626 NOR2X1_431/Y OAI21X1_626/B INVX1_568/A gnd OAI21X1_626/Y vdd OAI21X1
XXOR2X1_262 BUFX2_228/A gnd gnd NOR2X1_323/B vdd XOR2X1
XINVX1_447 INVX1_447/A gnd INVX1_447/Y vdd INVX1
XXOR2X1_2 XOR2X1_2/A gnd gnd XOR2X1_2/Y vdd XOR2X1
XAOI21X1_399 NAND3X1_541/B OR2X2_158/Y INVX1_593/A gnd OR2X2_160/B vdd AOI21X1
XNAND2X1_163 OR2X2_61/A OR2X2_61/B gnd NAND2X1_163/Y vdd NAND2X1
XOR2X2_50 gnd OR2X2_50/B gnd OR2X2_50/Y vdd OR2X2
XAOI21X1_61 AOI21X1_61/A AOI21X1_61/B NOR2X1_63/B gnd INVX2_24/A vdd AOI21X1
XOAI21X1_590 bloque_bytes[65] INVX1_494/Y OAI21X1_590/C gnd OR2X2_143/A vdd OAI21X1
XDFFPOSX1_229 INVX1_156/A CLKBUF1_10/Y AOI21X1_353/C gnd vdd DFFPOSX1
XINVX1_411 INVX1_411/A gnd INVX1_411/Y vdd INVX1
XNAND2X1_704 INVX2_92/Y XNOR2X1_252/A gnd NAND2X1_704/Y vdd NAND2X1
XFILL_14_4_0 gnd vdd FILL
XXOR2X1_226 BUFX2_212/A gnd gnd NOR2X1_275/B vdd XOR2X1
XBUFX2_64 gnd gnd BUFX2_64/Y vdd BUFX2
XNAND2X1_127 OAI21X1_105/Y OR2X2_48/B gnd OR2X2_46/A vdd NAND2X1
XFILL_12_6_1 gnd vdd FILL
XAOI21X1_363 INVX1_509/Y bloque_bytes[17] AOI21X1_363/C gnd INVX1_511/A vdd AOI21X1
XNAND3X1_536 NAND3X1_535/C NAND3X1_535/A NOR3X1_97/Y gnd INVX1_598/A vdd NAND3X1
XDFFPOSX1_193 XOR2X1_91/B CLKBUF1_37/Y bloque_bytes[23] gnd vdd DFFPOSX1
XDFFPOSX1_5 BUFX2_4/A CLKBUF1_4/Y NOR3X1_4/Y gnd vdd DFFPOSX1
XOR2X2_14 OR2X2_14/A OR2X2_14/B gnd INVX1_27/A vdd OR2X2
XAOI21X1_25 AOI21X1_25/A AOI21X1_25/B NOR2X1_33/B gnd INVX2_15/A vdd AOI21X1
XOAI21X1_554 INVX1_460/A INVX1_461/A INVX1_462/A gnd INVX1_464/A vdd OAI21X1
XINVX1_375 INVX1_375/A gnd INVX1_375/Y vdd INVX1
XBUFX2_28 gnd gnd BUFX2_28/Y vdd BUFX2
XFILL_4_0_0 gnd vdd FILL
XFILL_22_1_1 gnd vdd FILL
XNAND2X1_668 bloque_bytes[4] OR2X2_153/B gnd AOI21X1_383/B vdd NAND2X1
XXOR2X1_190 BUFX2_192/A gnd gnd XOR2X1_190/Y vdd XOR2X1
XNAND2X1_88 AOI21X1_53/A AOI21X1_53/B gnd INVX2_22/A vdd NAND2X1
XFILL_2_2_1 gnd vdd FILL
XAOI21X1_327 AOI21X1_327/A AOI21X1_327/B BUFX4_13/Y gnd DFFPOSX1_65/D vdd AOI21X1
XNAND3X1_500 INVX1_483/A INVX1_492/Y NOR3X1_90/Y gnd AOI21X1_346/B vdd NAND3X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XOAI21X1_73 INVX2_22/Y AND2X2_24/B INVX1_49/A gnd OAI21X1_74/B vdd OAI21X1
XDFFPOSX1_157 INVX1_57/A CLKBUF1_33/Y bloque_bytes[51] gnd vdd DFFPOSX1
XDFFPOSX1_91 MUX2X1_2/B CLKBUF1_13/Y INVX1_585/Y gnd vdd DFFPOSX1
XXOR2X1_154 BUFX2_177/A gnd gnd NOR2X1_180/B vdd XOR2X1
XBUFX2_6 BUFX2_6/A gnd hash[5] vdd BUFX2
XINVX1_339 INVX1_339/A gnd INVX1_339/Y vdd INVX1
XOAI21X1_518 NOR3X1_81/C OAI21X1_512/C INVX1_427/A gnd NOR2X1_329/A vdd OAI21X1
XNAND2X1_632 AND2X2_168/Y AND2X2_169/Y gnd NOR3X1_91/B vdd NAND2X1
XNAND2X1_52 INVX1_28/Y OR2X2_15/A gnd NAND2X1_53/A vdd NAND2X1
XOAI21X1_37 AND2X2_13/Y NOR2X1_34/Y INVX1_26/Y gnd NAND3X1_37/A vdd OAI21X1
XFILL_11_9_0 gnd vdd FILL
XDFFPOSX1_55 INVX2_88/A CLKBUF1_24/Y NOR2X1_377/Y gnd vdd DFFPOSX1
XNAND3X1_464 INVX1_439/A OAI21X1_533/Y NAND2X1_576/Y gnd NAND3X1_464/Y vdd NAND3X1
XAOI21X1_291 INVX1_407/A NAND3X1_440/Y INVX1_402/Y gnd NOR2X1_316/B vdd AOI21X1
XDFFPOSX1_121 XOR2X1_318/B CLKBUF1_5/Y bloque_bytes[95] gnd vdd DFFPOSX1
XINVX1_303 INVX1_303/A gnd INVX1_303/Y vdd INVX1
XOAI21X1_482 BUFX2_220/A NOR2X1_306/B INVX1_387/Y gnd OAI21X1_482/Y vdd OAI21X1
XXOR2X1_98 XOR2X1_98/A XOR2X1_98/B gnd XOR2X1_98/Y vdd XOR2X1
XXOR2X1_118 XOR2X1_118/A BUFX2_157/A gnd XOR2X1_118/Y vdd XOR2X1
XNAND2X1_596 INVX1_457/Y NOR2X1_351/Y gnd AOI21X1_317/B vdd NAND2X1
XAOI21X1_255 AOI21X1_255/A AOI21X1_255/B INVX1_313/Y gnd AOI21X1_256/A vdd AOI21X1
XFILL_1_5_0 gnd vdd FILL
XFILL_19_6_1 gnd vdd FILL
XFILL_21_4_0 gnd vdd FILL
XNAND3X1_428 INVX1_386/A INVX1_384/Y INVX1_385/Y gnd NAND3X1_433/C vdd NAND3X1
XNAND2X1_16 INVX1_10/A INVX2_5/Y gnd AND2X2_1/A vdd NAND2X1
XDFFPOSX1_19 BUFX2_18/A CLKBUF1_42/Y NOR3X1_18/Y gnd vdd DFFPOSX1
XAND2X2_198 gnd gnd gnd AND2X2_198/Y vdd AND2X2
XXOR2X1_62 OR2X2_60/A gnd gnd XOR2X1_62/Y vdd XOR2X1
XINVX1_267 INVX1_267/A gnd INVX1_267/Y vdd INVX1
XOAI21X1_446 gnd NOR2X1_276/B INVX1_341/Y gnd OAI21X1_446/Y vdd OAI21X1
XNAND3X1_93 NAND3X1_93/A XNOR2X1_43/A XOR2X1_50/B gnd NAND3X1_93/Y vdd NAND3X1
XFILL_13_2 gnd vdd FILL
XOR2X2_145 OR2X2_145/A INVX1_501/A gnd OR2X2_145/Y vdd OR2X2
XNAND2X1_560 INVX1_425/A NOR2X1_330/Y gnd NAND2X1_560/Y vdd NAND2X1
XAOI21X1_219 INVX1_236/A NAND3X1_323/Y INVX1_231/Y gnd NOR2X1_208/B vdd AOI21X1
XNAND3X1_392 AOI22X1_15/B INVX1_333/A INVX1_331/Y gnd AOI21X1_265/B vdd NAND3X1
XFILL_29_1_1 gnd vdd FILL
XFILL_9_2_1 gnd vdd FILL
XINVX1_231 INVX1_231/A gnd INVX1_231/Y vdd INVX1
XXOR2X1_26 XOR2X1_26/A OR2X2_20/A gnd OR2X2_28/B vdd XOR2X1
XNAND3X1_57 NAND3X1_57/A XNOR2X1_25/A XOR2X1_30/B gnd AOI21X1_46/B vdd NAND3X1
XAND2X2_162 BUFX4_31/Y AND2X2_162/B gnd AND2X2_162/Y vdd AND2X2
XNAND2X1_524 NAND2X1_524/A NAND2X1_524/B gnd XOR2X1_260/B vdd NAND2X1
XOAI21X1_410 OAI21X1_410/A INVX1_318/A INVX1_317/Y gnd AND2X2_125/A vdd OAI21X1
XNOR2X1_443 INVX1_585/A NOR2X1_350/Y gnd INVX1_586/A vdd NOR2X1
XAOI21X1_183 NOR3X1_53/Y NOR2X1_163/Y NOR2X1_161/A gnd AOI21X1_183/Y vdd AOI21X1
XOR2X2_109 BUFX2_164/A OR2X2_109/B gnd OR2X2_109/Y vdd OR2X2
XNAND2X1_5 INVX1_3/A INVX2_4/Y gnd AOI21X1_1/B vdd NAND2X1
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XNAND3X1_356 INVX1_280/Y INVX1_279/A NAND3X1_356/C gnd AND2X2_117/B vdd NAND3X1
XOAI22X1_4 INVX2_4/Y INVX1_3/A INVX2_5/Y INVX1_4/A gnd NOR2X1_9/B vdd OAI22X1
XINVX1_195 INVX1_195/A gnd INVX1_195/Y vdd INVX1
XOAI21X1_374 AOI21X1_242/Y INVX1_278/A INVX1_281/A gnd OAI21X1_374/Y vdd OAI21X1
XAND2X2_126 AND2X2_126/A INVX1_320/Y gnd NOR3X1_72/A vdd AND2X2
XFILL_35_2 gnd vdd FILL
XNAND3X1_21 NAND3X1_21/A XNOR2X1_7/A XOR2X1_10/B gnd AOI21X1_22/B vdd NAND3X1
XNOR2X1_407 INVX2_81/Y OR2X2_130/A gnd NOR2X1_407/Y vdd NOR2X1
XFILL_18_9_0 gnd vdd FILL
XNAND2X1_488 XOR2X1_242/B NOR2X1_280/Y gnd AOI21X1_272/C vdd NAND2X1
XAND2X2_99 AND2X2_99/A AND2X2_99/B gnd NOR3X1_58/C vdd AND2X2
XNAND3X1_320 INVX1_230/A NAND2X1_365/Y INVX2_61/Y gnd OAI21X1_328/B vdd NAND3X1
XAOI21X1_147 NOR3X1_47/Y NOR2X1_133/Y NOR2X1_131/A gnd OAI21X1_204/C vdd AOI21X1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XNOR2X1_371 BUFX4_14/Y INVX1_481/Y gnd NOR2X1_371/Y vdd NOR2X1
XOAI21X1_338 gnd NOR2X1_215/B INVX1_245/A gnd INVX2_62/A vdd OAI21X1
XINVX1_159 INVX1_159/A gnd INVX1_159/Y vdd INVX1
XFILL_28_4_0 gnd vdd FILL
XFILL_8_5_0 gnd vdd FILL
XFILL_26_6_1 gnd vdd FILL
XNAND2X1_452 OAI21X1_409/Y NAND2X1_452/B gnd NOR2X1_260/B vdd NAND2X1
XFILL_6_7_1 gnd vdd FILL
XAOI21X1_111 NOR3X1_41/Y NOR2X1_103/Y NOR2X1_101/A gnd OAI21X1_153/C vdd AOI21X1
XAND2X2_63 gnd OR2X2_82/B gnd NOR3X1_46/C vdd AND2X2
XNAND3X1_284 INVX1_179/A AOI21X1_196/A OR2X2_124/Y gnd NAND3X1_285/B vdd NAND3X1
XINVX1_123 INVX1_123/A gnd INVX1_123/Y vdd INVX1
XOAI21X1_302 gnd NOR2X1_192/B INVX1_208/A gnd INVX1_211/A vdd OAI21X1
XNAND2X1_416 NAND2X1_416/A INVX1_278/Y gnd INVX1_279/A vdd NAND2X1
XNOR2X1_335 gnd XOR2X1_271/Y gnd NOR2X1_335/Y vdd NOR2X1
XFILL_36_1_1 gnd vdd FILL
XAND2X2_27 gnd OR2X2_34/B gnd NOR3X1_34/C vdd AND2X2
XBUFX2_249 BUFX2_249/A gnd BUFX2_249/Y vdd BUFX2
XNAND3X1_248 INVX1_157/A NAND3X1_248/B OR2X2_108/Y gnd NAND3X1_249/B vdd NAND3X1
XOAI21X1_266 NOR3X1_56/Y NOR2X1_173/A NAND3X1_276/A gnd NAND2X1_310/B vdd OAI21X1
XBUFX4_12 BUFX4_8/A gnd MUX2X1_8/S vdd BUFX4
XNOR2X1_299 gnd XOR2X1_244/Y gnd NOR2X1_299/Y vdd NOR2X1
XNAND2X1_380 NAND2X1_380/A NAND3X1_331/Y gnd XOR2X1_196/A vdd NAND2X1
XINVX2_87 bloque_bytes[38] gnd INVX2_87/Y vdd INVX2
XNAND3X1_212 INVX1_135/A AOI21X1_148/A OR2X2_92/Y gnd NAND3X1_213/B vdd NAND3X1
XFILL_25_9_0 gnd vdd FILL
XBUFX2_213 BUFX2_213/A gnd BUFX2_213/Y vdd BUFX2
XXNOR2X1_251 vdd vdd gnd XNOR2X1_252/A vdd XNOR2X1
XNOR2X1_66 INVX1_62/Y NOR2X1_66/B gnd NOR2X1_66/Y vdd NOR2X1
XNAND2X1_344 NAND2X1_344/A NAND3X1_306/B gnd INVX1_251/A vdd NAND2X1
XINVX2_51 INVX2_51/A gnd INVX2_51/Y vdd INVX2
XOAI21X1_230 NOR3X1_52/Y NOR2X1_153/A NOR3X1_51/Y gnd OAI21X1_230/Y vdd OAI21X1
XNOR2X1_263 gnd XOR2X1_217/Y gnd AND2X2_127/A vdd NOR2X1
XINVX1_592 INVX1_592/A gnd INVX1_592/Y vdd INVX1
XBUFX2_177 BUFX2_177/A gnd BUFX2_177/Y vdd BUFX2
XNAND3X1_176 INVX1_113/A NAND3X1_176/B OR2X2_76/Y gnd NAND3X1_177/B vdd NAND3X1
XFILL_35_4_0 gnd vdd FILL
XFILL_33_6_1 gnd vdd FILL
XNOR2X1_30 gnd OR2X2_11/B gnd NOR2X1_30/Y vdd NOR2X1
XOAI21X1_194 NOR2X1_127/A INVX1_130/Y INVX1_131/Y gnd OAI21X1_194/Y vdd OAI21X1
XXNOR2X1_215 bloque_bytes[41] bloque_bytes[1] gnd XNOR2X1_215/Y vdd XNOR2X1
XINVX2_15 INVX2_15/A gnd INVX2_15/Y vdd INVX2
XNAND2X1_308 gnd OR2X2_122/B gnd AOI21X1_191/A vdd NAND2X1
XNOR2X1_227 gnd XOR2X1_190/Y gnd AND2X2_115/A vdd NOR2X1
XBUFX2_141 gnd gnd BUFX2_141/Y vdd BUFX2
XNAND3X1_140 INVX1_91/A AOI21X1_100/A OR2X2_60/Y gnd NAND3X1_140/Y vdd NAND3X1
XCLKBUF1_18 BUFX4_4/Y gnd CLKBUF1_18/Y vdd CLKBUF1
XINVX1_556 INVX1_556/A gnd INVX1_556/Y vdd INVX1
XXNOR2X1_179 XNOR2X1_178/Y OAI21X1_428/Y gnd INVX1_338/A vdd XNOR2X1
XOAI21X1_158 INVX2_37/Y AND2X2_54/B OR2X2_70/Y gnd OAI21X1_158/Y vdd OAI21X1
XNOR2X1_191 gnd NOR2X1_191/B gnd AND2X2_103/A vdd NOR2X1
XNAND2X1_272 INVX1_162/A NAND2X1_272/B gnd OAI21X1_233/A vdd NAND2X1
XNOR3X1_71 NOR3X1_71/A NOR3X1_71/B NOR3X1_71/C gnd NOR3X1_71/Y vdd NOR3X1
XNAND3X1_104 INVX1_69/A AOI21X1_76/A OR2X2_44/Y gnd NAND3X1_104/Y vdd NAND3X1
XINVX1_520 INVX1_520/A gnd INVX1_520/Y vdd INVX1
XDFFPOSX1_338 INVX1_396/A CLKBUF1_51/Y NAND2X1_683/Y gnd vdd DFFPOSX1
XBUFX2_105 gnd gnd BUFX2_105/Y vdd BUFX2
XOAI21X1_122 AND2X2_43/Y NOR2X1_84/Y INVX1_81/Y gnd OAI21X1_122/Y vdd OAI21X1
XXNOR2X1_65 XOR2X1_71/Y XOR2X1_59/Y gnd XNOR2X1_66/A vdd XNOR2X1
XXNOR2X1_143 XNOR2X1_143/A AND2X2_96/Y gnd XOR2X1_166/A vdd XNOR2X1
XNAND2X1_236 OR2X2_92/A OR2X2_92/B gnd AOI21X1_148/A vdd NAND2X1
XNOR2X1_155 NOR2X1_155/A INVX1_159/Y gnd NOR2X1_155/Y vdd NOR2X1
XFILL_32_9_0 gnd vdd FILL
XNOR3X1_35 INVX1_66/Y NOR3X1_35/B NOR3X1_35/C gnd NOR3X1_35/Y vdd NOR3X1
XDFFPOSX1_302 INVX1_310/A CLKBUF1_34/Y INVX1_551/Y gnd vdd DFFPOSX1
XINVX1_484 INVX1_484/A gnd INVX1_484/Y vdd INVX1
XXOR2X1_299 bloque_bytes[65] bloque_bytes[25] gnd NOR2X1_411/B vdd XOR2X1
XXNOR2X1_29 XOR2X1_31/Y XOR2X1_19/Y gnd XNOR2X1_30/A vdd XNOR2X1
XXNOR2X1_107 NAND2X1_237/Y AND2X2_72/Y gnd XOR2X1_126/A vdd XNOR2X1
XNOR2X1_119 gnd OR2X2_82/B gnd NOR3X1_46/B vdd NOR2X1
XNAND2X1_200 AND2X2_60/B AND2X2_60/A gnd AOI21X1_125/C vdd NAND2X1
XOR2X2_87 OR2X2_87/A OR2X2_87/B gnd OR2X2_87/Y vdd OR2X2
XDFFPOSX1_266 INVX1_225/A CLKBUF1_18/Y XNOR2X1_235/A gnd vdd DFFPOSX1
XAOI21X1_98 AOI21X1_98/A OR2X2_59/Y INVX1_90/A gnd AOI21X1_98/Y vdd AOI21X1
XINVX1_448 INVX1_448/A gnd INVX1_448/Y vdd INVX1
XOAI21X1_627 NOR2X1_432/Y OAI21X1_627/B INVX1_569/A gnd OAI21X1_627/Y vdd OAI21X1
XXOR2X1_263 BUFX2_229/A gnd gnd NOR2X1_324/B vdd XOR2X1
XXOR2X1_3 XOR2X1_3/A gnd gnd OR2X2_9/B vdd XOR2X1
XAOI21X1_400 AOI21X1_400/A AOI21X1_400/B AOI21X1_400/C gnd NAND3X1_547/B vdd AOI21X1
XNAND2X1_164 NAND3X1_143/Y NAND3X1_145/Y gnd INVX2_34/A vdd NAND2X1
XFILL_26_1 gnd vdd FILL
XOR2X2_51 gnd OR2X2_51/B gnd OR2X2_51/Y vdd OR2X2
XAOI21X1_62 NAND3X1_83/B OR2X2_35/Y INVX1_57/A gnd AOI21X1_62/Y vdd AOI21X1
XFILL_16_2_0 gnd vdd FILL
XOAI21X1_591 bloque_bytes[66] INVX1_495/Y OAI21X1_591/C gnd OAI21X1_591/Y vdd OAI21X1
XDFFPOSX1_230 INVX1_157/A CLKBUF1_10/Y AOI21X1_354/C gnd vdd DFFPOSX1
XINVX1_412 INVX1_412/A gnd INVX1_412/Y vdd INVX1
XNAND2X1_705 gnd gnd gnd NAND2X1_705/Y vdd NAND2X1
XFILL_14_4_1 gnd vdd FILL
XBUFX2_65 gnd gnd BUFX2_65/Y vdd BUFX2
XXOR2X1_227 BUFX2_213/A gnd gnd NOR2X1_276/B vdd XOR2X1
XNAND3X1_537 INVX1_592/A NAND3X1_537/B OR2X2_157/Y gnd AOI21X1_395/B vdd NAND3X1
XNAND2X1_128 INVX1_72/Y OR2X2_47/A gnd NAND2X1_129/A vdd NAND2X1
XAOI21X1_364 INVX1_512/Y bloque_bytes[18] OAI21X1_603/Y gnd INVX1_514/A vdd AOI21X1
XAOI21X1_26 NAND3X1_28/B OR2X2_11/Y INVX1_24/A gnd AOI21X1_26/Y vdd AOI21X1
XDFFPOSX1_194 INVX2_38/A CLKBUF1_10/Y bloque_bytes[8] gnd vdd DFFPOSX1
XDFFPOSX1_6 BUFX2_5/A CLKBUF1_35/Y NOR3X1_5/Y gnd vdd DFFPOSX1
XOR2X2_15 OR2X2_15/A INVX1_28/Y gnd OR2X2_15/Y vdd OR2X2
XXOR2X1_191 BUFX2_193/A gnd gnd NOR2X1_228/B vdd XOR2X1
XOAI21X1_555 INVX1_460/A INVX1_461/A INVX1_462/Y gnd OAI21X1_555/Y vdd OAI21X1
XINVX1_376 INVX1_376/A gnd INVX1_376/Y vdd INVX1
XFILL_4_0_1 gnd vdd FILL
XNAND2X1_669 INVX1_564/Y AOI21X1_374/Y gnd AOI21X1_383/A vdd NAND2X1
XBUFX2_29 gnd gnd BUFX2_29/Y vdd BUFX2
XNAND2X1_89 NAND3X1_73/A OR2X2_32/B gnd OR2X2_30/A vdd NAND2X1
XOAI21X1_74 OAI21X1_74/A OAI21X1_74/B INVX1_51/Y gnd OAI21X1_74/Y vdd OAI21X1
XNAND3X1_501 INVX2_84/Y NOR2X1_406/Y NOR3X1_94/Y gnd NAND3X1_501/Y vdd NAND3X1
XAOI21X1_328 AND2X2_161/B INVX2_82/Y AOI21X1_328/C gnd DFFPOSX1_66/D vdd AOI21X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XDFFPOSX1_158 INVX1_58/A CLKBUF1_33/Y bloque_bytes[52] gnd vdd DFFPOSX1
XDFFPOSX1_92 MUX2X1_3/B CLKBUF1_35/Y DFFPOSX1_92/D gnd vdd DFFPOSX1
XINVX1_340 INVX1_340/A gnd INVX1_340/Y vdd INVX1
XOAI21X1_519 NOR2X1_329/Y NOR2X1_328/B AOI22X1_20/C gnd XOR2X1_278/A vdd OAI21X1
XNAND2X1_633 NOR2X1_387/Y NOR2X1_388/Y gnd NOR3X1_94/C vdd NAND2X1
XXOR2X1_155 BUFX2_178/A gnd gnd NOR2X1_183/B vdd XOR2X1
XBUFX2_7 BUFX2_7/A gnd hash[6] vdd BUFX2
XAOI21X1_292 NAND3X1_446/B NAND3X1_441/Y INVX1_402/A gnd NOR2X1_316/A vdd AOI21X1
XNAND2X1_53 NAND2X1_53/A OR2X2_15/Y gnd OR2X2_16/A vdd NAND2X1
XDFFPOSX1_122 INVX2_11/A CLKBUF1_5/Y bloque_bytes[80] gnd vdd DFFPOSX1
XOAI21X1_38 OAI21X1_35/A AOI21X1_34/C NOR2X1_35/Y gnd NOR2X1_36/B vdd OAI21X1
XFILL_11_9_1 gnd vdd FILL
XDFFPOSX1_56 INVX2_89/A CLKBUF1_24/Y NOR2X1_378/Y gnd vdd DFFPOSX1
XFILL_13_7_0 gnd vdd FILL
XNAND3X1_465 INVX1_440/A AOI21X1_309/B INVX1_439/Y gnd INVX1_446/A vdd NAND3X1
XINVX1_304 NOR3X1_69/B gnd INVX1_304/Y vdd INVX1
XOAI21X1_483 BUFX2_220/A NOR2X1_306/B INVX1_387/A gnd AOI22X1_18/B vdd OAI21X1
XXOR2X1_99 XOR2X1_99/A XOR2X1_99/B gnd XOR2X1_99/Y vdd XOR2X1
XXOR2X1_119 XOR2X1_119/A BUFX2_158/A gnd XOR2X1_119/Y vdd XOR2X1
XNAND2X1_597 NAND3X1_477/Y INVX1_465/A gnd NAND2X1_597/Y vdd NAND2X1
XFILL_21_4_1 gnd vdd FILL
XFILL_23_2_0 gnd vdd FILL
XNAND3X1_429 INVX1_388/A NAND3X1_429/B INVX1_383/Y gnd AOI22X1_18/C vdd NAND3X1
XAOI21X1_256 AOI21X1_256/A AOI21X1_256/B NAND2X1_450/Y gnd OAI21X1_410/A vdd AOI21X1
XNAND2X1_17 MUX2X1_18/B INVX2_4/Y gnd AND2X2_1/B vdd NAND2X1
XFILL_1_5_1 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XDFFPOSX1_20 BUFX2_19/A CLKBUF1_48/Y NOR3X1_19/Y gnd vdd DFFPOSX1
XNAND3X1_94 OR2X2_40/Y INVX1_65/A NAND3X1_94/C gnd NAND3X1_94/Y vdd NAND3X1
XXOR2X1_63 OR2X2_61/A gnd gnd OR2X2_57/B vdd XOR2X1
XOAI21X1_447 BUFX2_213/A XOR2X1_231/Y INVX1_353/A gnd OAI21X1_447/Y vdd OAI21X1
XINVX1_268 INVX1_268/A gnd INVX1_268/Y vdd INVX1
XOR2X2_146 OR2X2_151/A INVX1_502/A gnd OR2X2_146/Y vdd OR2X2
XNAND2X1_561 INVX1_425/Y NOR2X1_330/Y gnd INVX1_428/A vdd NAND2X1
XAOI21X1_220 OAI21X1_327/Y NAND3X1_324/Y INVX1_231/A gnd NOR2X1_208/A vdd AOI21X1
XNAND3X1_393 INVX1_323/Y NAND3X1_386/Y NOR3X1_72/Y gnd AOI21X1_264/B vdd NAND3X1
XINVX1_232 BUFX2_183/A gnd INVX1_232/Y vdd INVX1
XAND2X2_163 BUFX4_32/Y AND2X2_163/B gnd AND2X2_163/Y vdd AND2X2
XOAI21X1_411 NOR2X1_257/A NOR3X1_69/Y AOI21X1_257/Y gnd NAND3X1_382/C vdd OAI21X1
XXOR2X1_27 XOR2X1_27/A OR2X2_21/A gnd OR2X2_29/B vdd XOR2X1
XNAND3X1_58 OR2X2_24/Y INVX1_43/A OAI21X1_57/Y gnd NAND3X1_58/Y vdd NAND3X1
XOR2X2_110 OR2X2_110/A OR2X2_110/B gnd INVX1_159/A vdd OR2X2
XNOR2X1_444 XOR2X1_296/Y NOR2X1_444/B gnd NOR2X1_444/Y vdd NOR2X1
XNAND2X1_525 INVX1_379/A NOR2X1_300/Y gnd NAND2X1_525/Y vdd NAND2X1
XAOI21X1_184 NAND3X1_264/B OR2X2_116/Y INVX1_168/A gnd OR2X2_118/B vdd AOI21X1
XNAND2X1_6 NOR2X1_4/A INVX2_6/Y gnd NAND2X1_6/Y vdd NAND2X1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XNAND3X1_357 INVX1_278/Y INVX1_281/Y AND2X2_117/A gnd NAND2X1_418/B vdd NAND3X1
XOAI22X1_5 INVX2_6/Y INVX2_10/A INVX1_9/A INVX2_7/Y gnd NOR2X1_15/A vdd OAI22X1
XINVX1_196 INVX1_196/A gnd INVX1_196/Y vdd INVX1
XNOR2X1_408 bloque_bytes[53] bloque_bytes[13] gnd NOR2X1_408/Y vdd NOR2X1
XFILL_20_7_0 gnd vdd FILL
XOAI21X1_375 gnd XOR2X1_198/Y INVX1_282/A gnd NAND2X1_420/A vdd OAI21X1
XAND2X2_127 AND2X2_127/A INVX1_321/Y gnd NOR3X1_72/C vdd AND2X2
XFILL_35_3 gnd vdd FILL
XFILL_0_8_0 gnd vdd FILL
XNAND3X1_22 OR2X2_8/Y INVX1_21/A NAND3X1_22/C gnd NAND2X1_38/A vdd NAND3X1
XFILL_18_9_1 gnd vdd FILL
XNAND2X1_489 INVX1_353/Y NOR2X1_283/Y gnd NAND2X1_490/B vdd NAND2X1
XNAND3X1_321 INVX1_230/A OAI21X1_324/Y NAND3X1_321/C gnd AOI21X1_223/A vdd NAND3X1
XAOI21X1_148 AOI21X1_148/A OR2X2_92/Y INVX1_135/A gnd OR2X2_94/B vdd AOI21X1
XINVX1_42 OR2X2_24/Y gnd INVX1_42/Y vdd INVX1
XINVX1_160 INVX1_160/A gnd INVX1_160/Y vdd INVX1
XFILL_30_2_0 gnd vdd FILL
XNOR2X1_372 BUFX4_17/Y INVX1_482/Y gnd NOR2X1_372/Y vdd NOR2X1
XOAI21X1_339 NOR3X1_64/C INVX2_62/Y NOR3X1_64/A gnd AND2X2_112/A vdd OAI21X1
XNAND2X1_453 INVX1_314/Y NOR2X1_260/B gnd NAND2X1_454/A vdd NAND2X1
XFILL_28_4_1 gnd vdd FILL
XAOI21X1_112 NAND2X1_179/Y OR2X2_68/Y INVX1_102/A gnd OR2X2_70/B vdd AOI21X1
XFILL_8_5_1 gnd vdd FILL
XNAND3X1_285 NAND3X1_287/A NAND3X1_285/B AOI21X1_194/Y gnd AND2X2_96/A vdd NAND3X1
XAND2X2_64 gnd OR2X2_83/B gnd AND2X2_64/Y vdd AND2X2
XOAI21X1_303 NOR3X1_59/A NOR3X1_59/B OAI21X1_309/B gnd NOR2X1_194/A vdd OAI21X1
XINVX1_124 INVX1_124/A gnd INVX1_124/Y vdd INVX1
XNAND2X1_417 NAND3X1_355/Y AOI22X1_12/C gnd NAND2X1_417/Y vdd NAND2X1
XNOR2X1_336 gnd NOR2X1_336/B gnd NOR2X1_336/Y vdd NOR2X1
XAND2X2_28 gnd OR2X2_35/B gnd AND2X2_28/Y vdd AND2X2
XNAND3X1_249 NAND3X1_251/A NAND3X1_249/B NAND3X1_249/C gnd AND2X2_84/A vdd NAND3X1
XBUFX2_250 XOR2X1_30/Y gnd BUFX2_250/Y vdd BUFX2
XBUFX4_13 INVX8_2/Y gnd BUFX4_13/Y vdd BUFX4
XINVX2_88 INVX2_88/A gnd INVX2_88/Y vdd INVX2
XOAI21X1_267 OAI21X1_267/A XNOR2X1_142/B INVX1_184/A gnd XOR2X1_160/A vdd OAI21X1
XNOR2X1_300 gnd NOR2X1_300/B gnd NOR2X1_300/Y vdd NOR2X1
XNAND2X1_381 INVX1_244/Y AND2X2_110/A gnd NAND2X1_382/B vdd NAND2X1
XNAND3X1_213 NAND3X1_213/A NAND3X1_213/B AOI21X1_146/Y gnd AND2X2_72/A vdd NAND3X1
XFILL_25_9_1 gnd vdd FILL
XFILL_27_7_0 gnd vdd FILL
XBUFX2_214 BUFX2_214/A gnd BUFX2_214/Y vdd BUFX2
XXNOR2X1_252 XNOR2X1_252/A INVX2_92/Y gnd XOR2X1_2/A vdd XNOR2X1
XNOR2X1_67 NOR2X1_67/A NOR2X1_66/Y gnd XOR2X1_58/A vdd NOR2X1
XFILL_7_8_0 gnd vdd FILL
XOAI21X1_231 NOR3X1_52/C NOR3X1_52/B INVX1_155/Y gnd NAND3X1_242/A vdd OAI21X1
XNAND2X1_345 INVX1_207/Y AND2X2_103/A gnd NAND3X1_306/C vdd NAND2X1
XINVX2_52 INVX2_52/A gnd INVX2_52/Y vdd INVX2
XNOR2X1_264 gnd NOR2X1_264/B gnd NOR2X1_264/Y vdd NOR2X1
XNOR2X1_31 NOR2X1_31/A INVX2_15/A gnd XOR2X1_20/B vdd NOR2X1
XINVX1_593 INVX1_593/A gnd INVX1_593/Y vdd INVX1
XBUFX2_178 BUFX2_178/A gnd BUFX2_178/Y vdd BUFX2
XXNOR2X1_216 bloque_bytes[42] bloque_bytes[2] gnd XNOR2X1_216/Y vdd XNOR2X1
XNAND3X1_177 NAND3X1_179/A NAND3X1_177/B NAND3X1_177/C gnd AND2X2_60/A vdd NAND3X1
XFILL_35_4_1 gnd vdd FILL
XOAI21X1_195 NOR3X1_47/C NOR3X1_47/B INVX1_132/Y gnd NAND2X1_231/A vdd OAI21X1
XINVX2_16 INVX2_16/A gnd INVX2_16/Y vdd INVX2
XNAND2X1_309 NAND3X1_278/Y NAND2X1_309/B gnd XNOR2X1_142/A vdd NAND2X1
XNOR2X1_228 gnd NOR2X1_228/B gnd NOR2X1_228/Y vdd NOR2X1
XINVX1_557 bloque_bytes[0] gnd INVX1_557/Y vdd INVX1
XNAND3X1_141 OAI21X1_135/Y NAND3X1_140/Y AOI21X1_98/Y gnd AND2X2_48/A vdd NAND3X1
XCLKBUF1_19 BUFX4_4/Y gnd CLKBUF1_19/Y vdd CLKBUF1
XBUFX2_142 gnd gnd BUFX2_142/Y vdd BUFX2
XXNOR2X1_180 NOR2X1_278/A XNOR2X1_180/B gnd BUFX2_222/A vdd XNOR2X1
XOAI21X1_159 OAI21X1_159/A OAI21X1_158/Y INVX1_106/Y gnd NAND3X1_166/C vdd OAI21X1
XFILL_11_0_0 gnd vdd FILL
XNOR2X1_192 gnd NOR2X1_192/B gnd NOR2X1_192/Y vdd NOR2X1
XNAND2X1_273 gnd AND2X2_82/B gnd NAND3X1_245/B vdd NAND2X1
XNOR3X1_72 NOR3X1_72/A INVX2_66/Y NOR3X1_72/C gnd NOR3X1_72/Y vdd NOR3X1
XINVX1_521 bloque_bytes[61] gnd INVX1_521/Y vdd INVX1
XNAND3X1_105 NAND3X1_107/A NAND3X1_104/Y AOI21X1_74/Y gnd AND2X2_36/A vdd NAND3X1
XDFFPOSX1_339 INVX1_397/A CLKBUF1_8/Y NAND2X1_684/Y gnd vdd DFFPOSX1
XBUFX2_106 gnd gnd BUFX2_106/Y vdd BUFX2
XOAI21X1_123 XNOR2X1_62/A AOI21X1_94/C NOR2X1_85/Y gnd NOR2X1_86/B vdd OAI21X1
XXNOR2X1_66 XNOR2X1_66/A OR2X2_55/Y gnd INVX1_87/A vdd XNOR2X1
XXNOR2X1_144 XNOR2X1_144/A INVX2_58/Y gnd XOR2X1_167/A vdd XNOR2X1
XFILL_34_7_0 gnd vdd FILL
XNOR2X1_156 INVX1_161/Y NOR2X1_156/B gnd NOR2X1_156/Y vdd NOR2X1
XNAND2X1_237 INVX2_45/Y OAI21X1_204/Y gnd NAND2X1_237/Y vdd NAND2X1
XFILL_32_9_1 gnd vdd FILL
XNOR3X1_36 INVX1_67/Y NOR3X1_36/B NOR3X1_36/C gnd NOR2X1_73/B vdd NOR3X1
XDFFPOSX1_303 INVX1_311/A CLKBUF1_34/Y INVX1_552/Y gnd vdd DFFPOSX1
XINVX1_485 INVX1_485/A gnd NOR3X1_95/A vdd INVX1
XXOR2X1_300 bloque_bytes[43] bloque_bytes[3] gnd XOR2X1_300/Y vdd XOR2X1
XXNOR2X1_108 XNOR2X1_108/A INVX2_46/Y gnd XOR2X1_127/A vdd XNOR2X1
XXNOR2X1_30 XNOR2X1_30/A OR2X2_23/Y gnd INVX1_43/A vdd XNOR2X1
XNOR2X1_120 gnd OR2X2_83/B gnd NOR2X1_120/Y vdd NOR2X1
XNAND2X1_201 OR2X2_77/A OR2X2_77/B gnd NAND2X1_201/Y vdd NAND2X1
XFILL_4_1 gnd vdd FILL
XOR2X2_88 OR2X2_88/A OR2X2_88/B gnd OR2X2_88/Y vdd OR2X2
XOAI21X1_628 NOR2X1_433/Y OAI21X1_628/B INVX1_570/A gnd OAI21X1_628/Y vdd OAI21X1
XDFFPOSX1_267 INVX1_226/A CLKBUF1_32/Y XNOR2X1_236/A gnd vdd DFFPOSX1
XAOI21X1_99 NOR3X1_39/Y NOR2X1_93/Y NOR2X1_91/A gnd AOI21X1_99/Y vdd AOI21X1
XINVX1_449 INVX1_449/A gnd INVX1_449/Y vdd INVX1
XXOR2X1_264 BUFX2_230/A gnd gnd NOR2X1_327/B vdd XOR2X1
XAOI21X1_401 OR2X2_160/B OR2X2_160/A AND2X2_197/B gnd NOR2X1_452/A vdd AOI21X1
XXOR2X1_4 XOR2X1_4/A gnd gnd AND2X2_9/B vdd XOR2X1
XNAND2X1_165 OAI21X1_139/Y OR2X2_64/B gnd OR2X2_62/A vdd NAND2X1
XFILL_18_0_0 gnd vdd FILL
XDFFPOSX1_231 INVX1_158/A CLKBUF1_36/Y INVX1_574/A gnd vdd DFFPOSX1
XMUX2X1_10 BUFX2_10/A INVX1_3/A MUX2X1_9/S gnd NOR3X1_10/B vdd MUX2X1
XOR2X2_52 OR2X2_52/A OR2X2_52/B gnd OR2X2_52/Y vdd OR2X2
XAOI21X1_63 NOR3X1_33/Y NOR2X1_63/Y NOR2X1_61/A gnd OAI21X1_85/C vdd AOI21X1
XOAI21X1_592 bloque_bytes[67] INVX1_496/Y OAI21X1_592/C gnd NOR2X1_412/B vdd OAI21X1
XFILL_16_2_1 gnd vdd FILL
XINVX1_413 INVX1_413/A gnd INVX1_413/Y vdd INVX1
XNAND2X1_706 NAND3X1_533/B NAND3X1_533/A gnd XNOR2X1_253/A vdd NAND2X1
XBUFX2_66 gnd gnd BUFX2_66/Y vdd BUFX2
XXOR2X1_228 BUFX2_214/A gnd gnd NOR2X1_279/B vdd XOR2X1
XNAND3X1_538 INVX1_592/Y NAND3X1_537/B OR2X2_157/Y gnd AOI21X1_396/B vdd NAND3X1
XNAND2X1_129 NAND2X1_129/A OR2X2_47/Y gnd OR2X2_48/A vdd NAND2X1
XAOI21X1_365 INVX1_515/Y bloque_bytes[19] AOI21X1_365/C gnd INVX1_517/A vdd AOI21X1
XOR2X2_16 OR2X2_16/A OR2X2_16/B gnd INVX1_31/A vdd OR2X2
XAOI21X1_27 NOR3X1_27/Y NOR2X1_33/Y NOR2X1_31/A gnd OAI21X1_34/C vdd AOI21X1
XDFFPOSX1_195 INVX1_110/A CLKBUF1_10/Y bloque_bytes[9] gnd vdd DFFPOSX1
XDFFPOSX1_7 BUFX2_6/A CLKBUF1_4/Y NOR3X1_6/Y gnd vdd DFFPOSX1
XINVX1_377 INVX1_377/A gnd INVX1_377/Y vdd INVX1
XNAND2X1_670 XNOR2X1_234/Y INVX1_546/A gnd NAND2X1_670/Y vdd NAND2X1
XXOR2X1_192 BUFX2_194/A gnd gnd XOR2X1_192/Y vdd XOR2X1
XOAI21X1_556 NOR3X1_85/C OAI21X1_556/B INVX1_465/A gnd NOR2X1_353/A vdd OAI21X1
XBUFX2_30 gnd gnd BUFX2_30/Y vdd BUFX2
XNAND2X1_90 OR2X2_31/B OR2X2_31/A gnd NAND2X1_91/A vdd NAND2X1
XOAI21X1_75 NOR2X1_57/A INVX1_53/Y INVX1_54/Y gnd NAND2X1_95/B vdd OAI21X1
XNAND3X1_502 INVX2_80/A NOR2X1_406/Y NOR3X1_90/Y gnd AOI21X1_348/B vdd NAND3X1
XAOI21X1_329 INVX1_476/Y NAND2X1_616/Y OAI21X1_574/Y gnd AOI21X1_329/Y vdd AOI21X1
XINVX2_3 target[4] gnd INVX2_3/Y vdd INVX2
XDFFPOSX1_93 MUX2X1_4/B CLKBUF1_4/Y NAND2X1_700/Y gnd vdd DFFPOSX1
XDFFPOSX1_159 INVX1_59/A CLKBUF1_7/Y bloque_bytes[53] gnd vdd DFFPOSX1
XINVX1_341 INVX1_341/A gnd INVX1_341/Y vdd INVX1
XOAI21X1_520 BUFX2_228/A NOR2X1_330/B INVX1_425/Y gnd NAND3X1_456/B vdd OAI21X1
XNAND2X1_634 INVX1_483/A INVX1_484/A gnd NOR2X1_406/A vdd NAND2X1
XXOR2X1_156 XOR2X1_156/A BUFX2_171/A gnd INVX1_195/A vdd XOR2X1
XBUFX2_8 BUFX2_8/A gnd hash[7] vdd BUFX2
XNAND2X1_54 OR2X2_16/B OR2X2_16/A gnd NAND2X1_55/A vdd NAND2X1
XFILL_13_7_1 gnd vdd FILL
XFILL_15_5_0 gnd vdd FILL
XAOI21X1_293 INVX1_402/A NAND3X1_439/B INVX1_401/Y gnd NOR3X1_79/C vdd AOI21X1
XNAND3X1_466 INVX1_441/Y INVX1_442/Y INVX1_443/Y gnd NAND3X1_466/Y vdd NAND3X1
XOAI21X1_39 INVX2_16/Y AND2X2_12/B INVX1_27/A gnd OAI21X1_39/Y vdd OAI21X1
XDFFPOSX1_123 INVX1_11/A CLKBUF1_16/Y bloque_bytes[81] gnd vdd DFFPOSX1
XDFFPOSX1_57 OR2X2_144/B CLKBUF1_6/Y NOR2X1_379/Y gnd vdd DFFPOSX1
XXOR2X1_120 XOR2X1_120/A XOR2X1_120/B gnd BUFX2_166/A vdd XOR2X1
XINVX1_305 INVX1_305/A gnd INVX1_305/Y vdd INVX1
XOAI21X1_484 gnd NOR2X1_300/B INVX1_379/Y gnd OAI21X1_484/Y vdd OAI21X1
XFILL_25_0_0 gnd vdd FILL
XNOR2X1_1 target[7] NOR2X1_1/B gnd INVX1_2/A vdd NOR2X1
XNAND2X1_598 INVX1_463/A NOR2X1_354/Y gnd NAND2X1_598/Y vdd NAND2X1
XFILL_3_3_1 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XFILL_23_2_1 gnd vdd FILL
XNAND2X1_18 OAI21X1_7/Y NOR2X1_11/Y gnd AOI21X1_9/A vdd NAND2X1
XNAND3X1_430 INVX1_388/A OAI21X1_482/Y NAND3X1_430/C gnd NAND2X1_524/A vdd NAND3X1
XAOI21X1_257 AOI21X1_257/A AOI21X1_257/B NAND2X1_455/Y gnd AOI21X1_257/Y vdd AOI21X1
XINVX1_269 INVX1_269/A gnd INVX1_269/Y vdd INVX1
XOAI21X1_448 OAI21X1_448/A INVX1_356/A INVX1_355/Y gnd AND2X2_133/A vdd OAI21X1
XDFFPOSX1_21 BUFX2_20/A CLKBUF1_42/Y NOR3X1_20/Y gnd vdd DFFPOSX1
XNAND3X1_95 INVX1_66/A NAND3X1_95/B OR2X2_41/Y gnd NAND3X1_96/A vdd NAND3X1
XXOR2X1_64 XOR2X1_78/B gnd gnd OR2X2_58/B vdd XOR2X1
XNAND2X1_562 NAND2X1_562/A NAND2X1_562/B gnd XOR2X1_278/B vdd NAND2X1
XAOI21X1_221 INVX1_231/A NAND3X1_322/B INVX1_230/Y gnd NOR3X1_61/C vdd AOI21X1
XOR2X2_147 OR2X2_137/Y INVX1_503/A gnd OR2X2_147/Y vdd OR2X2
XNAND3X1_394 INVX1_326/A NAND3X1_394/B NAND3X1_389/Y gnd NAND2X1_474/A vdd NAND3X1
XAND2X2_164 INVX8_2/A AND2X2_164/B gnd AND2X2_164/Y vdd AND2X2
XINVX1_233 INVX1_233/A gnd INVX1_233/Y vdd INVX1
XOAI21X1_412 OAI21X1_412/A INVX1_316/A INVX1_319/A gnd OAI21X1_412/Y vdd OAI21X1
XXOR2X1_28 XOR2X1_28/A XOR2X1_28/B gnd XOR2X1_28/Y vdd XOR2X1
XNAND3X1_59 INVX1_44/A NAND3X1_59/B OR2X2_25/Y gnd OAI21X1_62/C vdd NAND3X1
XNOR2X1_445 gnd gnd gnd NOR3X1_97/B vdd NOR2X1
XOR2X2_111 OR2X2_111/A INVX1_160/Y gnd OR2X2_111/Y vdd OR2X2
XNAND2X1_526 XOR2X1_260/B NOR2X1_304/Y gnd AOI21X1_288/C vdd NAND2X1
XAOI21X1_185 AOI21X1_185/A AOI21X1_185/B OAI21X1_256/B gnd NAND3X1_272/B vdd AOI21X1
XNAND3X1_358 INVX2_64/A NAND3X1_358/B NAND3X1_358/C gnd NOR3X1_67/A vdd NAND3X1
XNAND2X1_7 NOR2X1_2/Y NAND2X1_7/B gnd AOI21X1_5/B vdd NAND2X1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XFILL_22_5_0 gnd vdd FILL
XOAI22X1_6 INVX2_8/Y INVX1_5/A INVX1_6/A INVX2_9/Y gnd OAI22X1_6/Y vdd OAI22X1
XNAND3X1_23 INVX1_22/A NAND2X1_40/Y OR2X2_9/Y gnd NAND2X1_41/B vdd NAND3X1
XFILL_2_6_0 gnd vdd FILL
XNOR2X1_409 INVX1_549/A OR2X2_140/A gnd INVX1_534/A vdd NOR2X1
XINVX1_197 INVX1_197/A gnd INVX1_197/Y vdd INVX1
XFILL_20_7_1 gnd vdd FILL
XOAI21X1_376 gnd NOR2X1_239/B INVX1_283/A gnd INVX2_64/A vdd OAI21X1
XAND2X2_128 AND2X2_128/A NOR3X1_71/A gnd BUFX2_216/A vdd AND2X2
XFILL_0_8_1 gnd vdd FILL
XNAND2X1_490 OAI21X1_447/Y NAND2X1_490/B gnd NOR2X1_284/B vdd NAND2X1
XNAND3X1_322 INVX1_231/A NAND3X1_322/B INVX1_230/Y gnd INVX1_237/A vdd NAND3X1
XAOI21X1_149 AOI21X1_149/A AOI21X1_149/B OAI21X1_205/B gnd NAND3X1_218/B vdd AOI21X1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XOAI21X1_340 gnd XOR2X1_182/Y INVX1_246/A gnd INVX1_249/A vdd OAI21X1
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XFILL_32_0_0 gnd vdd FILL
XFILL_30_2_1 gnd vdd FILL
XNOR2X1_373 BUFX4_15/Y INVX2_78/Y gnd NOR2X1_373/Y vdd NOR2X1
XNAND2X1_454 NAND2X1_454/A INVX1_316/Y gnd INVX1_317/A vdd NAND2X1
XAOI21X1_113 NAND3X1_161/Y NAND3X1_163/Y AOI21X1_113/C gnd NAND3X1_164/B vdd AOI21X1
XAND2X2_65 OR2X2_84/A OR2X2_84/B gnd AND2X2_65/Y vdd AND2X2
XNAND3X1_286 INVX1_180/Y NAND3X1_286/B OR2X2_125/Y gnd NAND3X1_287/C vdd NAND3X1
XINVX1_125 INVX1_125/A gnd INVX1_125/Y vdd INVX1
XOAI21X1_304 NOR3X1_60/A NOR3X1_60/C INVX2_60/A gnd NOR2X1_193/A vdd OAI21X1
XNOR2X1_337 NOR2X1_337/A INVX1_437/Y gnd NOR2X1_337/Y vdd NOR2X1
XNAND2X1_418 OAI21X1_374/Y NAND2X1_418/B gnd XOR2X1_214/A vdd NAND2X1
XAND2X2_29 OR2X2_36/A OR2X2_36/B gnd AND2X2_29/Y vdd AND2X2
XBUFX2_251 OR2X2_44/A gnd BUFX2_251/Y vdd BUFX2
XNAND3X1_250 INVX1_158/Y NAND3X1_252/B OR2X2_109/Y gnd NAND3X1_251/C vdd NAND3X1
XBUFX4_14 INVX8_2/Y gnd BUFX4_14/Y vdd BUFX4
XINVX2_89 INVX2_89/A gnd INVX2_89/Y vdd INVX2
XFILL_17_1 gnd vdd FILL
XOAI21X1_268 AND2X2_94/Y NOR2X1_170/Y INVX1_178/Y gnd AOI21X1_192/A vdd OAI21X1
XNAND2X1_382 OAI21X1_337/Y NAND2X1_382/B gnd INVX1_289/A vdd NAND2X1
XNOR2X1_301 NOR2X1_301/A INVX1_380/Y gnd NOR2X1_301/Y vdd NOR2X1
XFILL_27_7_1 gnd vdd FILL
XFILL_29_5_0 gnd vdd FILL
XFILL_7_8_1 gnd vdd FILL
XFILL_9_6_0 gnd vdd FILL
XNAND3X1_214 INVX1_136/Y NAND2X1_239/Y OR2X2_93/Y gnd NAND3X1_214/Y vdd NAND3X1
XBUFX2_215 BUFX2_215/A gnd BUFX2_215/Y vdd BUFX2
XXNOR2X1_253 XNOR2X1_253/A NAND2X1_704/Y gnd XOR2X1_3/A vdd XNOR2X1
XNOR2X1_68 gnd OR2X2_41/B gnd NOR3X1_35/B vdd NOR2X1
XOAI21X1_232 NOR3X1_52/Y NOR2X1_153/A NAND2X1_269/B gnd NAND2X1_272/B vdd OAI21X1
XINVX2_53 INVX2_53/A gnd INVX2_53/Y vdd INVX2
XNAND2X1_346 INVX1_208/Y NOR2X1_192/Y gnd NAND2X1_347/B vdd NAND2X1
XNOR2X1_265 NOR2X1_265/A INVX1_323/Y gnd NOR2X1_265/Y vdd NOR2X1
XNAND3X1_178 INVX1_114/Y NAND2X1_201/Y OR2X2_77/Y gnd NAND3X1_178/Y vdd NAND3X1
XINVX1_594 INVX1_594/A gnd INVX1_594/Y vdd INVX1
XNOR2X1_32 XOR2X1_2/A OR2X2_12/B gnd NOR2X1_32/Y vdd NOR2X1
XXNOR2X1_217 bloque_bytes[47] bloque_bytes[7] gnd XNOR2X1_217/Y vdd XNOR2X1
XBUFX2_179 BUFX2_179/A gnd BUFX2_179/Y vdd BUFX2
XINVX2_17 INVX2_17/A gnd INVX2_17/Y vdd INVX2
XOAI21X1_196 NOR3X1_48/Y NOR2X1_133/A NOR3X1_47/Y gnd NAND2X1_233/B vdd OAI21X1
XNOR2X1_229 NOR2X1_229/A INVX1_266/Y gnd NOR2X1_230/B vdd NOR2X1
XNAND2X1_310 INVX1_184/A NAND2X1_310/B gnd OAI21X1_267/A vdd NAND2X1
XCLKBUF1_20 BUFX4_6/Y gnd CLKBUF1_20/Y vdd CLKBUF1
XNAND3X1_142 INVX1_92/Y NAND2X1_163/Y OR2X2_61/Y gnd NAND3X1_142/Y vdd NAND3X1
XINVX1_558 INVX1_558/A gnd INVX1_558/Y vdd INVX1
XBUFX2_143 gnd gnd BUFX2_143/Y vdd BUFX2
XOAI21X1_160 NOR2X1_107/A INVX1_108/Y INVX1_109/Y gnd OAI21X1_160/Y vdd OAI21X1
XXNOR2X1_181 NOR2X1_281/Y NOR2X1_280/Y gnd XOR2X1_247/A vdd XNOR2X1
XFILL_11_0_1 gnd vdd FILL
XNOR2X1_193 NOR2X1_193/A INVX1_209/Y gnd NOR2X1_194/B vdd NOR2X1
XNAND2X1_274 OR2X2_108/A OR2X2_108/B gnd NAND3X1_248/B vdd NAND2X1
XDFFPOSX1_340 INVX1_398/A CLKBUF1_45/Y NAND2X1_685/Y gnd vdd DFFPOSX1
XNOR3X1_73 NOR3X1_73/A INVX1_342/A NOR3X1_73/C gnd NOR3X1_73/Y vdd NOR3X1
XNAND3X1_106 INVX1_70/Y NAND3X1_106/B OR2X2_45/Y gnd NAND3X1_107/C vdd NAND3X1
XINVX1_522 INVX1_522/A gnd INVX1_522/Y vdd INVX1
XXNOR2X1_145 BUFX2_173/A XOR2X1_148/Y gnd OR2X2_127/A vdd XNOR2X1
XBUFX2_107 gnd gnd BUFX2_107/Y vdd BUFX2
XFILL_36_5_0 gnd vdd FILL
XOAI21X1_124 INVX2_31/Y AND2X2_42/B INVX1_82/A gnd OAI21X1_125/B vdd OAI21X1
XXNOR2X1_67 gnd XOR2X1_62/Y gnd XNOR2X1_67/Y vdd XNOR2X1
XFILL_34_7_1 gnd vdd FILL
XNOR2X1_157 NOR2X1_157/A NOR2X1_156/Y gnd XOR2X1_148/A vdd NOR2X1
XNAND2X1_238 AND2X2_72/B AND2X2_72/A gnd OAI21X1_205/B vdd NAND2X1
XNOR3X1_37 INVX1_77/Y NOR3X1_37/B NOR3X1_37/C gnd NOR3X1_37/Y vdd NOR3X1
XINVX1_486 MUX2X1_3/S gnd INVX1_486/Y vdd INVX1
XDFFPOSX1_304 INVX1_315/A CLKBUF1_17/Y INVX1_553/Y gnd vdd DFFPOSX1
XXOR2X1_301 bloque_bytes[44] bloque_bytes[4] gnd NOR2X1_413/A vdd XOR2X1
XXNOR2X1_109 BUFX2_157/A XOR2X1_108/Y gnd OR2X2_95/A vdd XNOR2X1
XXNOR2X1_31 gnd XOR2X1_22/Y gnd AOI21X1_57/B vdd XNOR2X1
XNOR2X1_121 NOR2X1_121/A INVX2_42/A gnd XOR2X1_110/B vdd NOR2X1
XFILL_10_3_0 gnd vdd FILL
XNAND2X1_202 NAND3X1_179/Y NAND3X1_181/Y gnd INVX2_40/A vdd NAND2X1
XFILL_4_2 gnd vdd FILL
XOAI21X1_629 AOI21X1_393/Y NOR2X1_434/Y INVX1_573/A gnd OAI21X1_629/Y vdd OAI21X1
XOR2X2_89 gnd OR2X2_89/B gnd OR2X2_89/Y vdd OR2X2
XDFFPOSX1_268 INVX1_227/A CLKBUF1_27/Y NAND2X1_652/Y gnd vdd DFFPOSX1
XINVX1_450 INVX1_450/A gnd INVX1_450/Y vdd INVX1
XXOR2X1_265 XOR2X1_265/A BUFX2_223/A gnd INVX1_423/A vdd XOR2X1
XAOI21X1_402 NOR2X1_452/Y AOI21X1_402/B INVX1_597/A gnd NOR2X1_454/A vdd AOI21X1
XXOR2X1_5 XOR2X1_5/A gnd gnd OR2X2_11/B vdd XOR2X1
XNAND2X1_166 OR2X2_63/B OR2X2_63/A gnd NAND2X1_166/Y vdd NAND2X1
XAOI21X1_64 NAND3X1_84/B OR2X2_36/Y INVX1_58/A gnd OR2X2_38/B vdd AOI21X1
XDFFPOSX1_232 INVX1_160/A CLKBUF1_14/Y INVX1_575/A gnd vdd DFFPOSX1
XFILL_18_0_1 gnd vdd FILL
XMUX2X1_11 BUFX2_11/A NOR2X1_5/A BUFX4_9/Y gnd NOR3X1_11/B vdd MUX2X1
XOR2X2_53 OR2X2_53/A OR2X2_53/B gnd OR2X2_53/Y vdd OR2X2
XOAI21X1_593 bloque_bytes[68] INVX1_497/Y OAI21X1_593/C gnd NOR2X1_413/B vdd OAI21X1
XXOR2X1_229 XOR2X1_229/A BUFX2_207/A gnd INVX1_347/A vdd XOR2X1
XINVX1_414 INVX1_414/A gnd INVX1_414/Y vdd INVX1
XNAND2X1_707 gnd gnd gnd AOI21X1_394/A vdd NAND2X1
XBUFX2_67 gnd gnd BUFX2_67/Y vdd BUFX2
XNAND3X1_539 INVX1_593/Y NAND3X1_541/B OR2X2_158/Y gnd NAND3X1_539/Y vdd NAND3X1
XNAND2X1_130 OR2X2_48/B OR2X2_48/A gnd NAND2X1_130/Y vdd NAND2X1
XAOI21X1_366 INVX1_518/Y bloque_bytes[20] AOI21X1_366/C gnd INVX1_520/A vdd AOI21X1
XOR2X2_17 gnd OR2X2_17/B gnd OR2X2_17/Y vdd OR2X2
XAOI21X1_28 NAND3X1_30/B OR2X2_12/Y INVX1_25/A gnd OR2X2_14/B vdd AOI21X1
XDFFPOSX1_8 BUFX2_7/A CLKBUF1_43/Y NOR3X1_7/Y gnd vdd DFFPOSX1
XINVX1_378 INVX1_378/A gnd INVX1_378/Y vdd INVX1
XOAI21X1_557 NOR2X1_353/Y NOR2X1_352/B AOI22X1_22/C gnd XOR2X1_296/A vdd OAI21X1
XDFFPOSX1_196 INVX1_111/A CLKBUF1_10/Y bloque_bytes[10] gnd vdd DFFPOSX1
XBUFX2_31 gnd gnd BUFX2_31/Y vdd BUFX2
XNAND2X1_671 bloque_bytes[6] OR2X2_140/A gnd AOI21X1_384/A vdd NAND2X1
XXOR2X1_193 XOR2X1_193/A INVX1_251/A gnd INVX1_271/A vdd XOR2X1
XAOI21X1_330 AND2X2_162/B NOR2X1_389/Y AOI21X1_330/C gnd AOI21X1_330/Y vdd AOI21X1
XNAND2X1_91 NAND2X1_91/A OR2X2_31/Y gnd OR2X2_32/A vdd NAND2X1
XDFFPOSX1_160 INVX1_61/A CLKBUF1_7/Y bloque_bytes[54] gnd vdd DFFPOSX1
XOAI21X1_76 AND2X2_26/Y NOR2X1_58/Y INVX1_55/Y gnd OAI21X1_76/Y vdd OAI21X1
XNAND3X1_503 XNOR2X1_208/Y NAND3X1_503/B AOI21X1_370/Y gnd AOI21X1_379/C vdd NAND3X1
XDFFPOSX1_94 MUX2X1_5/B CLKBUF1_35/Y NAND2X1_701/Y gnd vdd DFFPOSX1
XINVX2_4 target[1] gnd INVX2_4/Y vdd INVX2
XINVX1_342 INVX1_342/A gnd INVX1_342/Y vdd INVX1
XOAI21X1_521 BUFX2_228/A NOR2X1_330/B INVX1_425/A gnd AOI22X1_20/B vdd OAI21X1
XBUFX2_9 BUFX2_9/A gnd hash[8] vdd BUFX2
XNAND2X1_635 BUFX4_30/Y NAND3X1_501/Y gnd NAND2X1_635/Y vdd NAND2X1
XXOR2X1_157 XOR2X1_157/A OR2X2_125/A gnd NOR2X1_186/B vdd XOR2X1
XFILL_17_3_0 gnd vdd FILL
XNAND2X1_55 NAND2X1_55/A INVX1_31/A gnd INVX1_29/A vdd NAND2X1
XFILL_15_5_1 gnd vdd FILL
XAOI21X1_294 OAI21X1_503/Y AOI21X1_294/B INVX2_70/A gnd AOI21X1_294/Y vdd AOI21X1
XNAND3X1_467 INVX1_443/A INVX1_441/Y INVX1_442/Y gnd NAND3X1_467/Y vdd NAND3X1
XDFFPOSX1_124 INVX1_12/A CLKBUF1_5/Y bloque_bytes[82] gnd vdd DFFPOSX1
XOAI21X1_40 AOI21X1_34/Y OAI21X1_39/Y INVX1_29/Y gnd OAI21X1_40/Y vdd OAI21X1
XDFFPOSX1_58 INVX1_472/A CLKBUF1_15/Y NOR2X1_382/Y gnd vdd DFFPOSX1
XXOR2X1_121 BUFX2_158/A XOR2X1_121/B gnd XOR2X1_121/Y vdd XOR2X1
XINVX1_306 INVX1_306/A gnd INVX1_306/Y vdd INVX1
XOAI21X1_485 BUFX2_221/A XOR2X1_249/Y INVX1_391/A gnd XNOR2X1_191/B vdd OAI21X1
XFILL_25_0_1 gnd vdd FILL
XNOR2X1_2 NOR2X1_2/A NOR2X1_2/B gnd NOR2X1_2/Y vdd NOR2X1
XNAND2X1_599 INVX1_463/Y NOR2X1_354/Y gnd INVX1_466/A vdd NAND2X1
XFILL_5_1_1 gnd vdd FILL
XDFFPOSX1_22 BUFX2_21/A CLKBUF1_43/Y NOR3X1_21/Y gnd vdd DFFPOSX1
XNAND2X1_19 NOR2X1_13/Y NOR2X1_14/Y gnd NOR2X1_16/A vdd NAND2X1
XNAND3X1_431 AOI22X1_18/B INVX1_390/A INVX1_388/Y gnd NAND2X1_524/B vdd NAND3X1
XAOI21X1_258 INVX1_318/Y NAND3X1_382/C INVX1_317/A gnd OAI21X1_412/A vdd AOI21X1
XINVX1_270 BUFX2_191/A gnd INVX1_270/Y vdd INVX1
XOAI21X1_449 NOR2X1_281/A NOR3X1_73/Y AOI21X1_273/Y gnd OAI21X1_449/Y vdd OAI21X1
XNAND3X1_96 NAND3X1_96/A OAI21X1_93/Y NAND3X1_96/C gnd XNOR2X1_52/B vdd NAND3X1
XXOR2X1_65 BUFX2_262/A gnd gnd OR2X2_59/B vdd XOR2X1
XOR2X2_148 OR2X2_138/Y INVX1_504/A gnd OR2X2_148/Y vdd OR2X2
XNAND2X1_563 INVX1_417/A NOR2X1_324/Y gnd NAND2X1_563/Y vdd NAND2X1
XAOI21X1_222 AOI21X1_222/A NAND2X1_373/Y INVX2_61/A gnd AOI21X1_223/B vdd AOI21X1
XFILL_14_8_0 gnd vdd FILL
XNAND3X1_395 INVX1_337/Y INVX1_336/A AOI21X1_266/B gnd AND2X2_129/B vdd NAND3X1
XXOR2X1_29 XOR2X1_29/A XOR2X1_15/A gnd XOR2X1_29/Y vdd XOR2X1
XNOR2X1_446 gnd gnd gnd NOR3X1_98/B vdd NOR2X1
XINVX1_234 INVX1_234/A gnd INVX1_234/Y vdd INVX1
XAND2X2_165 BUFX4_31/Y AND2X2_165/B gnd AND2X2_165/Y vdd AND2X2
XOAI21X1_413 gnd NOR2X1_262/B INVX1_320/A gnd NAND2X1_458/A vdd OAI21X1
XNAND3X1_60 OAI21X1_62/C NAND3X1_60/B NAND3X1_60/C gnd OAI21X1_68/B vdd NAND3X1
XOR2X2_112 OR2X2_112/A OR2X2_112/B gnd INVX1_163/A vdd OR2X2
XNAND2X1_527 INVX1_391/Y NOR2X1_307/Y gnd NAND2X1_528/B vdd NAND2X1
XAOI21X1_186 OR2X2_118/B OR2X2_118/A AND2X2_90/B gnd NOR2X1_165/A vdd AOI21X1
XNAND3X1_359 INVX1_287/A NAND2X1_423/B INVX2_64/Y gnd OAI21X1_385/B vdd NAND3X1
XNAND2X1_8 target[5] INVX2_1/Y gnd OAI21X1_3/C vdd NAND2X1
XFILL_4_4_0 gnd vdd FILL
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XINVX1_198 AOI22X1_8/D gnd INVX1_198/Y vdd INVX1
XFILL_22_5_1 gnd vdd FILL
XFILL_24_3_0 gnd vdd FILL
XOAI21X1_377 NOR3X1_68/C INVX2_64/Y NOR3X1_68/A gnd AND2X2_120/A vdd OAI21X1
XOAI22X1_7 INVX1_5/Y target[7] INVX1_6/Y target[6] gnd NOR2X1_13/B vdd OAI22X1
XNAND3X1_24 NAND2X1_41/B NAND2X1_41/A NAND3X1_24/C gnd XNOR2X1_16/B vdd NAND3X1
XFILL_2_6_1 gnd vdd FILL
XNOR2X1_410 NOR2X1_410/A NOR2X1_410/B gnd NOR2X1_410/Y vdd NOR2X1
XAND2X2_129 AND2X2_129/A AND2X2_129/B gnd XOR2X1_240/A vdd AND2X2
XNAND2X1_491 INVX1_352/Y NOR2X1_284/B gnd NAND2X1_491/Y vdd NAND2X1
XAOI21X1_150 OR2X2_94/B OR2X2_94/A AND2X2_72/B gnd NOR2X1_135/A vdd AOI21X1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XNAND3X1_323 INVX1_232/Y INVX1_233/Y INVX1_234/Y gnd NAND3X1_323/Y vdd NAND3X1
XFILL_32_0_1 gnd vdd FILL
XOAI21X1_341 NOR3X1_63/A INVX1_247/A OAI21X1_347/B gnd NOR2X1_218/A vdd OAI21X1
XINVX1_162 INVX1_162/A gnd INVX1_162/Y vdd INVX1
XNOR2X1_374 BUFX4_15/Y INVX2_79/Y gnd NOR2X1_374/Y vdd NOR2X1
XNAND2X1_455 NAND3X1_381/Y AOI22X1_14/C gnd NAND2X1_455/Y vdd NAND2X1
XAOI21X1_114 OR2X2_70/B OR2X2_70/A AND2X2_54/B gnd NOR2X1_105/A vdd AOI21X1
XNAND3X1_287 NAND3X1_287/A NAND3X1_287/B NAND3X1_287/C gnd AOI21X1_197/A vdd NAND3X1
XAND2X2_66 AND2X2_66/A AND2X2_66/B gnd AND2X2_66/Y vdd AND2X2
XINVX1_126 OR2X2_86/Y gnd INVX1_126/Y vdd INVX1
XOAI21X1_305 gnd XOR2X1_165/Y INVX1_210/Y gnd NAND3X1_308/B vdd OAI21X1
XNOR2X1_338 NOR2X1_338/A NOR2X1_337/Y gnd BUFX2_245/A vdd NOR2X1
XFILL_21_8_0 gnd vdd FILL
XNAND2X1_419 INVX1_282/Y NOR2X1_238/Y gnd NAND3X1_358/B vdd NAND2X1
XFILL_1_9_0 gnd vdd FILL
XBUFX2_252 OR2X2_45/A gnd BUFX2_252/Y vdd BUFX2
XAND2X2_30 AND2X2_30/A AND2X2_30/B gnd AND2X2_30/Y vdd AND2X2
XNAND3X1_251 NAND3X1_251/A NAND3X1_251/B NAND3X1_251/C gnd AOI21X1_173/A vdd NAND3X1
XBUFX4_15 INVX8_2/Y gnd BUFX4_15/Y vdd BUFX4
XFILL_17_2 gnd vdd FILL
XOAI21X1_269 AND2X2_94/Y NOR2X1_170/Y INVX1_178/A gnd AOI21X1_193/A vdd OAI21X1
XNAND2X1_383 INVX1_245/Y AND2X2_111/A gnd NAND3X1_332/C vdd NAND2X1
XNOR2X1_302 NOR2X1_302/A NOR2X1_301/Y gnd BUFX2_229/A vdd NOR2X1
XFILL_31_3_0 gnd vdd FILL
XINVX2_90 gnd gnd INVX2_90/Y vdd INVX2
XFILL_29_5_1 gnd vdd FILL
XXNOR2X1_254 XNOR2X1_254/A XNOR2X1_254/B gnd XOR2X1_4/A vdd XNOR2X1
XFILL_9_6_1 gnd vdd FILL
XNOR2X1_69 gnd OR2X2_42/B gnd NOR3X1_36/B vdd NOR2X1
XNAND3X1_215 NAND3X1_213/A NAND3X1_215/B NAND3X1_214/Y gnd AOI21X1_149/A vdd NAND3X1
XBUFX2_216 BUFX2_216/A gnd BUFX2_216/Y vdd BUFX2
XOAI21X1_233 OAI21X1_233/A NAND3X1_240/Y INVX1_162/A gnd XOR2X1_140/A vdd OAI21X1
XNOR2X1_266 NOR2X1_266/A NOR2X1_265/Y gnd BUFX2_217/A vdd NOR2X1
XINVX2_54 INVX2_54/A gnd INVX2_54/Y vdd INVX2
XNAND2X1_347 INVX1_211/A NAND2X1_347/B gnd NOR3X1_59/B vdd NAND2X1
XINVX1_595 INVX1_595/A gnd INVX1_595/Y vdd INVX1
XBUFX2_180 BUFX2_180/A gnd BUFX2_180/Y vdd BUFX2
XNAND3X1_179 NAND3X1_179/A OAI21X1_172/Y NAND3X1_178/Y gnd NAND3X1_179/Y vdd NAND3X1
XNOR2X1_33 NOR2X1_33/A NOR2X1_33/B gnd NOR2X1_33/Y vdd NOR2X1
XXNOR2X1_218 bloque_bytes[39] OR2X2_144/B gnd AND2X2_182/B vdd XNOR2X1
XINVX2_18 INVX2_18/A gnd INVX2_18/Y vdd INVX2
XNAND2X1_311 gnd OR2X2_123/B gnd NAND3X1_281/B vdd NAND2X1
XOAI21X1_197 NOR3X1_48/C NOR3X1_48/B INVX1_133/Y gnd NAND3X1_206/A vdd OAI21X1
XNOR2X1_230 NOR2X1_230/A NOR2X1_230/B gnd BUFX2_205/A vdd NOR2X1
XOR2X2_1 gnd OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XBUFX2_144 gnd gnd BUFX2_144/Y vdd BUFX2
XNAND3X1_143 OAI21X1_135/Y OAI21X1_138/Y NAND3X1_142/Y gnd NAND3X1_143/Y vdd NAND3X1
XCLKBUF1_21 BUFX4_4/Y gnd CLKBUF1_21/Y vdd CLKBUF1
XINVX1_559 bloque_bytes[1] gnd INVX1_559/Y vdd INVX1
XFILL_28_8_0 gnd vdd FILL
XFILL_8_9_0 gnd vdd FILL
XOAI21X1_161 AND2X2_56/Y NOR3X1_43/B INVX1_110/Y gnd OAI21X1_161/Y vdd OAI21X1
XXNOR2X1_182 NOR2X1_285/Y XNOR2X1_182/B gnd XNOR2X1_183/A vdd XNOR2X1
XNOR2X1_194 NOR2X1_194/A NOR2X1_194/B gnd BUFX2_189/A vdd NOR2X1
XNAND2X1_275 INVX2_51/Y NAND3X1_254/C gnd XNOR2X1_125/A vdd NAND2X1
XDFFPOSX1_341 INVX1_400/A CLKBUF1_40/Y NAND2X1_686/Y gnd vdd DFFPOSX1
XNOR3X1_74 NOR3X1_74/A INVX2_67/Y NOR3X1_74/C gnd NOR3X1_74/Y vdd NOR3X1
XNAND3X1_107 NAND3X1_107/A NAND3X1_107/B NAND3X1_107/C gnd AOI21X1_77/A vdd NAND3X1
XXNOR2X1_146 XOR2X1_161/Y XOR2X1_149/Y gnd XNOR2X1_147/A vdd XNOR2X1
XINVX1_523 INVX1_523/A gnd INVX1_523/Y vdd INVX1
XFILL_36_5_1 gnd vdd FILL
XBUFX2_108 gnd gnd BUFX2_108/Y vdd BUFX2
XOAI21X1_125 AOI21X1_94/Y OAI21X1_125/B INVX1_84/Y gnd NAND3X1_130/C vdd OAI21X1
XNOR2X1_158 gnd OR2X2_113/B gnd NOR3X1_53/B vdd NOR2X1
XXNOR2X1_68 XNOR2X1_67/Y INVX2_32/Y gnd OR2X2_76/A vdd XNOR2X1
XNOR3X1_38 INVX1_78/Y NOR2X1_79/Y NOR3X1_38/C gnd NOR3X1_38/Y vdd NOR3X1
XNAND2X1_239 OR2X2_93/A OR2X2_93/B gnd NAND2X1_239/Y vdd NAND2X1
XINVX1_487 inicio gnd INVX1_487/Y vdd INVX1
XDFFPOSX1_305 XNOR2X1_174/B CLKBUF1_27/Y NAND3X1_513/Y gnd vdd DFFPOSX1
XXNOR2X1_32 AOI21X1_57/B INVX2_20/Y gnd OR2X2_44/A vdd XNOR2X1
XXOR2X1_302 bloque_bytes[45] bloque_bytes[5] gnd NOR2X1_414/A vdd XOR2X1
XXNOR2X1_110 XOR2X1_121/Y XOR2X1_109/Y gnd XNOR2X1_110/Y vdd XNOR2X1
XNAND2X1_203 OAI21X1_173/Y OR2X2_80/B gnd OR2X2_78/A vdd NAND2X1
XNOR2X1_122 OR2X2_84/A OR2X2_84/B gnd NOR2X1_122/Y vdd NOR2X1
XFILL_10_3_1 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XDFFPOSX1_269 INVX1_229/A CLKBUF1_31/Y NAND2X1_653/Y gnd vdd DFFPOSX1
XOR2X2_90 gnd OR2X2_90/B gnd OR2X2_90/Y vdd OR2X2
XXOR2X1_266 XOR2X1_266/A BUFX2_224/A gnd NOR2X1_330/B vdd XOR2X1
XOAI21X1_630 INVX1_579/A INVX1_580/Y INVX2_90/Y gnd AND2X2_188/A vdd OAI21X1
XINVX1_451 INVX1_451/A gnd INVX1_451/Y vdd INVX1
XXOR2X1_6 XOR2X1_6/A gnd gnd OR2X2_12/B vdd XOR2X1
XAOI21X1_403 INVX2_93/Y INVX1_598/Y NOR2X1_448/A gnd AOI21X1_403/Y vdd AOI21X1
XNAND2X1_167 NAND2X1_166/Y OR2X2_63/Y gnd OR2X2_64/A vdd NAND2X1
XFILL_35_8_0 gnd vdd FILL
XOR2X2_54 OR2X2_54/A OR2X2_54/B gnd INVX1_82/A vdd OR2X2
XAOI21X1_65 NAND3X1_89/Y AOI21X1_65/B AOI21X1_65/C gnd NAND3X1_92/B vdd AOI21X1
XDFFPOSX1_233 XOR2X1_141/B CLKBUF1_30/Y INVX1_543/A gnd vdd DFFPOSX1
XINVX1_415 INVX1_415/A gnd INVX1_415/Y vdd INVX1
XMUX2X1_12 BUFX2_12/A NOR2X1_4/A BUFX4_9/Y gnd MUX2X1_12/Y vdd MUX2X1
XNAND2X1_708 NAND2X1_708/A NAND2X1_708/B gnd XNOR2X1_254/A vdd NAND2X1
XOAI21X1_594 bloque_bytes[69] INVX1_498/Y OAI21X1_594/C gnd INVX1_576/A vdd OAI21X1
XXOR2X1_230 XOR2X1_230/A BUFX2_208/A gnd XOR2X1_230/Y vdd XOR2X1
XAOI21X1_367 INVX1_521/Y bloque_bytes[21] AOI21X1_367/C gnd INVX1_523/A vdd AOI21X1
XBUFX2_68 gnd gnd BUFX2_68/Y vdd BUFX2
XNAND3X1_540 AOI21X1_395/A NAND3X1_539/Y NAND3X1_540/C gnd AND2X2_197/B vdd NAND3X1
XNAND2X1_131 NAND2X1_130/Y OR2X2_48/Y gnd INVX1_73/A vdd NAND2X1
XDFFPOSX1_9 BUFX2_8/A CLKBUF1_4/Y NOR3X1_8/Y gnd vdd DFFPOSX1
XAOI21X1_29 AOI21X1_29/A AOI21X1_29/B OAI21X1_35/B gnd NAND3X1_38/B vdd AOI21X1
XOR2X2_18 gnd OR2X2_18/B gnd OR2X2_18/Y vdd OR2X2
XINVX1_379 INVX1_379/A gnd INVX1_379/Y vdd INVX1
XOAI21X1_558 BUFX2_236/A XOR2X1_284/Y INVX1_463/Y gnd OAI21X1_558/Y vdd OAI21X1
XDFFPOSX1_197 INVX1_112/A CLKBUF1_41/Y bloque_bytes[11] gnd vdd DFFPOSX1
XBUFX2_32 gnd gnd BUFX2_32/Y vdd BUFX2
XNAND2X1_672 bloque_bytes[7] OR2X2_141/A gnd AOI21X1_385/A vdd NAND2X1
XXOR2X1_194 XOR2X1_188/Y BUFX2_188/A gnd XOR2X1_194/Y vdd XOR2X1
XNAND2X1_92 OR2X2_32/B OR2X2_32/A gnd NAND2X1_93/A vdd NAND2X1
XAOI21X1_331 AND2X2_163/B NOR2X1_390/Y INVX1_477/A gnd NOR3X1_87/B vdd AOI21X1
XNAND3X1_504 XNOR2X1_209/Y NAND3X1_504/B AOI21X1_371/Y gnd NAND3X1_504/Y vdd NAND3X1
XDFFPOSX1_161 XOR2X1_51/B CLKBUF1_7/Y bloque_bytes[55] gnd vdd DFFPOSX1
XOAI21X1_77 NOR2X1_63/B NOR2X1_63/A NOR3X1_33/Y gnd OAI21X1_77/Y vdd OAI21X1
XDFFPOSX1_95 MUX2X1_6/B CLKBUF1_35/Y XNOR2X1_249/Y gnd vdd DFFPOSX1
XINVX2_5 target[0] gnd INVX2_5/Y vdd INVX2
XXOR2X1_158 XOR2X1_158/A BUFX2_173/A gnd NOR2X1_187/B vdd XOR2X1
XFILL_19_1_0 gnd vdd FILL
XINVX1_343 INVX1_343/A gnd INVX1_343/Y vdd INVX1
XOAI21X1_522 gnd NOR2X1_324/B INVX1_417/Y gnd AOI21X1_302/A vdd OAI21X1
XNAND2X1_636 INVX2_80/A INVX2_81/A gnd NAND2X1_636/Y vdd NAND2X1
XFILL_17_3_1 gnd vdd FILL
XOAI21X1_41 NOR2X1_37/A INVX1_31/Y INVX1_32/Y gnd OAI21X1_41/Y vdd OAI21X1
XNAND2X1_56 INVX2_16/A AND2X2_12/Y gnd AOI21X1_34/C vdd NAND2X1
XAOI21X1_295 NAND3X1_445/B AOI21X1_294/Y INVX1_408/Y gnd AOI21X1_296/A vdd AOI21X1
XNAND3X1_468 INVX1_445/A NAND3X1_466/Y INVX1_440/Y gnd AOI22X1_21/C vdd NAND3X1
XDFFPOSX1_125 INVX1_13/A CLKBUF1_16/Y bloque_bytes[83] gnd vdd DFFPOSX1
XDFFPOSX1_59 AND2X2_158/B CLKBUF1_38/Y NOR2X1_384/Y gnd vdd DFFPOSX1
XOAI21X1_486 OAI21X1_486/A INVX1_394/A INVX1_393/Y gnd AND2X2_141/A vdd OAI21X1
XINVX1_307 INVX1_307/A gnd INVX1_307/Y vdd INVX1
XXOR2X1_122 OR2X2_108/A gnd gnd XOR2X1_122/Y vdd XOR2X1
XNOR2X1_3 INVX1_3/A INVX2_4/Y gnd NOR2X1_3/Y vdd NOR2X1
XNAND2X1_600 NAND3X1_482/Y NAND3X1_483/Y gnd XOR2X1_296/B vdd NAND2X1
XAOI21X1_259 INVX1_331/A NAND3X1_388/Y INVX1_326/Y gnd NOR2X1_268/B vdd AOI21X1
XNAND2X1_20 INVX2_11/Y XNOR2X1_5/A gnd XNOR2X1_6/B vdd NAND2X1
XDFFPOSX1_23 BUFX2_22/A CLKBUF1_43/Y NOR3X1_22/Y gnd vdd DFFPOSX1
XNAND3X1_432 INVX1_380/Y AOI21X1_287/A NOR3X1_78/Y gnd AOI21X1_288/B vdd NAND3X1
XINVX1_271 INVX1_271/A gnd INVX1_271/Y vdd INVX1
XOAI21X1_450 OAI21X1_450/A INVX1_354/A INVX1_357/A gnd OAI21X1_450/Y vdd OAI21X1
XXOR2X1_66 XOR2X1_66/A OR2X2_52/A gnd OR2X2_60/B vdd XOR2X1
XNAND3X1_97 INVX1_67/A NAND3X1_97/B OR2X2_42/Y gnd AOI21X1_72/C vdd NAND3X1
XOR2X2_149 OR2X2_149/A OR2X2_149/B gnd OR2X2_149/Y vdd OR2X2
XFILL_30_1 gnd vdd FILL
XNAND2X1_564 XOR2X1_278/B NOR2X1_328/Y gnd AOI21X1_304/C vdd NAND2X1
XAOI21X1_223 AOI21X1_223/A AOI21X1_223/B INVX1_237/Y gnd AOI21X1_224/A vdd AOI21X1
XNAND3X1_396 INVX1_335/Y INVX1_338/Y AND2X2_129/A gnd NAND3X1_396/Y vdd NAND3X1
XFILL_14_8_1 gnd vdd FILL
XFILL_16_6_0 gnd vdd FILL
XXOR2X1_30 XOR2X1_30/A XOR2X1_30/B gnd XOR2X1_30/Y vdd XOR2X1
XNAND3X1_61 INVX1_45/A NAND2X1_80/Y OR2X2_26/Y gnd AOI21X1_48/C vdd NAND3X1
XNOR2X1_447 vdd gnd gnd NOR2X1_447/Y vdd NOR2X1
XINVX1_235 INVX1_235/A gnd INVX1_235/Y vdd INVX1
XAND2X2_166 INVX8_1/A AND2X2_166/B gnd AND2X2_166/Y vdd AND2X2
XOAI21X1_414 gnd XOR2X1_217/Y INVX1_321/A gnd INVX2_66/A vdd OAI21X1
XOR2X2_113 gnd OR2X2_113/B gnd OR2X2_113/Y vdd OR2X2
XNAND2X1_9 target[4] INVX2_2/Y gnd NAND2X1_9/Y vdd NAND2X1
XNAND2X1_528 XNOR2X1_191/B NAND2X1_528/B gnd NOR2X1_308/B vdd NAND2X1
XAOI21X1_187 NOR2X1_165/Y NAND3X1_272/Y INVX1_172/A gnd NOR2X1_167/A vdd AOI21X1
XNAND3X1_360 INVX1_287/A NAND3X1_360/B NAND2X1_424/Y gnd NAND3X1_360/Y vdd NAND3X1
XFILL_24_3_1 gnd vdd FILL
XFILL_26_1_0 gnd vdd FILL
XOAI22X1_8 INVX4_1/Y INVX1_7/A INVX1_8/A INVX2_3/Y gnd OAI22X1_8/Y vdd OAI22X1
XFILL_4_4_1 gnd vdd FILL
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XFILL_6_2_0 gnd vdd FILL
XINVX1_199 INVX1_199/A gnd INVX1_199/Y vdd INVX1
XOAI21X1_378 gnd XOR2X1_200/Y INVX1_284/A gnd INVX1_287/A vdd OAI21X1
XAND2X2_130 NOR2X1_274/Y INVX1_339/Y gnd NOR3X1_74/A vdd AND2X2
XNAND3X1_25 INVX1_23/A NAND3X1_25/B OR2X2_10/Y gnd NAND3X1_26/C vdd NAND3X1
XNOR2X1_411 NOR2X1_411/A NOR2X1_411/B gnd NOR2X1_411/Y vdd NOR2X1
XOAI22X1_10 INVX2_10/Y target[3] INVX1_9/Y target[2] gnd NOR2X1_15/B vdd OAI22X1
XNAND2X1_492 NAND2X1_491/Y INVX1_354/Y gnd INVX1_355/A vdd NAND2X1
XAOI21X1_151 NOR2X1_135/Y AOI21X1_151/B INVX1_139/A gnd NOR2X1_137/A vdd AOI21X1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XNAND3X1_324 INVX1_234/A INVX1_232/Y INVX1_233/Y gnd NAND3X1_324/Y vdd NAND3X1
XNOR2X1_375 BUFX4_15/Y NOR3X1_92/A gnd NOR2X1_375/Y vdd NOR2X1
XINVX1_163 INVX1_163/A gnd INVX1_163/Y vdd INVX1
XOAI21X1_342 NOR3X1_64/A NOR3X1_64/C INVX2_62/A gnd NOR2X1_217/A vdd OAI21X1
XNAND2X1_456 OAI21X1_412/Y NAND3X1_383/Y gnd XOR2X1_232/A vdd NAND2X1
XAOI21X1_115 NOR2X1_105/Y AOI21X1_115/B INVX1_106/A gnd NOR2X1_107/A vdd AOI21X1
XAND2X2_67 OR2X2_85/A OR2X2_85/B gnd AND2X2_67/Y vdd AND2X2
XNAND3X1_288 INVX1_180/A NAND3X1_286/B OR2X2_125/Y gnd OR2X2_128/B vdd NAND3X1
XINVX1_127 INVX1_127/A gnd OR2X2_87/B vdd INVX1
XOAI21X1_306 gnd XOR2X1_165/Y INVX1_210/A gnd INVX1_212/A vdd OAI21X1
XFILL_23_6_0 gnd vdd FILL
XNOR2X1_339 gnd NOR2X1_339/B gnd NOR2X1_339/Y vdd NOR2X1
XNAND2X1_420 NAND2X1_420/A NAND3X1_358/B gnd BUFX2_207/A vdd NAND2X1
XFILL_3_7_0 gnd vdd FILL
XFILL_21_8_1 gnd vdd FILL
XFILL_1_9_1 gnd vdd FILL
XAND2X2_31 OR2X2_37/A OR2X2_37/B gnd AND2X2_31/Y vdd AND2X2
XBUFX2_253 BUFX2_253/A gnd BUFX2_253/Y vdd BUFX2
XNAND3X1_252 INVX1_158/A NAND3X1_252/B OR2X2_109/Y gnd OR2X2_112/B vdd NAND3X1
XBUFX4_16 INVX8_2/Y gnd BUFX4_16/Y vdd BUFX4
XOAI21X1_270 AND2X2_95/Y NOR2X1_172/Y INVX1_179/A gnd NAND3X1_283/C vdd OAI21X1
XFILL_33_1_0 gnd vdd FILL
XNAND2X1_384 INVX1_246/Y NOR2X1_216/Y gnd NAND2X1_385/B vdd NAND2X1
XNOR2X1_303 gnd XOR2X1_246/Y gnd NOR2X1_303/Y vdd NOR2X1
XFILL_31_3_1 gnd vdd FILL
XINVX2_91 INVX2_91/A gnd INVX2_91/Y vdd INVX2
XNAND3X1_216 INVX1_136/A NAND2X1_239/Y OR2X2_93/Y gnd OR2X2_96/B vdd NAND3X1
XXNOR2X1_255 XNOR2X1_255/A AND2X2_197/Y gnd XOR2X1_6/A vdd XNOR2X1
XNOR2X1_70 gnd OR2X2_43/B gnd NOR2X1_70/Y vdd NOR2X1
XBUFX2_217 BUFX2_217/A gnd BUFX2_217/Y vdd BUFX2
XINVX2_55 INVX2_55/A gnd INVX2_55/Y vdd INVX2
XOAI21X1_234 AND2X2_82/Y NOR2X1_150/Y INVX1_156/Y gnd AOI21X1_168/A vdd OAI21X1
XNOR2X1_267 gnd NOR2X1_267/B gnd NOR2X1_267/Y vdd NOR2X1
XNAND2X1_348 INVX1_210/A NOR2X1_195/Y gnd NAND3X1_308/C vdd NAND2X1
XINVX1_596 INVX1_596/A gnd OR2X2_161/B vdd INVX1
XBUFX2_181 BUFX2_181/A gnd BUFX2_181/Y vdd BUFX2
XNAND3X1_180 INVX1_114/A NAND2X1_201/Y OR2X2_77/Y gnd OR2X2_80/B vdd NAND3X1
XNOR2X1_34 XOR2X1_3/A OR2X2_13/B gnd NOR2X1_34/Y vdd NOR2X1
XXNOR2X1_219 bloque_bytes[24] INVX1_501/A gnd NAND3X1_503/B vdd XNOR2X1
XOAI21X1_198 NOR3X1_48/Y NOR2X1_133/A NAND2X1_231/B gnd OAI21X1_198/Y vdd OAI21X1
XINVX2_19 INVX2_19/A gnd INVX2_19/Y vdd INVX2
XNAND2X1_312 BUFX2_171/A OR2X2_124/B gnd AOI21X1_196/A vdd NAND2X1
XNOR2X1_231 gnd XOR2X1_192/Y gnd NOR2X1_231/Y vdd NOR2X1
XOR2X2_2 gnd OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XBUFX2_145 gnd gnd BUFX2_145/Y vdd BUFX2
XNAND3X1_144 INVX1_92/A NAND2X1_163/Y OR2X2_61/Y gnd OR2X2_64/B vdd NAND3X1
XCLKBUF1_22 BUFX4_4/Y gnd CLKBUF1_22/Y vdd CLKBUF1
XINVX1_560 INVX1_560/A gnd INVX1_560/Y vdd INVX1
XXNOR2X1_183 XNOR2X1_183/A OAI21X1_447/Y gnd INVX1_357/A vdd XNOR2X1
XFILL_30_6_0 gnd vdd FILL
XFILL_28_8_1 gnd vdd FILL
XFILL_8_9_1 gnd vdd FILL
XNOR2X1_195 gnd XOR2X1_165/Y gnd NOR2X1_195/Y vdd NOR2X1
XOAI21X1_162 NOR3X1_44/Y NOR2X1_113/A NOR3X1_43/Y gnd NAND2X1_195/B vdd OAI21X1
XNAND2X1_276 AND2X2_84/B AND2X2_84/A gnd OAI21X1_239/B vdd NAND2X1
XINVX1_524 bloque_bytes[62] gnd INVX1_524/Y vdd INVX1
XNAND3X1_108 INVX1_70/A NAND3X1_106/B OR2X2_45/Y gnd OR2X2_48/B vdd NAND3X1
XBUFX2_109 gnd gnd BUFX2_109/Y vdd BUFX2
XDFFPOSX1_342 INVX1_405/A CLKBUF1_45/Y NAND2X1_687/Y gnd vdd DFFPOSX1
XNOR3X1_75 NOR3X1_75/A INVX1_361/A NOR3X1_75/C gnd NOR3X1_75/Y vdd NOR3X1
XXNOR2X1_147 XNOR2X1_147/A OR2X2_127/Y gnd INVX1_186/A vdd XNOR2X1
XXNOR2X1_69 XNOR2X1_69/A XNOR2X1_69/B gnd OR2X2_77/A vdd XNOR2X1
XOAI21X1_126 NOR2X1_87/A INVX1_86/Y INVX1_87/Y gnd NAND2X1_152/B vdd OAI21X1
XNOR2X1_159 gnd OR2X2_114/B gnd NOR3X1_54/B vdd NOR2X1
XNAND2X1_240 AOI21X1_149/A AOI21X1_149/B gnd INVX2_46/A vdd NAND2X1
XNOR3X1_39 INVX1_88/Y NOR2X1_88/Y NOR3X1_39/C gnd NOR3X1_39/Y vdd NOR3X1
XINVX1_488 INVX1_488/A gnd INVX1_488/Y vdd INVX1
XDFFPOSX1_306 INVX1_320/A CLKBUF1_46/Y OR2X2_145/A gnd vdd DFFPOSX1
XXNOR2X1_33 AOI21X1_57/C NAND3X1_60/C gnd OR2X2_45/A vdd XNOR2X1
XXOR2X1_303 bloque_bytes[46] bloque_bytes[6] gnd XOR2X1_303/Y vdd XOR2X1
XXNOR2X1_111 XNOR2X1_110/Y OR2X2_95/Y gnd INVX1_142/A vdd XNOR2X1
XNOR2X1_123 NOR2X1_123/A NOR3X1_46/Y gnd NOR2X1_123/Y vdd NOR2X1
XFILL_12_1_1 gnd vdd FILL
XNAND2X1_204 OR2X2_79/B OR2X2_79/A gnd NAND2X1_204/Y vdd NAND2X1
XDFFPOSX1_270 INVX1_234/A CLKBUF1_11/Y XNOR2X1_238/A gnd vdd DFFPOSX1
XOR2X2_91 gnd OR2X2_91/B gnd OR2X2_91/Y vdd OR2X2
XXOR2X1_267 XOR2X1_267/A BUFX2_225/A gnd NOR2X1_331/B vdd XOR2X1
XOAI21X1_631 OAI21X1_631/A INVX1_581/Y INVX1_582/Y gnd AND2X2_191/A vdd OAI21X1
XINVX1_452 INVX1_452/A gnd INVX1_452/Y vdd INVX1
XXOR2X1_7 XOR2X1_7/A vdd gnd OR2X2_13/B vdd XOR2X1
XAOI21X1_404 INVX2_92/Y XNOR2X1_252/A XNOR2X1_253/A gnd NAND3X1_548/A vdd AOI21X1
XNAND2X1_168 OR2X2_64/B OR2X2_64/A gnd NAND2X1_168/Y vdd NAND2X1
XFILL_35_8_1 gnd vdd FILL
XAOI21X1_66 OR2X2_38/B OR2X2_38/A AND2X2_30/B gnd NOR2X1_65/A vdd AOI21X1
XOR2X2_55 OR2X2_55/A OR2X2_55/B gnd OR2X2_55/Y vdd OR2X2
XOAI21X1_595 bloque_bytes[70] INVX1_499/Y OAI21X1_595/C gnd INVX1_577/A vdd OAI21X1
XDFFPOSX1_234 INVX2_53/A CLKBUF1_47/Y INVX1_507/A gnd vdd DFFPOSX1
XINVX1_416 INVX1_416/A gnd INVX1_416/Y vdd INVX1
XMUX2X1_13 BUFX2_13/A INVX2_2/A BUFX4_9/Y gnd NOR3X1_13/B vdd MUX2X1
XNAND2X1_709 INVX1_598/A NAND2X1_709/B gnd OAI21X1_639/A vdd NAND2X1
XBUFX2_69 gnd gnd BUFX2_69/Y vdd BUFX2
XXOR2X1_231 AND2X2_125/Y BUFX2_209/A gnd XOR2X1_231/Y vdd XOR2X1
XNAND2X1_132 INVX2_28/A AND2X2_36/Y gnd AOI21X1_82/C vdd NAND2X1
XAOI21X1_368 INVX1_524/Y bloque_bytes[22] AOI21X1_368/C gnd INVX1_526/A vdd AOI21X1
XNAND3X1_541 INVX1_593/A NAND3X1_541/B OR2X2_158/Y gnd NAND3X1_542/B vdd NAND3X1
XDFFPOSX1_198 INVX1_113/A CLKBUF1_41/Y bloque_bytes[12] gnd vdd DFFPOSX1
XOR2X2_19 gnd OR2X2_19/B gnd OR2X2_19/Y vdd OR2X2
XAOI21X1_30 OR2X2_14/B OR2X2_14/A AND2X2_12/B gnd NOR2X1_35/A vdd AOI21X1
XFILL_11_4_0 gnd vdd FILL
XINVX1_380 INVX1_380/A gnd INVX1_380/Y vdd INVX1
XOAI21X1_559 BUFX2_236/A XOR2X1_284/Y INVX1_463/A gnd AOI22X1_22/B vdd OAI21X1
XXOR2X1_195 AND2X2_109/Y BUFX2_189/A gnd XOR2X1_195/Y vdd XOR2X1
XNAND2X1_673 INVX1_544/A OAI21X1_591/Y gnd NAND2X1_673/Y vdd NAND2X1
XBUFX2_33 gnd gnd BUFX2_33/Y vdd BUFX2
XNAND2X1_93 NAND2X1_93/A OR2X2_32/Y gnd INVX1_51/A vdd NAND2X1
XOAI21X1_78 NOR3X1_34/C NOR3X1_34/B INVX1_56/Y gnd OAI21X1_78/Y vdd OAI21X1
XAOI21X1_332 AND2X2_164/B NOR2X1_395/B INVX1_478/A gnd NOR3X1_88/B vdd AOI21X1
XNAND3X1_505 XNOR2X1_210/Y XNOR2X1_221/Y NAND2X1_652/B gnd AOI21X1_381/C vdd NAND3X1
XINVX2_6 target[3] gnd INVX2_6/Y vdd INVX2
XDFFPOSX1_162 INVX2_26/A CLKBUF1_12/Y bloque_bytes[40] gnd vdd DFFPOSX1
XDFFPOSX1_96 MUX2X1_7/B CLKBUF1_35/Y NAND2X1_703/Y gnd vdd DFFPOSX1
XINVX1_344 INVX1_344/A gnd INVX1_344/Y vdd INVX1
XFILL_1_0_0 gnd vdd FILL
XNAND2X1_637 INVX2_80/A NOR2X1_406/Y gnd OR2X2_130/A vdd NAND2X1
XXOR2X1_159 XOR2X1_159/A BUFX2_174/A gnd NOR2X1_189/B vdd XOR2X1
XFILL_19_1_1 gnd vdd FILL
XOAI21X1_523 BUFX2_229/A NOR2X1_331/B INVX1_429/A gnd XNOR2X1_199/B vdd OAI21X1
XNAND2X1_57 NAND2X1_57/A OAI21X1_41/Y gnd XOR2X1_29/A vdd NAND2X1
XOAI21X1_42 AND2X2_14/Y NOR3X1_29/B INVX1_33/Y gnd NAND3X1_42/B vdd OAI21X1
XDFFPOSX1_60 AND2X2_159/B CLKBUF1_37/Y DFFPOSX1_60/D gnd vdd DFFPOSX1
XAOI21X1_296 AOI21X1_296/A AOI21X1_296/B AOI21X1_296/C gnd OAI21X1_505/A vdd AOI21X1
XNAND3X1_469 INVX1_445/A OAI21X1_539/Y NAND2X1_579/Y gnd NAND3X1_469/Y vdd NAND3X1
XDFFPOSX1_126 INVX1_14/A CLKBUF1_5/Y bloque_bytes[84] gnd vdd DFFPOSX1
XOAI21X1_487 NOR2X1_305/A NOR3X1_77/Y AOI21X1_289/Y gnd NAND3X1_434/C vdd OAI21X1
XINVX1_308 BUFX2_203/A gnd INVX1_308/Y vdd INVX1
XXOR2X1_123 BUFX2_164/A gnd gnd OR2X2_105/B vdd XOR2X1
XNAND2X1_601 INVX1_455/A NOR2X1_348/Y gnd NAND2X1_601/Y vdd NAND2X1
XNOR2X1_4 NOR2X1_4/A INVX2_6/Y gnd NOR2X1_4/Y vdd NOR2X1
XNAND2X1_21 gnd OR2X2_1/B gnd NAND3X1_5/B vdd NAND2X1
XNAND3X1_433 INVX1_383/A OAI21X1_479/Y NAND3X1_433/C gnd NAND2X1_531/A vdd NAND3X1
XAOI21X1_260 NAND3X1_394/B NAND3X1_389/Y INVX1_326/A gnd NOR2X1_268/A vdd AOI21X1
XFILL_8_1 gnd vdd FILL
XDFFPOSX1_24 BUFX2_23/A CLKBUF1_43/Y NOR3X1_23/Y gnd vdd DFFPOSX1
XXOR2X1_67 XOR2X1_67/A OR2X2_53/A gnd OR2X2_61/B vdd XOR2X1
XINVX1_272 INVX1_272/A gnd INVX1_272/Y vdd INVX1
XOAI21X1_451 gnd XOR2X1_234/Y INVX1_358/A gnd NAND2X1_496/A vdd OAI21X1
XNAND3X1_98 NAND3X1_99/B NAND3X1_96/A AOI21X1_72/C gnd NAND3X1_98/Y vdd NAND3X1
XOR2X2_150 OR2X2_145/A OR2X2_150/B gnd OR2X2_150/Y vdd OR2X2
XNAND2X1_565 INVX1_429/Y NOR2X1_331/Y gnd NAND2X1_565/Y vdd NAND2X1
XFILL_30_2 gnd vdd FILL
XAOI21X1_224 AOI21X1_224/A AOI21X1_224/B AOI21X1_224/C gnd OAI21X1_334/A vdd AOI21X1
XFILL_16_6_1 gnd vdd FILL
XFILL_18_4_0 gnd vdd FILL
XNAND3X1_397 INVX2_67/A NAND3X1_397/B NAND2X1_478/Y gnd NOR3X1_73/A vdd NAND3X1
XINVX1_236 INVX1_236/A gnd INVX1_236/Y vdd INVX1
XOAI21X1_415 NOR3X1_72/C INVX2_66/Y NOR3X1_72/A gnd AND2X2_128/A vdd OAI21X1
XNOR2X1_448 NOR2X1_448/A INVX2_93/A gnd XOR2X1_317/B vdd NOR2X1
XXOR2X1_31 XOR2X1_15/A XOR2X1_31/B gnd XOR2X1_31/Y vdd XOR2X1
XNAND3X1_62 NAND3X1_63/B OAI21X1_62/C AOI21X1_48/C gnd NAND2X1_81/A vdd NAND3X1
XAND2X2_167 BUFX4_32/Y AND2X2_167/B gnd AND2X2_167/Y vdd AND2X2
XNAND2X1_529 INVX1_390/Y NOR2X1_308/B gnd NAND2X1_529/Y vdd NAND2X1
XOR2X2_114 gnd OR2X2_114/B gnd OR2X2_114/Y vdd OR2X2
XAOI21X1_188 INVX2_54/Y INVX1_173/Y NOR2X1_161/A gnd AOI21X1_190/A vdd AOI21X1
XFILL_6_2_1 gnd vdd FILL
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XFILL_8_0_0 gnd vdd FILL
XNAND3X1_361 INVX1_288/A AOI21X1_245/B INVX1_287/Y gnd INVX1_294/A vdd NAND3X1
XFILL_26_1_1 gnd vdd FILL
XOAI22X1_9 INVX1_7/Y target[5] INVX1_8/Y target[4] gnd NOR2X1_14/B vdd OAI22X1
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XOAI21X1_379 NOR3X1_67/A NOR3X1_67/B OAI21X1_385/B gnd NOR2X1_242/A vdd OAI21X1
XAND2X2_131 NOR2X1_275/Y INVX1_340/Y gnd NOR3X1_74/C vdd AND2X2
XNAND3X1_26 NAND3X1_26/A NAND2X1_41/B NAND3X1_26/C gnd NAND3X1_26/Y vdd NAND3X1
XNOR2X1_412 XOR2X1_300/Y NOR2X1_412/B gnd INVX1_538/A vdd NOR2X1
XNAND2X1_493 NAND3X1_407/Y AOI22X1_16/C gnd AOI21X1_273/C vdd NAND2X1
XNAND3X1_325 INVX1_236/A NAND3X1_323/Y INVX1_231/Y gnd AOI22X1_10/C vdd NAND3X1
XAOI21X1_152 INVX2_45/Y INVX1_140/Y NOR2X1_131/A gnd AOI21X1_152/Y vdd AOI21X1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XNOR2X1_376 BUFX4_15/Y INVX1_484/Y gnd NOR2X1_376/Y vdd NOR2X1
XFILL_15_9_0 gnd vdd FILL
XINVX1_164 INVX1_164/A gnd INVX1_164/Y vdd INVX1
XOAI21X1_343 gnd XOR2X1_183/Y INVX1_248/Y gnd OAI21X1_343/Y vdd OAI21X1
XNAND2X1_457 INVX1_320/Y AND2X2_126/A gnd NAND3X1_384/B vdd NAND2X1
XAOI21X1_116 INVX2_36/Y INVX1_107/Y NOR2X1_101/A gnd AOI21X1_118/A vdd AOI21X1
XNAND3X1_289 NAND3X1_289/A OR2X2_128/B OR2X2_126/B gnd AOI21X1_197/B vdd NAND3X1
XAND2X2_68 gnd OR2X2_89/B gnd NOR3X1_47/C vdd AND2X2
XINVX1_128 INVX1_128/A gnd INVX1_128/Y vdd INVX1
XOAI21X1_307 BUFX2_179/A INVX1_214/A INVX1_215/A gnd INVX1_217/A vdd OAI21X1
XFILL_25_4_0 gnd vdd FILL
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XFILL_5_5_0 gnd vdd FILL
XFILL_23_6_1 gnd vdd FILL
XNAND2X1_421 INVX1_283/Y NOR2X1_239/Y gnd NAND3X1_358/C vdd NAND2X1
XNOR2X1_340 NOR2X1_340/A NOR2X1_340/B gnd NOR2X1_340/Y vdd NOR2X1
XFILL_3_7_1 gnd vdd FILL
XAND2X2_32 gnd OR2X2_41/B gnd NOR3X1_35/C vdd AND2X2
XBUFX2_254 XOR2X1_61/A gnd BUFX2_254/Y vdd BUFX2
XNAND3X1_253 NAND3X1_253/A OR2X2_112/B OR2X2_110/B gnd AOI21X1_173/B vdd NAND3X1
XBUFX4_17 INVX8_2/Y gnd BUFX4_17/Y vdd BUFX4
XOAI21X1_271 AND2X2_95/Y NOR2X1_172/Y INVX1_179/Y gnd NAND3X1_287/A vdd OAI21X1
XNOR2X1_304 NOR2X1_304/A NOR2X1_304/B gnd NOR2X1_304/Y vdd NOR2X1
XFILL_33_1_1 gnd vdd FILL
XINVX2_92 INVX2_92/A gnd INVX2_92/Y vdd INVX2
XNAND2X1_385 INVX1_249/A NAND2X1_385/B gnd INVX1_247/A vdd NAND2X1
XNAND3X1_217 NAND3X1_217/A OR2X2_96/B OR2X2_94/B gnd AOI21X1_149/B vdd NAND3X1
XBUFX2_218 BUFX2_218/A gnd BUFX2_218/Y vdd BUFX2
XXNOR2X1_256 XNOR2X1_256/A INVX2_94/Y gnd XOR2X1_7/A vdd XNOR2X1
XNOR2X1_71 NOR2X1_71/A INVX2_27/A gnd NOR2X1_71/Y vdd NOR2X1
XNAND2X1_349 INVX1_210/Y NOR2X1_195/Y gnd NAND3X1_309/B vdd NAND2X1
XINVX2_56 INVX2_56/A gnd INVX2_56/Y vdd INVX2
XOAI21X1_235 AND2X2_82/Y NOR2X1_150/Y INVX1_156/A gnd AOI21X1_169/A vdd OAI21X1
XNOR2X1_268 NOR2X1_268/A NOR2X1_268/B gnd NOR2X1_268/Y vdd NOR2X1
XINVX1_597 INVX1_597/A gnd INVX1_597/Y vdd INVX1
XBUFX2_182 BUFX2_182/A gnd BUFX2_182/Y vdd BUFX2
XFILL_22_9_0 gnd vdd FILL
XNAND3X1_181 OAI21X1_173/Y OR2X2_80/B OR2X2_78/B gnd NAND3X1_181/Y vdd NAND3X1
XNOR2X1_35 NOR2X1_35/A INVX1_27/Y gnd NOR2X1_35/Y vdd NOR2X1
XOAI21X1_199 OAI21X1_199/A XNOR2X1_106/B INVX1_140/A gnd XOR2X1_120/A vdd OAI21X1
XXNOR2X1_220 bloque_bytes[25] INVX1_502/A gnd NAND3X1_504/B vdd XNOR2X1
XINVX2_20 INVX2_20/A gnd INVX2_20/Y vdd INVX2
XNAND2X1_313 INVX2_57/Y NAND2X1_313/B gnd XNOR2X1_143/A vdd NAND2X1
XNOR2X1_232 NOR2X1_232/A NOR2X1_232/B gnd NOR2X1_232/Y vdd NOR2X1
XNAND3X1_145 OAI21X1_139/Y OR2X2_64/B OR2X2_62/B gnd NAND3X1_145/Y vdd NAND3X1
XFILL_32_4_0 gnd vdd FILL
XFILL_30_6_1 gnd vdd FILL
XBUFX2_146 gnd gnd BUFX2_146/Y vdd BUFX2
XOR2X2_3 gnd OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XCLKBUF1_23 BUFX4_5/Y gnd CLKBUF1_23/Y vdd CLKBUF1
XINVX1_561 INVX1_561/A gnd INVX1_561/Y vdd INVX1
XXNOR2X1_184 NOR2X1_290/A XNOR2X1_184/B gnd BUFX2_226/A vdd XNOR2X1
XNOR2X1_196 NOR2X1_196/A NOR2X1_196/B gnd NOR2X1_196/Y vdd NOR2X1
XOAI21X1_163 AND2X2_57/Y NOR3X1_44/B INVX1_111/Y gnd NAND3X1_170/A vdd OAI21X1
XNAND2X1_277 BUFX2_164/A OR2X2_109/B gnd NAND3X1_252/B vdd NAND2X1
XNOR3X1_76 NOR3X1_76/A INVX2_68/Y NOR3X1_76/C gnd NOR3X1_76/Y vdd NOR3X1
XNAND3X1_109 OAI21X1_105/Y OR2X2_48/B OR2X2_46/B gnd AOI21X1_77/B vdd NAND3X1
XINVX1_525 INVX1_525/A gnd INVX1_525/Y vdd INVX1
XBUFX2_110 gnd gnd BUFX2_110/Y vdd BUFX2
XDFFPOSX1_343 INVX1_406/A CLKBUF1_45/Y NAND3X1_514/Y gnd vdd DFFPOSX1
XXNOR2X1_148 NOR2X1_182/A XNOR2X1_148/B gnd BUFX2_186/A vdd XNOR2X1
XXNOR2X1_70 XNOR2X1_70/A XNOR2X1_70/B gnd XOR2X1_98/B vdd XNOR2X1
XOAI21X1_127 NOR3X1_39/C NOR2X1_88/Y INVX1_88/Y gnd NAND3X1_132/B vdd OAI21X1
XNOR2X1_160 gnd OR2X2_115/B gnd NOR2X1_160/Y vdd NOR2X1
XNAND2X1_241 NAND3X1_217/A OR2X2_96/B gnd OR2X2_94/A vdd NAND2X1
XNOR3X1_40 INVX1_89/Y NOR2X1_89/Y AND2X2_45/Y gnd NOR3X1_40/Y vdd NOR3X1
XDFFPOSX1_307 INVX1_321/A CLKBUF1_8/Y OR2X2_151/A gnd vdd DFFPOSX1
XINVX1_489 INVX1_489/A gnd INVX1_489/Y vdd INVX1
XXOR2X1_304 bloque_bytes[29] INVX1_533/A gnd NOR2X1_426/A vdd XOR2X1
XXNOR2X1_112 gnd XOR2X1_112/Y gnd NAND2X1_248/B vdd XNOR2X1
XFILL_21_1 gnd vdd FILL
XXNOR2X1_34 NAND3X1_75/B OAI21X1_68/B gnd BUFX2_253/A vdd XNOR2X1
XFILL_29_9_0 gnd vdd FILL
XNOR2X1_124 OR2X2_85/A OR2X2_85/B gnd NOR2X1_124/Y vdd NOR2X1
XNAND2X1_205 NAND2X1_204/Y OR2X2_79/Y gnd OR2X2_80/A vdd NAND2X1
XDFFPOSX1_271 INVX1_235/A CLKBUF1_31/Y NOR2X1_426/B gnd vdd DFFPOSX1
XOR2X2_92 OR2X2_92/A OR2X2_92/B gnd OR2X2_92/Y vdd OR2X2
XINVX1_453 INVX1_453/A gnd INVX1_453/Y vdd INVX1
XXOR2X1_268 XOR2X1_268/A BUFX2_226/A gnd NOR2X1_333/B vdd XOR2X1
XOAI21X1_632 INVX1_585/A NOR2X1_350/Y INVX1_587/A gnd OAI21X1_632/Y vdd OAI21X1
XXOR2X1_8 XOR2X1_8/A vdd gnd XOR2X1_8/Y vdd XOR2X1
XAOI21X1_405 AOI21X1_403/Y NAND3X1_548/Y OAI21X1_648/B gnd OAI21X1_650/A vdd AOI21X1
XNAND2X1_169 NAND2X1_168/Y OR2X2_64/Y gnd INVX1_95/A vdd NAND2X1
XAOI21X1_67 NOR2X1_65/Y AOI21X1_67/B INVX1_62/A gnd NOR2X1_67/A vdd AOI21X1
XOR2X2_56 OR2X2_56/A OR2X2_56/B gnd OR2X2_56/Y vdd OR2X2
XDFFPOSX1_235 INVX1_165/A CLKBUF1_47/Y INVX1_510/A gnd vdd DFFPOSX1
XOAI21X1_596 bloque_bytes[71] INVX1_500/Y OAI21X1_596/C gnd OR2X2_144/A vdd OAI21X1
XINVX1_417 INVX1_417/A gnd INVX1_417/Y vdd INVX1
XMUX2X1_14 BUFX2_14/A INVX2_1/A BUFX4_9/Y gnd MUX2X1_14/Y vdd MUX2X1
XNAND2X1_710 vdd gnd gnd NAND3X1_537/B vdd NAND2X1
XBUFX2_70 gnd gnd BUFX2_70/Y vdd BUFX2
XXOR2X1_232 XOR2X1_232/A BUFX2_210/A gnd XOR2X1_232/Y vdd XOR2X1
XNAND3X1_542 NAND3X1_544/A NAND3X1_542/B NAND3X1_542/C gnd AND2X2_197/A vdd NAND3X1
XNAND2X1_133 NAND3X1_112/Y OAI21X1_109/Y gnd XOR2X1_69/A vdd NAND2X1
XAOI21X1_369 INVX1_527/Y bloque_bytes[23] OAI21X1_608/Y gnd INVX1_529/A vdd AOI21X1
XAOI21X1_31 NOR2X1_35/Y NAND3X1_38/Y INVX1_29/A gnd NOR2X1_37/A vdd AOI21X1
XFILL_13_2_0 gnd vdd FILL
XDFFPOSX1_199 INVX1_114/A CLKBUF1_10/Y bloque_bytes[13] gnd vdd DFFPOSX1
XOR2X2_20 OR2X2_20/A OR2X2_20/B gnd OR2X2_20/Y vdd OR2X2
XFILL_11_4_1 gnd vdd FILL
XXOR2X1_196 XOR2X1_196/A BUFX2_190/A gnd XOR2X1_196/Y vdd XOR2X1
XOAI21X1_560 gnd NOR2X1_348/B INVX1_455/Y gnd AOI21X1_318/A vdd OAI21X1
XINVX1_381 INVX1_381/A gnd INVX1_381/Y vdd INVX1
XNAND2X1_674 INVX1_544/Y NAND2X1_659/B gnd AOI21X1_388/B vdd NAND2X1
XBUFX2_34 gnd gnd BUFX2_34/Y vdd BUFX2
XNAND2X1_94 INVX2_22/A AND2X2_24/Y gnd NAND2X1_94/Y vdd NAND2X1
XOAI21X1_79 NOR2X1_63/B NOR2X1_63/A NAND3X1_77/Y gnd OAI21X1_79/Y vdd OAI21X1
XAOI21X1_333 INVX2_75/A INVX2_83/A OAI21X1_576/Y gnd AOI21X1_333/Y vdd AOI21X1
XNAND3X1_506 XNOR2X1_211/Y NAND3X1_506/B NAND2X1_653/B gnd AOI21X1_382/C vdd NAND3X1
XDFFPOSX1_97 MUX2X1_8/B CLKBUF1_4/Y DFFPOSX1_97/D gnd vdd DFFPOSX1
XINVX2_7 target[2] gnd INVX2_7/Y vdd INVX2
XDFFPOSX1_163 INVX1_66/A CLKBUF1_12/Y bloque_bytes[41] gnd vdd DFFPOSX1
XFILL_36_9_0 gnd vdd FILL
XINVX1_345 INVX1_345/A gnd INVX1_345/Y vdd INVX1
XOAI21X1_524 AOI21X1_304/Y INVX1_432/A INVX1_431/Y gnd AND2X2_149/A vdd OAI21X1
XFILL_1_0_1 gnd vdd FILL
XNAND2X1_638 bloque_bytes[72] bloque_bytes[32] gnd AOI21X1_370/A vdd NAND2X1
XXOR2X1_160 XOR2X1_160/A XOR2X1_160/B gnd BUFX2_182/A vdd XOR2X1
XAOI21X1_297 NAND3X1_443/Y NAND3X1_444/Y NAND2X1_550/Y gnd OAI21X1_506/C vdd AOI21X1
XOAI21X1_43 NOR2X1_43/B NOR2X1_43/A NOR3X1_29/Y gnd NAND2X1_62/B vdd OAI21X1
XNAND2X1_58 INVX2_17/Y NAND2X1_58/B gnd NAND3X1_42/C vdd NAND2X1
XDFFPOSX1_127 INVX1_15/A CLKBUF1_38/Y bloque_bytes[85] gnd vdd DFFPOSX1
XDFFPOSX1_61 INVX2_74/A CLKBUF1_9/Y AOI21X1_324/Y gnd vdd DFFPOSX1
XNAND3X1_470 AOI22X1_21/B INVX1_447/A INVX1_445/Y gnd NAND3X1_470/Y vdd NAND3X1
XOAI21X1_488 OAI21X1_488/A INVX1_392/A INVX1_395/A gnd NAND2X1_532/A vdd OAI21X1
XINVX1_309 INVX1_309/A gnd INVX1_309/Y vdd INVX1
XXOR2X1_124 BUFX2_165/A gnd gnd AND2X2_81/B vdd XOR2X1
XNOR2X1_5 NOR2X1_5/A INVX2_7/Y gnd NOR2X1_5/Y vdd NOR2X1
XNAND2X1_602 XOR2X1_296/B NOR2X1_352/Y gnd NAND2X1_602/Y vdd NAND2X1
XNAND2X1_22 NAND3X1_6/B NAND3X1_6/A gnd XNOR2X1_6/A vdd NAND2X1
XFILL_8_2 gnd vdd FILL
XFILL_10_7_0 gnd vdd FILL
XAOI21X1_261 INVX1_326/A AOI21X1_261/B INVX1_325/Y gnd NOR3X1_71/C vdd AOI21X1
XNAND3X1_434 INVX1_394/Y INVX1_393/A NAND3X1_434/C gnd AND2X2_141/B vdd NAND3X1
XINVX1_273 INVX1_273/A gnd INVX1_273/Y vdd INVX1
XDFFPOSX1_25 BUFX2_24/A CLKBUF1_43/Y NOR3X1_24/Y gnd vdd DFFPOSX1
XAOI21X1_1 AOI21X1_1/A AOI21X1_1/B NOR2X1_3/Y gnd OAI21X1_2/B vdd AOI21X1
XXOR2X1_68 NOR2X1_77/Y XOR2X1_54/A gnd XOR2X1_68/Y vdd XOR2X1
XNAND3X1_99 AOI21X1_72/C NAND3X1_99/B NOR3X1_35/Y gnd INVX1_74/A vdd NAND3X1
XOAI21X1_452 gnd NOR2X1_287/B INVX1_359/A gnd INVX2_68/A vdd OAI21X1
XNAND2X1_566 XNOR2X1_199/B NAND2X1_565/Y gnd NOR2X1_332/B vdd NAND2X1
XFILL_20_2_0 gnd vdd FILL
XOR2X2_151 OR2X2_151/A OR2X2_151/B gnd OR2X2_151/Y vdd OR2X2
XFILL_0_3_0 gnd vdd FILL
XAOI21X1_225 NAND2X1_372/A NAND2X1_372/B AOI21X1_225/C gnd OAI21X1_335/C vdd AOI21X1
XFILL_18_4_1 gnd vdd FILL
XNAND3X1_398 INVX1_344/A NAND2X1_480/B INVX2_67/Y gnd OAI21X1_442/B vdd NAND3X1
XAND2X2_168 AND2X2_159/B INVX2_74/A gnd AND2X2_168/Y vdd AND2X2
XINVX1_237 INVX1_237/A gnd INVX1_237/Y vdd INVX1
XOAI21X1_416 gnd NOR2X1_264/B INVX1_322/A gnd INVX1_325/A vdd OAI21X1
XNOR2X1_449 gnd gnd gnd NOR2X1_449/Y vdd NOR2X1
XNAND3X1_63 AOI21X1_48/C NAND3X1_63/B NOR3X1_31/Y gnd INVX1_52/A vdd NAND3X1
XXOR2X1_32 OR2X2_36/A gnd gnd XOR2X1_32/Y vdd XOR2X1
XOR2X2_115 gnd OR2X2_115/B gnd OR2X2_115/Y vdd OR2X2
XNAND2X1_530 NAND2X1_529/Y INVX1_392/Y gnd INVX1_393/A vdd NAND2X1
XAOI21X1_189 INVX2_53/Y XNOR2X1_131/A NAND2X1_288/Y gnd AOI21X1_189/Y vdd AOI21X1
XINVX1_83 INVX1_83/A gnd OR2X2_55/B vdd INVX1
XFILL_8_0_1 gnd vdd FILL
XNAND3X1_362 INVX1_289/Y INVX1_290/Y INVX1_291/Y gnd NAND3X1_362/Y vdd NAND3X1
XINVX1_201 INVX1_201/A gnd INVX1_201/Y vdd INVX1
XNOR2X1_413 NOR2X1_413/A NOR2X1_413/B gnd INVX1_539/A vdd NOR2X1
XOAI21X1_380 NOR3X1_68/A NOR3X1_68/C INVX2_64/A gnd NOR2X1_241/A vdd OAI21X1
XAND2X2_132 AND2X2_132/A NOR3X1_73/A gnd BUFX2_220/A vdd AND2X2
XNAND3X1_27 NAND3X1_26/C NAND3X1_26/A NOR3X1_27/Y gnd INVX1_30/A vdd NAND3X1
XNAND2X1_494 OAI21X1_450/Y NAND3X1_409/Y gnd XOR2X1_250/A vdd NAND2X1
XNAND3X1_326 INVX1_236/A NAND3X1_326/B NAND3X1_326/C gnd NAND2X1_372/A vdd NAND3X1
XAOI21X1_153 INVX2_44/Y XNOR2X1_104/A AOI21X1_153/C gnd NAND3X1_219/A vdd AOI21X1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_165 INVX1_165/A gnd INVX1_165/Y vdd INVX1
XFILL_17_7_0 gnd vdd FILL
XOAI21X1_344 gnd XOR2X1_183/Y INVX1_248/A gnd INVX1_250/A vdd OAI21X1
XNOR2X1_377 BUFX4_15/Y INVX2_80/Y gnd NOR2X1_377/Y vdd NOR2X1
XFILL_15_9_1 gnd vdd FILL
XNAND2X1_458 NAND2X1_458/A NAND3X1_384/B gnd BUFX2_215/A vdd NAND2X1
XAOI21X1_117 INVX2_35/Y XNOR2X1_77/A XNOR2X1_78/A gnd NAND3X1_165/A vdd AOI21X1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XNAND3X1_290 INVX2_57/Y NAND3X1_290/B NAND2X1_313/B gnd AOI21X1_199/B vdd NAND3X1
XAND2X2_69 gnd OR2X2_90/B gnd NOR3X1_48/C vdd AND2X2
XFILL_7_3_0 gnd vdd FILL
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XOAI21X1_308 BUFX2_179/A INVX1_214/A INVX1_215/Y gnd AOI21X1_212/A vdd OAI21X1
XFILL_25_4_1 gnd vdd FILL
XFILL_27_2_0 gnd vdd FILL
XFILL_5_5_1 gnd vdd FILL
XNAND2X1_422 INVX1_284/Y NOR2X1_240/Y gnd NAND2X1_423/B vdd NAND2X1
XNOR2X1_341 NOR2X1_341/A NOR3X1_83/Y gnd NOR2X1_341/Y vdd NOR2X1
XAND2X2_33 gnd OR2X2_42/B gnd NOR3X1_36/C vdd AND2X2
XNAND3X1_254 INVX2_51/Y NAND3X1_254/B NAND3X1_254/C gnd AOI21X1_175/B vdd NAND3X1
XBUFX2_255 OR2X2_52/A gnd BUFX2_255/Y vdd BUFX2
XINVX2_93 INVX2_93/A gnd INVX2_93/Y vdd INVX2
XOAI21X1_272 OAI21X1_267/A XNOR2X1_142/B OAI21X1_272/C gnd NAND2X1_313/B vdd OAI21X1
XNOR2X1_305 NOR2X1_305/A NOR3X1_77/Y gnd NOR2X1_305/Y vdd NOR2X1
XBUFX4_18 BUFX4_18/A gnd NOR3X1_3/C vdd BUFX4
XNAND2X1_386 INVX1_248/A NOR2X1_219/Y gnd NAND3X1_334/C vdd NAND2X1
XNAND3X1_218 INVX2_45/Y NAND3X1_218/B OAI21X1_204/Y gnd AOI21X1_151/B vdd NAND3X1
XBUFX2_219 BUFX2_219/A gnd BUFX2_219/Y vdd BUFX2
XXNOR2X1_257 gnd gnd gnd OR2X2_161/A vdd XNOR2X1
XNOR2X1_72 OR2X2_44/A OR2X2_44/B gnd NOR2X1_72/Y vdd NOR2X1
XOAI21X1_236 AND2X2_83/Y NOR2X1_152/Y INVX1_157/A gnd NAND3X1_247/C vdd OAI21X1
XINVX2_57 INVX2_57/A gnd INVX2_57/Y vdd INVX2
XNAND2X1_350 NAND2X1_350/A INVX1_218/A gnd XNOR2X1_152/B vdd NAND2X1
XNOR2X1_269 NOR2X1_269/A NOR3X1_71/Y gnd NOR2X1_269/Y vdd NOR2X1
XFILL_22_9_1 gnd vdd FILL
XFILL_24_7_0 gnd vdd FILL
XNOR2X1_36 INVX1_29/Y NOR2X1_36/B gnd NOR2X1_37/B vdd NOR2X1
XINVX1_598 INVX1_598/A gnd INVX1_598/Y vdd INVX1
XFILL_4_8_0 gnd vdd FILL
XBUFX2_183 BUFX2_183/A gnd BUFX2_183/Y vdd BUFX2
XXNOR2X1_221 bloque_bytes[26] INVX1_531/A gnd XNOR2X1_221/Y vdd XNOR2X1
XNAND3X1_182 INVX2_39/Y NAND3X1_182/B OAI21X1_170/Y gnd AOI21X1_127/B vdd NAND3X1
XNAND3X1_1 NAND2X1_3/A NAND2X1_3/B NOR2X1_9/Y gnd NOR2X1_10/B vdd NAND3X1
XOAI21X1_200 AND2X2_70/Y NOR2X1_130/Y INVX1_134/Y gnd AOI21X1_144/A vdd OAI21X1
XNOR2X1_233 NOR2X1_233/A NOR3X1_65/Y gnd NOR2X1_233/Y vdd NOR2X1
XINVX2_21 INVX2_21/A gnd INVX2_21/Y vdd INVX2
XNAND2X1_314 AND2X2_96/B AND2X2_96/A gnd OAI21X1_273/B vdd NAND2X1
XFILL_34_2_0 gnd vdd FILL
XBUFX2_147 gnd gnd BUFX2_147/Y vdd BUFX2
XCLKBUF1_24 BUFX4_3/Y gnd CLKBUF1_24/Y vdd CLKBUF1
XINVX1_562 bloque_bytes[3] gnd INVX1_562/Y vdd INVX1
XNAND3X1_146 INVX2_33/Y NAND3X1_146/B NAND3X1_146/C gnd AOI21X1_103/B vdd NAND3X1
XFILL_32_4_1 gnd vdd FILL
XOR2X2_4 gnd OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XXNOR2X1_185 NOR2X1_293/Y NOR2X1_292/Y gnd XOR2X1_256/A vdd XNOR2X1
XNOR2X1_197 NOR2X1_197/A NOR3X1_59/Y gnd NOR2X1_197/Y vdd NOR2X1
XNAND2X1_278 AOI21X1_173/A AOI21X1_173/B gnd INVX2_52/A vdd NAND2X1
XOAI21X1_164 NOR3X1_44/Y NOR2X1_113/A NAND3X1_170/B gnd NAND2X1_196/B vdd OAI21X1
XDFFPOSX1_344 INVX1_410/A CLKBUF1_19/Y NAND2X1_689/Y gnd vdd DFFPOSX1
XNOR3X1_77 NOR3X1_77/A INVX1_380/A NOR3X1_77/C gnd NOR3X1_77/Y vdd NOR3X1
XNAND3X1_110 INVX2_27/Y AOI21X1_77/Y NAND3X1_110/C gnd AOI21X1_79/B vdd NAND3X1
XINVX1_526 INVX1_526/A gnd INVX1_526/Y vdd INVX1
XBUFX2_111 gnd gnd BUFX2_111/Y vdd BUFX2
XXNOR2X1_149 NOR2X1_185/Y NOR2X1_184/Y gnd XOR2X1_175/A vdd XNOR2X1
XXNOR2X1_71 XNOR2X1_71/A AND2X2_48/Y gnd XOR2X1_86/A vdd XNOR2X1
XOAI21X1_128 NOR3X1_40/Y NOR2X1_93/A NOR3X1_39/Y gnd NAND2X1_157/B vdd OAI21X1
XNOR2X1_161 NOR2X1_161/A INVX2_54/A gnd XOR2X1_150/B vdd NOR2X1
XNAND2X1_242 OR2X2_95/B OR2X2_95/A gnd NAND2X1_243/A vdd NAND2X1
XNOR3X1_41 INVX1_99/Y NOR3X1_41/B NOR3X1_41/C gnd NOR3X1_41/Y vdd NOR3X1
XDFFPOSX1_308 INVX1_322/A CLKBUF1_39/Y INVX1_554/Y gnd vdd DFFPOSX1
XINVX1_490 INVX1_490/A gnd INVX1_490/Y vdd INVX1
XXNOR2X1_113 NAND2X1_248/B INVX2_47/Y gnd AND2X2_89/A vdd XNOR2X1
XFILL_21_2 gnd vdd FILL
XFILL_31_7_0 gnd vdd FILL
XXOR2X1_305 AND2X2_188/A BUFX2_243/A gnd XOR2X1_305/Y vdd XOR2X1
XXNOR2X1_35 OAI21X1_69/A AND2X2_24/Y gnd XOR2X1_46/A vdd XNOR2X1
XNOR2X1_125 NOR2X1_125/A INVX1_126/Y gnd NOR2X1_125/Y vdd NOR2X1
XFILL_29_9_1 gnd vdd FILL
XNAND2X1_206 OR2X2_80/B OR2X2_80/A gnd NAND2X1_206/Y vdd NAND2X1
XDFFPOSX1_272 INVX1_239/A CLKBUF1_33/Y INVX1_534/Y gnd vdd DFFPOSX1
XOR2X2_93 OR2X2_93/A OR2X2_93/B gnd OR2X2_93/Y vdd OR2X2
XOAI21X1_633 INVX1_586/Y INVX1_587/A INVX1_588/A gnd OAI21X1_633/Y vdd OAI21X1
XINVX1_454 INVX1_454/A gnd INVX1_454/Y vdd INVX1
XXOR2X1_269 XOR2X1_269/A XOR2X1_269/B gnd XOR2X1_275/A vdd XOR2X1
XXOR2X1_9 XOR2X1_9/A vdd gnd XOR2X1_9/Y vdd XOR2X1
XNAND2X1_170 INVX2_34/A AND2X2_48/Y gnd OAI21X1_140/B vdd NAND2X1
XAOI21X1_68 INVX2_24/Y INVX1_63/Y NOR2X1_61/A gnd AOI21X1_68/Y vdd AOI21X1
XDFFPOSX1_236 INVX1_166/A CLKBUF1_47/Y INVX1_513/A gnd vdd DFFPOSX1
XMUX2X1_15 BUFX2_15/A XOR2X1_1/B BUFX4_8/Y gnd MUX2X1_15/Y vdd MUX2X1
XOAI21X1_597 bloque_bytes[74] INVX2_85/Y OAI21X1_597/C gnd OR2X2_139/A vdd OAI21X1
XOR2X2_57 gnd OR2X2_57/B gnd OR2X2_57/Y vdd OR2X2
XINVX1_418 INVX1_418/A gnd INVX1_418/Y vdd INVX1
XXOR2X1_233 XOR2X1_233/A XOR2X1_233/B gnd XOR2X1_233/Y vdd XOR2X1
XNAND2X1_711 gnd gnd gnd NAND3X1_541/B vdd NAND2X1
XBUFX2_71 gnd gnd BUFX2_71/Y vdd BUFX2
XNAND3X1_543 INVX1_594/Y NAND3X1_545/B OR2X2_159/Y gnd NAND3X1_544/C vdd NAND3X1
XNAND2X1_134 INVX2_29/Y AOI21X1_93/B gnd XNOR2X1_60/B vdd NAND2X1
XAOI21X1_370 AOI21X1_370/A OR2X2_131/Y INVX1_501/A gnd AOI21X1_370/Y vdd AOI21X1
XAOI21X1_32 INVX2_15/Y INVX1_30/Y NOR2X1_31/A gnd AOI21X1_32/Y vdd AOI21X1
XOR2X2_21 OR2X2_21/A OR2X2_21/B gnd OR2X2_21/Y vdd OR2X2
XFILL_13_2_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XDFFPOSX1_200 INVX1_116/A CLKBUF1_36/Y bloque_bytes[14] gnd vdd DFFPOSX1
XINVX1_382 INVX1_382/A gnd INVX1_382/Y vdd INVX1
XXOR2X1_197 XOR2X1_197/A XOR2X1_197/B gnd XOR2X1_197/Y vdd XOR2X1
XNAND2X1_675 INVX1_571/Y INVX1_550/A gnd NAND2X1_675/Y vdd NAND2X1
XOAI21X1_561 BUFX2_237/A NOR2X1_355/B INVX1_467/A gnd OAI21X1_561/Y vdd OAI21X1
XAOI21X1_334 NOR2X1_400/Y INVX2_83/A BUFX4_16/Y gnd AND2X2_170/B vdd AOI21X1
XBUFX2_35 gnd gnd BUFX2_35/Y vdd BUFX2
XNAND2X1_95 NAND2X1_95/A NAND2X1_95/B gnd XOR2X1_49/A vdd NAND2X1
XOAI21X1_80 OAI21X1_85/A OAI21X1_85/B INVX1_63/A gnd XOR2X1_50/A vdd OAI21X1
XNAND3X1_507 NAND2X1_654/A NAND3X1_507/B AOI21X1_374/Y gnd XNOR2X1_242/A vdd NAND3X1
XDFFPOSX1_98 INVX1_4/A CLKBUF1_41/Y INVX1_578/Y gnd vdd DFFPOSX1
XINVX2_8 target[7] gnd INVX2_8/Y vdd INVX2
XDFFPOSX1_164 INVX1_67/A CLKBUF1_47/Y bloque_bytes[42] gnd vdd DFFPOSX1
XFILL_36_9_1 gnd vdd FILL
XINVX1_346 INVX1_346/A gnd INVX1_346/Y vdd INVX1
XOAI21X1_525 NOR2X1_329/A NOR3X1_81/Y OAI21X1_525/C gnd OAI21X1_525/Y vdd OAI21X1
XXOR2X1_161 BUFX2_174/A XOR2X1_161/B gnd XOR2X1_161/Y vdd XOR2X1
XNAND2X1_639 AOI21X1_370/A OR2X2_131/Y gnd NAND2X1_639/Y vdd NAND2X1
XNAND2X1_59 gnd OR2X2_17/B gnd NAND3X1_41/B vdd NAND2X1
XAOI21X1_298 INVX1_413/Y NAND3X1_447/C INVX1_412/A gnd OAI21X1_507/A vdd AOI21X1
XNAND3X1_471 INVX1_437/Y NAND3X1_464/Y NOR3X1_84/Y gnd AOI21X1_312/B vdd NAND3X1
XDFFPOSX1_128 INVX1_17/A CLKBUF1_5/Y bloque_bytes[86] gnd vdd DFFPOSX1
XOAI21X1_44 NOR3X1_30/C NOR3X1_30/B INVX1_34/Y gnd NAND3X1_44/A vdd OAI21X1
XDFFPOSX1_62 INVX1_473/A CLKBUF1_38/Y NOR2X1_385/Y gnd vdd DFFPOSX1
XXOR2X1_125 BUFX2_166/A gnd gnd AND2X2_82/B vdd XOR2X1
XOAI21X1_489 gnd NOR2X1_310/B INVX1_396/A gnd OAI21X1_489/Y vdd OAI21X1
XINVX1_310 INVX1_310/A gnd INVX1_310/Y vdd INVX1
XFILL_12_5_0 gnd vdd FILL
XNOR2X1_6 target[5] INVX2_1/Y gnd NOR2X1_6/Y vdd NOR2X1
XNAND2X1_603 INVX1_467/Y NOR2X1_355/Y gnd NAND2X1_603/Y vdd NAND2X1
XNAND2X1_23 gnd OR2X2_2/B gnd NAND3X1_7/B vdd NAND2X1
XFILL_10_7_1 gnd vdd FILL
XDFFPOSX1_26 INVX1_507/A CLKBUF1_20/Y NOR2X1_358/Y gnd vdd DFFPOSX1
XAOI21X1_262 OAI21X1_427/Y NAND2X1_468/Y INVX2_66/A gnd AOI21X1_263/B vdd AOI21X1
XNAND3X1_435 INVX1_392/Y INVX1_395/Y AND2X2_141/A gnd NAND2X1_532/B vdd NAND3X1
XINVX1_274 INVX1_274/A gnd INVX1_274/Y vdd INVX1
XOAI21X1_453 NOR3X1_76/C INVX2_68/Y NOR3X1_76/A gnd AND2X2_136/A vdd OAI21X1
XAOI21X1_2 NAND2X1_6/Y NOR2X1_5/Y NOR2X1_4/Y gnd AOI21X1_2/Y vdd AOI21X1
XXOR2X1_69 XOR2X1_69/A XOR2X1_71/A gnd XOR2X1_69/Y vdd XOR2X1
XFILL_22_0_0 gnd vdd FILL
XNAND2X1_567 INVX1_428/Y NOR2X1_332/B gnd NAND2X1_567/Y vdd NAND2X1
XFILL_2_1_0 gnd vdd FILL
XAOI21X1_226 INVX1_242/Y AOI21X1_226/B INVX1_241/A gnd OAI21X1_336/A vdd AOI21X1
XFILL_20_2_1 gnd vdd FILL
XOR2X2_152 OR2X2_137/Y OR2X2_152/B gnd OR2X2_152/Y vdd OR2X2
XFILL_0_3_1 gnd vdd FILL
XNAND3X1_399 INVX1_344/A OAI21X1_438/Y NAND3X1_399/C gnd NAND3X1_399/Y vdd NAND3X1
XAND2X2_169 INVX1_474/A AND2X2_169/B gnd AND2X2_169/Y vdd AND2X2
XINVX1_238 INVX1_238/A gnd INVX1_238/Y vdd INVX1
XOAI21X1_417 NOR3X1_71/A NOR3X1_71/B OAI21X1_423/B gnd NOR2X1_266/A vdd OAI21X1
XNAND3X1_64 INVX1_46/A NAND3X1_64/B OR2X2_27/Y gnd NAND3X1_64/Y vdd NAND3X1
XNOR2X1_450 NOR2X1_450/A NOR3X1_98/Y gnd NOR2X1_450/Y vdd NOR2X1
XXOR2X1_33 OR2X2_37/A gnd gnd OR2X2_33/B vdd XOR2X1
XOR2X2_116 AND2X2_89/A AND2X2_89/B gnd OR2X2_116/Y vdd OR2X2
XNAND2X1_531 NAND2X1_531/A AOI22X1_18/C gnd AOI21X1_289/C vdd NAND2X1
XAOI21X1_190 AOI21X1_190/A NAND3X1_273/Y AOI21X1_190/C gnd OAI21X1_261/A vdd AOI21X1
XNAND3X1_363 INVX1_291/A INVX1_289/Y INVX1_290/Y gnd NAND3X1_363/Y vdd NAND3X1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XNAND3X1_28 INVX1_24/A NAND3X1_28/B OR2X2_11/Y gnd AOI21X1_24/B vdd NAND3X1
XINVX1_202 INVX1_202/A gnd INVX1_202/Y vdd INVX1
XNOR2X1_414 NOR2X1_414/A INVX1_576/A gnd INVX1_540/A vdd NOR2X1
XOAI21X1_381 gnd XOR2X1_201/Y INVX1_286/Y gnd NAND3X1_360/B vdd OAI21X1
XAND2X2_133 AND2X2_133/A AND2X2_133/B gnd AND2X2_133/Y vdd AND2X2
XNAND2X1_495 INVX1_358/Y NOR2X1_286/Y gnd NAND3X1_410/B vdd NAND2X1
XNAND3X1_327 AOI22X1_10/B INVX1_238/A INVX1_236/Y gnd NAND2X1_372/B vdd NAND3X1
XAOI21X1_154 AOI21X1_152/Y NAND3X1_219/Y AOI21X1_154/C gnd OAI21X1_210/A vdd AOI21X1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_166 INVX1_166/A gnd INVX1_166/Y vdd INVX1
XFILL_17_7_1 gnd vdd FILL
XOAI21X1_345 INVX1_251/A INVX1_252/A INVX1_253/A gnd INVX1_255/A vdd OAI21X1
XFILL_19_5_0 gnd vdd FILL
XNOR2X1_378 BUFX4_17/Y INVX2_81/Y gnd NOR2X1_378/Y vdd NOR2X1
XFILL_12_1 gnd vdd FILL
XNAND2X1_459 INVX1_321/Y AND2X2_127/A gnd NAND3X1_384/C vdd NAND2X1
XAOI21X1_118 AOI21X1_118/A AOI21X1_118/B NAND2X1_189/Y gnd OAI21X1_159/A vdd AOI21X1
XAND2X2_70 gnd OR2X2_91/B gnd AND2X2_70/Y vdd AND2X2
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XNAND3X1_291 AOI21X1_201/Y XNOR2X1_142/A XOR2X1_160/B gnd AOI21X1_202/B vdd NAND3X1
XFILL_27_2_1 gnd vdd FILL
XFILL_29_0_0 gnd vdd FILL
XFILL_7_3_1 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XINVX1_130 OR2X2_88/Y gnd INVX1_130/Y vdd INVX1
XOAI21X1_309 NOR3X1_59/C OAI21X1_309/B INVX1_218/A gnd NOR2X1_197/A vdd OAI21X1
XNOR2X1_342 BUFX2_232/A NOR2X1_342/B gnd NOR2X1_342/Y vdd NOR2X1
XNAND2X1_423 INVX1_287/A NAND2X1_423/B gnd NOR3X1_67/B vdd NAND2X1
XBUFX2_256 OR2X2_53/A gnd BUFX2_256/Y vdd BUFX2
XAND2X2_34 gnd OR2X2_43/B gnd AND2X2_34/Y vdd AND2X2
XNAND3X1_255 AOI21X1_177/Y XNOR2X1_124/A XOR2X1_140/B gnd AOI21X1_178/B vdd NAND3X1
XINVX2_94 INVX2_94/A gnd INVX2_94/Y vdd INVX2
XOAI21X1_273 XNOR2X1_143/A OAI21X1_273/B AND2X2_96/B gnd XNOR2X1_144/A vdd OAI21X1
XNAND2X1_387 INVX1_248/Y NOR2X1_219/Y gnd NAND2X1_387/Y vdd NAND2X1
XFILL_34_1 gnd vdd FILL
XNOR2X1_306 BUFX2_220/A NOR2X1_306/B gnd NOR2X1_306/Y vdd NOR2X1
XBUFX4_19 BUFX4_18/A gnd NOR3X1_9/C vdd BUFX4
XNAND3X1_219 NAND3X1_219/A XNOR2X1_106/A XOR2X1_120/B gnd NAND3X1_219/Y vdd NAND3X1
XBUFX2_220 BUFX2_220/A gnd BUFX2_220/Y vdd BUFX2
XXNOR2X1_258 XOR2X1_318/Y gnd gnd XNOR2X1_258/Y vdd XNOR2X1
XNOR2X1_73 NOR2X1_73/A NOR2X1_73/B gnd NOR2X1_73/Y vdd NOR2X1
XOAI21X1_237 AND2X2_83/Y NOR2X1_152/Y INVX1_157/Y gnd NAND3X1_251/A vdd OAI21X1
XNAND2X1_351 INVX1_216/A NOR2X1_198/Y gnd NAND3X1_313/C vdd NAND2X1
XINVX2_58 INVX2_58/A gnd INVX2_58/Y vdd INVX2
XFILL_26_5_0 gnd vdd FILL
XNOR2X1_270 BUFX2_208/A XOR2X1_221/Y gnd NOR2X1_270/Y vdd NOR2X1
XINVX1_599 INVX1_599/A gnd INVX1_599/Y vdd INVX1
XFILL_6_6_0 gnd vdd FILL
XFILL_24_7_1 gnd vdd FILL
XNAND3X1_183 AOI21X1_129/Y XNOR2X1_88/A XOR2X1_100/B gnd AOI21X1_130/B vdd NAND3X1
XNOR2X1_37 NOR2X1_37/A NOR2X1_37/B gnd XOR2X1_28/A vdd NOR2X1
XFILL_4_8_1 gnd vdd FILL
XBUFX2_184 BUFX2_184/A gnd BUFX2_184/Y vdd BUFX2
XXNOR2X1_222 bloque_bytes[27] INVX1_503/A gnd NAND3X1_506/B vdd XNOR2X1
XNAND3X1_2 NAND3X1_2/A NAND3X1_2/B NAND3X1_2/C gnd NAND3X1_2/Y vdd NAND3X1
XINVX2_22 INVX2_22/A gnd INVX2_22/Y vdd INVX2
XNOR2X1_234 BUFX2_192/A XOR2X1_194/Y gnd NOR2X1_234/Y vdd NOR2X1
XOAI21X1_201 AND2X2_70/Y NOR2X1_130/Y INVX1_134/A gnd AOI21X1_145/A vdd OAI21X1
XFILL_36_0_0 gnd vdd FILL
XNAND2X1_315 OR2X2_125/A OR2X2_125/B gnd NAND3X1_286/B vdd NAND2X1
XFILL_34_2_1 gnd vdd FILL
XCLKBUF1_25 BUFX4_7/Y gnd CLKBUF1_25/Y vdd CLKBUF1
XOR2X2_5 vdd OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XBUFX2_148 gnd gnd BUFX2_148/Y vdd BUFX2
XNAND3X1_147 NAND3X1_147/A XNOR2X1_70/A NOR2X1_91/Y gnd AOI21X1_106/B vdd NAND3X1
XINVX1_563 INVX1_563/A gnd INVX1_563/Y vdd INVX1
XOAI21X1_165 OAI21X1_165/A XNOR2X1_88/B INVX1_118/A gnd XOR2X1_100/A vdd OAI21X1
XXNOR2X1_186 NOR2X1_297/Y XNOR2X1_186/B gnd XNOR2X1_186/Y vdd XNOR2X1
XNOR2X1_198 BUFX2_180/A NOR2X1_198/B gnd NOR2X1_198/Y vdd NOR2X1
XNAND2X1_279 NAND3X1_253/A OR2X2_112/B gnd OR2X2_110/A vdd NAND2X1
XDFFPOSX1_345 XNOR2X1_194/B CLKBUF1_22/Y NAND2X1_690/Y gnd vdd DFFPOSX1
XNOR3X1_78 NOR3X1_78/A INVX2_69/Y NOR3X1_78/C gnd NOR3X1_78/Y vdd NOR3X1
XINVX1_527 bloque_bytes[63] gnd INVX1_527/Y vdd INVX1
XNAND3X1_111 AOI21X1_81/Y XNOR2X1_52/A NOR2X1_71/Y gnd AOI21X1_82/B vdd NAND3X1
XXNOR2X1_150 NOR2X1_189/Y XNOR2X1_150/B gnd XNOR2X1_151/A vdd XNOR2X1
XBUFX2_112 gnd gnd BUFX2_112/Y vdd BUFX2
XNOR2X1_162 AND2X2_89/A AND2X2_89/B gnd NOR2X1_162/Y vdd NOR2X1
XXNOR2X1_72 XNOR2X1_72/A INVX2_34/Y gnd XOR2X1_87/A vdd XNOR2X1
XOAI21X1_129 AND2X2_45/Y NOR2X1_89/Y INVX1_89/Y gnd OAI21X1_129/Y vdd OAI21X1
XNAND2X1_243 NAND2X1_243/A OR2X2_95/Y gnd OR2X2_96/A vdd NAND2X1
XNOR3X1_42 NOR3X1_42/A NOR3X1_42/B NOR3X1_42/C gnd NOR3X1_42/Y vdd NOR3X1
XINVX1_491 INVX1_491/A gnd INVX1_491/Y vdd INVX1
XDFFPOSX1_309 INVX1_324/A CLKBUF1_39/Y OR2X2_137/Y gnd vdd DFFPOSX1
XXNOR2X1_36 XNOR2X1_36/A INVX2_22/Y gnd XOR2X1_47/A vdd XNOR2X1
XXNOR2X1_114 XNOR2X1_114/A XNOR2X1_114/B gnd OR2X2_117/A vdd XNOR2X1
XFILL_33_5_0 gnd vdd FILL
XFILL_31_7_1 gnd vdd FILL
XXOR2X1_306 XOR2X1_306/A BUFX2_245/A gnd XOR2X1_306/Y vdd XOR2X1
XNOR2X1_126 INVX1_128/Y NOR2X1_126/B gnd NOR2X1_127/B vdd NOR2X1
XNAND2X1_207 NAND2X1_206/Y OR2X2_80/Y gnd INVX1_117/A vdd NAND2X1
XDFFPOSX1_273 XNOR2X1_158/B CLKBUF1_44/Y NAND2X1_656/Y gnd vdd DFFPOSX1
XOR2X2_94 OR2X2_94/A OR2X2_94/B gnd OR2X2_94/Y vdd OR2X2
XINVX1_455 INVX1_455/A gnd INVX1_455/Y vdd INVX1
XOAI21X1_634 NOR2X1_444/B XOR2X1_296/Y INVX1_589/A gnd NAND2X1_703/A vdd OAI21X1
XXOR2X1_270 BUFX2_231/A gnd gnd XOR2X1_270/Y vdd XOR2X1
XNAND2X1_171 NAND3X1_148/Y OAI21X1_143/Y gnd XOR2X1_89/A vdd NAND2X1
XAOI21X1_69 INVX2_23/Y AOI21X1_69/B NAND2X1_98/Y gnd NAND3X1_93/A vdd AOI21X1
XDFFPOSX1_237 INVX1_167/A CLKBUF1_47/Y INVX1_516/A gnd vdd DFFPOSX1
XMUX2X1_16 BUFX2_16/A NOR2X1_1/B BUFX4_9/Y gnd MUX2X1_16/Y vdd MUX2X1
XOAI21X1_598 bloque_bytes[77] INVX2_86/Y AOI21X1_359/Y gnd XNOR2X1_234/A vdd OAI21X1
XOR2X2_58 gnd OR2X2_58/B gnd OR2X2_58/Y vdd OR2X2
XXOR2X1_234 BUFX2_215/A gnd gnd XOR2X1_234/Y vdd XOR2X1
XINVX1_419 INVX1_419/A gnd INVX1_419/Y vdd INVX1
XNAND2X1_712 INVX2_93/Y NAND2X1_712/B gnd XNOR2X1_255/A vdd NAND2X1
XBUFX2_72 gnd gnd BUFX2_72/Y vdd BUFX2
XNAND3X1_544 NAND3X1_544/A NAND3X1_544/B NAND3X1_544/C gnd AOI21X1_400/A vdd NAND3X1
XNAND2X1_135 gnd OR2X2_49/B gnd NAND3X1_113/B vdd NAND2X1
XFILL_15_0_1 gnd vdd FILL
XAOI21X1_371 AOI21X1_371/A OR2X2_132/Y INVX1_502/A gnd AOI21X1_371/Y vdd AOI21X1
XAOI21X1_33 INVX2_14/Y XNOR2X1_14/A XNOR2X1_15/A gnd NAND3X1_39/A vdd AOI21X1
XOR2X2_22 OR2X2_22/A OR2X2_22/B gnd INVX1_38/A vdd OR2X2
XDFFPOSX1_201 XOR2X1_101/B CLKBUF1_9/Y bloque_bytes[15] gnd vdd DFFPOSX1
XINVX1_383 INVX1_383/A gnd INVX1_383/Y vdd INVX1
XOAI21X1_562 AOI21X1_320/Y INVX1_470/A INVX1_469/Y gnd AND2X2_157/A vdd OAI21X1
XBUFX2_36 gnd gnd BUFX2_36/Y vdd BUFX2
XNAND2X1_676 INVX1_572/Y INVX1_551/A gnd NAND2X1_676/Y vdd NAND2X1
XXOR2X1_198 INVX1_289/A gnd gnd XOR2X1_198/Y vdd XOR2X1
XAOI21X1_335 NOR2X1_400/Y INVX2_83/A AND2X2_165/B gnd NOR2X1_401/A vdd AOI21X1
XOAI21X1_81 AND2X2_28/Y NOR2X1_60/Y INVX1_57/Y gnd NAND3X1_85/A vdd OAI21X1
XNAND2X1_96 INVX2_23/Y AOI21X1_69/B gnd NAND3X1_78/C vdd NAND2X1
XDFFPOSX1_165 INVX1_68/A CLKBUF1_44/Y bloque_bytes[43] gnd vdd DFFPOSX1
XNAND3X1_508 INVX1_549/Y XNOR2X1_224/Y AOI21X1_378/Y gnd NAND3X1_508/Y vdd NAND3X1
XINVX2_9 target[6] gnd INVX2_9/Y vdd INVX2
XDFFPOSX1_99 INVX1_3/A CLKBUF1_41/Y NOR2X1_436/Y gnd vdd DFFPOSX1
XXOR2X1_162 BUFX2_179/A gnd gnd XOR2X1_162/Y vdd XOR2X1
XINVX1_347 INVX1_347/A gnd INVX1_347/Y vdd INVX1
XOAI21X1_526 AOI21X1_306/Y INVX1_430/A INVX1_433/A gnd OAI21X1_526/Y vdd OAI21X1
XNAND2X1_640 INVX1_501/Y NAND2X1_639/Y gnd OR2X2_150/B vdd NAND2X1
XOAI21X1_45 NOR2X1_43/B NOR2X1_43/A NAND3X1_42/A gnd NAND2X1_63/B vdd OAI21X1
XNAND2X1_60 NAND3X1_42/B NAND3X1_42/A gnd NAND2X1_60/Y vdd NAND2X1
XNAND3X1_472 INVX1_440/A OAI21X1_536/Y NAND3X1_467/Y gnd NAND2X1_588/A vdd NAND3X1
XAOI21X1_299 INVX1_426/A NAND3X1_455/B INVX1_421/Y gnd NOR2X1_328/B vdd AOI21X1
XDFFPOSX1_129 XOR2X1_11/B CLKBUF1_25/Y bloque_bytes[87] gnd vdd DFFPOSX1
XDFFPOSX1_63 INVX1_474/A CLKBUF1_38/Y DFFPOSX1_63/D gnd vdd DFFPOSX1
XINVX1_311 INVX1_311/A gnd INVX1_311/Y vdd INVX1
XFILL_14_3_0 gnd vdd FILL
XXOR2X1_126 XOR2X1_126/A AND2X2_77/A gnd OR2X2_108/B vdd XOR2X1
XOAI21X1_490 gnd NOR2X1_311/B INVX1_397/A gnd INVX2_70/A vdd OAI21X1
XNAND2X1_604 OAI21X1_561/Y NAND2X1_603/Y gnd NOR2X1_356/B vdd NAND2X1
XFILL_12_5_1 gnd vdd FILL
XNOR2X1_7 XOR2X1_1/B INVX2_9/Y gnd NOR2X1_7/Y vdd NOR2X1
XNAND2X1_24 NAND3X1_8/Y OAI21X1_9/Y gnd XNOR2X1_7/A vdd NAND2X1
XDFFPOSX1_27 INVX1_510/A CLKBUF1_20/Y AND2X2_158/Y gnd vdd DFFPOSX1
XAOI21X1_263 NAND3X1_386/Y AOI21X1_263/B INVX1_332/Y gnd AOI21X1_264/A vdd AOI21X1
XNAND3X1_436 INVX2_70/A NAND2X1_534/B NAND3X1_436/C gnd NOR3X1_79/A vdd NAND3X1
XINVX1_275 INVX1_275/A gnd INVX1_275/Y vdd INVX1
XOAI21X1_454 gnd XOR2X1_236/Y INVX1_360/A gnd INVX1_363/A vdd OAI21X1
XAOI21X1_3 INVX1_2/Y INVX1_1/A XOR2X1_1/Y gnd AOI21X1_3/Y vdd AOI21X1
XXOR2X1_70 XOR2X1_70/A NOR2X1_81/Y gnd XOR2X1_75/A vdd XOR2X1
XFILL_22_0_1 gnd vdd FILL
XOR2X2_153 OR2X2_138/Y OR2X2_153/B gnd OR2X2_153/Y vdd OR2X2
XNAND2X1_568 NAND2X1_567/Y INVX1_430/Y gnd INVX1_431/A vdd NAND2X1
XFILL_2_1_1 gnd vdd FILL
XAOI21X1_227 INVX1_255/A NAND3X1_336/Y INVX1_250/Y gnd NOR2X1_220/B vdd AOI21X1
XNAND3X1_400 INVX1_345/A NAND2X1_482/Y INVX1_344/Y gnd INVX1_351/A vdd NAND3X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XNOR2X1_451 gnd gnd gnd NOR2X1_451/Y vdd NOR2X1
XXOR2X1_34 BUFX2_249/A gnd gnd OR2X2_34/B vdd XOR2X1
XINVX1_239 INVX1_239/A gnd INVX1_239/Y vdd INVX1
XAND2X2_170 AND2X2_170/A AND2X2_170/B gnd AND2X2_170/Y vdd AND2X2
XOAI21X1_418 NOR3X1_72/A NOR3X1_72/C INVX2_66/A gnd NOR2X1_265/A vdd OAI21X1
XNAND3X1_65 INVX1_46/Y NAND3X1_64/B OR2X2_27/Y gnd NAND3X1_65/Y vdd NAND3X1
XOR2X2_117 OR2X2_117/A OR2X2_117/B gnd OR2X2_117/Y vdd OR2X2
XNAND2X1_532 NAND2X1_532/A NAND2X1_532/B gnd XOR2X1_268/A vdd NAND2X1
XAOI21X1_191 AOI21X1_191/A OR2X2_122/Y INVX1_177/A gnd NOR2X1_173/A vdd AOI21X1
XNAND3X1_364 INVX1_293/A NAND3X1_362/Y INVX1_288/Y gnd AOI22X1_13/C vdd NAND3X1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XFILL_11_8_0 gnd vdd FILL
XINVX1_203 INVX1_203/A gnd INVX1_203/Y vdd INVX1
XOAI21X1_382 gnd XOR2X1_201/Y INVX1_286/A gnd INVX1_288/A vdd OAI21X1
XNAND3X1_29 INVX1_24/Y NAND3X1_28/B OR2X2_11/Y gnd AOI21X1_25/B vdd NAND3X1
XNOR2X1_415 XOR2X1_303/Y INVX1_577/A gnd INVX1_541/A vdd NOR2X1
XAND2X2_134 NOR2X1_286/Y INVX1_358/Y gnd NOR3X1_76/A vdd AND2X2
XNAND2X1_496 NAND2X1_496/A NAND3X1_410/B gnd BUFX2_223/A vdd NAND2X1
XAOI21X1_155 AOI21X1_155/A OR2X2_98/Y INVX1_144/A gnd NOR2X1_143/A vdd AOI21X1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XNAND3X1_328 INVX1_228/Y AOI21X1_223/A NOR3X1_62/Y gnd AOI21X1_224/B vdd NAND3X1
XFILL_19_5_1 gnd vdd FILL
XFILL_21_3_0 gnd vdd FILL
XFILL_1_4_0 gnd vdd FILL
XINVX1_167 INVX1_167/A gnd INVX1_167/Y vdd INVX1
XOAI21X1_346 INVX1_251/A INVX1_252/A INVX1_253/Y gnd AOI21X1_228/A vdd OAI21X1
XNOR2X1_379 BUFX4_17/Y NOR3X1_95/A gnd NOR2X1_379/Y vdd NOR2X1
XFILL_12_2 gnd vdd FILL
XNAND2X1_460 INVX1_322/Y NOR2X1_264/Y gnd NAND2X1_460/Y vdd NAND2X1
XNAND3X1_292 INVX1_185/A INVX1_186/A NAND3X1_292/C gnd NAND2X1_323/A vdd NAND3X1
XAND2X2_71 OR2X2_92/A OR2X2_92/B gnd AND2X2_71/Y vdd AND2X2
XAOI21X1_119 NAND3X1_169/B OR2X2_74/Y INVX1_111/A gnd NOR2X1_113/A vdd AOI21X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XFILL_29_0_1 gnd vdd FILL
XINVX1_131 INVX1_131/A gnd INVX1_131/Y vdd INVX1
XOAI21X1_310 NOR2X1_197/Y NOR2X1_196/B AOI22X1_9/C gnd XOR2X1_179/A vdd OAI21X1
XNOR2X1_343 BUFX2_233/A NOR2X1_343/B gnd NOR2X1_343/Y vdd NOR2X1
XNAND2X1_424 INVX1_286/A NOR2X1_243/Y gnd NAND2X1_424/Y vdd NAND2X1
XBUFX2_257 XOR2X1_54/A gnd BUFX2_257/Y vdd BUFX2
XAND2X2_35 OR2X2_44/A OR2X2_44/B gnd AND2X2_35/Y vdd AND2X2
XNAND3X1_256 INVX1_163/A INVX1_164/A NAND3X1_256/C gnd NAND2X1_285/A vdd NAND3X1
XOAI21X1_274 AND2X2_97/Y NOR2X1_174/Y INVX1_180/A gnd NAND3X1_287/B vdd OAI21X1
XBUFX4_20 BUFX4_18/A gnd BUFX4_20/Y vdd BUFX4
XFILL_18_8_0 gnd vdd FILL
XNAND2X1_388 NAND3X1_334/Y INVX1_256/A gnd NAND2X1_388/Y vdd NAND2X1
XNOR2X1_307 BUFX2_221/A XOR2X1_249/Y gnd NOR2X1_307/Y vdd NOR2X1
XXNOR2X1_259 XNOR2X1_258/Y OR2X2_161/Y gnd INVX1_600/A vdd XNOR2X1
XNOR2X1_74 OR2X2_45/A OR2X2_45/B gnd NOR2X1_74/Y vdd NOR2X1
XNAND3X1_220 OR2X2_96/Y INVX1_142/A OAI21X1_210/Y gnd NAND2X1_247/A vdd NAND3X1
XBUFX2_221 BUFX2_221/A gnd BUFX2_221/Y vdd BUFX2
XOAI21X1_238 OAI21X1_233/A NAND3X1_240/Y OAI21X1_238/C gnd NAND3X1_254/C vdd OAI21X1
XNOR2X1_271 BUFX2_209/A NOR2X1_271/B gnd NOR2X1_271/Y vdd NOR2X1
XFILL_28_3_0 gnd vdd FILL
XFILL_8_4_0 gnd vdd FILL
XINVX2_59 INVX2_59/A gnd INVX2_59/Y vdd INVX2
XNAND2X1_352 INVX1_216/Y NOR2X1_198/Y gnd INVX1_219/A vdd NAND2X1
XFILL_26_5_1 gnd vdd FILL
XINVX1_600 INVX1_600/A gnd INVX1_600/Y vdd INVX1
XFILL_6_6_1 gnd vdd FILL
XBUFX2_185 BUFX2_185/A gnd BUFX2_185/Y vdd BUFX2
XNAND3X1_184 OR2X2_80/Y INVX1_120/A NAND3X1_184/C gnd NAND2X1_209/A vdd NAND3X1
XNOR2X1_38 gnd OR2X2_17/B gnd NOR3X1_29/B vdd NOR2X1
XXNOR2X1_223 bloque_bytes[28] INVX1_504/A gnd NAND3X1_507/B vdd XNOR2X1
XNAND3X1_3 NAND3X1_3/A NAND3X1_3/B AOI21X1_7/C gnd NOR2X1_11/B vdd NAND3X1
XINVX2_23 INVX2_23/A gnd INVX2_23/Y vdd INVX2
XNAND2X1_316 AOI21X1_197/A AOI21X1_197/B gnd INVX2_58/A vdd NAND2X1
XNOR2X1_235 BUFX2_193/A XOR2X1_195/Y gnd NOR2X1_235/Y vdd NOR2X1
XOAI21X1_202 AND2X2_71/Y NOR2X1_132/Y INVX1_135/A gnd NAND3X1_211/C vdd OAI21X1
XFILL_36_0_1 gnd vdd FILL
XBUFX2_149 gnd gnd BUFX2_149/Y vdd BUFX2
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XCLKBUF1_26 BUFX4_3/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XNAND3X1_148 OR2X2_64/Y INVX1_98/A NAND3X1_148/C gnd NAND3X1_148/Y vdd NAND3X1
XINVX1_564 bloque_bytes[4] gnd INVX1_564/Y vdd INVX1
XXNOR2X1_187 XNOR2X1_186/Y OAI21X1_466/Y gnd INVX1_376/A vdd XNOR2X1
XOAI21X1_166 AND2X2_58/Y NOR2X1_110/Y INVX1_112/Y gnd NAND3X1_175/A vdd OAI21X1
XNOR2X1_199 BUFX2_181/A XOR2X1_168/Y gnd NOR2X1_199/Y vdd NOR2X1
XNAND2X1_280 INVX1_160/Y OR2X2_111/A gnd NAND2X1_281/A vdd NAND2X1
XNAND3X1_112 OR2X2_48/Y INVX1_76/A NAND3X1_112/C gnd NAND3X1_112/Y vdd NAND3X1
XDFFPOSX1_346 INVX1_415/A CLKBUF1_51/Y OAI21X1_626/Y gnd vdd DFFPOSX1
XNOR3X1_79 NOR3X1_79/A INVX1_399/A NOR3X1_79/C gnd NOR3X1_79/Y vdd NOR3X1
XBUFX2_113 gnd gnd BUFX2_113/Y vdd BUFX2
XINVX1_528 INVX1_528/A gnd INVX1_528/Y vdd INVX1
XXNOR2X1_151 XNOR2X1_151/A XNOR2X1_151/B gnd INVX1_205/A vdd XNOR2X1
XFILL_25_8_0 gnd vdd FILL
XFILL_5_9_0 gnd vdd FILL
XXNOR2X1_73 XOR2X1_78/B XOR2X1_68/Y gnd OR2X2_63/A vdd XNOR2X1
XNOR2X1_163 NOR2X1_163/A NOR3X1_54/Y gnd NOR2X1_163/Y vdd NOR2X1
XOAI21X1_130 NOR3X1_40/Y NOR2X1_93/A NAND3X1_134/B gnd NAND2X1_158/B vdd OAI21X1
XNAND2X1_244 OR2X2_96/B OR2X2_96/A gnd NAND2X1_245/A vdd NAND2X1
XNOR3X1_43 INVX1_110/Y NOR3X1_43/B AND2X2_56/Y gnd NOR3X1_43/Y vdd NOR3X1
XINVX1_492 INVX1_492/A gnd INVX1_492/Y vdd INVX1
XFILL_35_3_0 gnd vdd FILL
XFILL_33_5_1 gnd vdd FILL
XDFFPOSX1_310 INVX1_329/A CLKBUF1_39/Y OR2X2_138/Y gnd vdd DFFPOSX1
XXNOR2X1_37 BUFX2_241/A XOR2X1_28/Y gnd OR2X2_31/A vdd XNOR2X1
XXNOR2X1_115 XNOR2X1_115/A XNOR2X1_115/B gnd BUFX2_169/A vdd XNOR2X1
XXOR2X1_307 XOR2X1_307/A BUFX2_246/A gnd XOR2X1_307/Y vdd XOR2X1
XNOR2X1_127 NOR2X1_127/A NOR2X1_127/B gnd XOR2X1_118/A vdd NOR2X1
XNAND2X1_208 INVX2_40/A AND2X2_60/Y gnd OAI21X1_174/B vdd NAND2X1
XDFFPOSX1_274 INVX1_244/A CLKBUF1_17/Y NOR2X1_431/B gnd vdd DFFPOSX1
XOAI21X1_635 NOR3X1_97/C NOR3X1_97/B INVX1_590/Y gnd NAND3X1_533/B vdd OAI21X1
XOR2X2_95 OR2X2_95/A OR2X2_95/B gnd OR2X2_95/Y vdd OR2X2
XXOR2X1_271 BUFX2_232/A gnd gnd XOR2X1_271/Y vdd XOR2X1
XINVX1_456 INVX1_456/A gnd INVX1_456/Y vdd INVX1
XNAND2X1_172 INVX2_35/Y XNOR2X1_77/A gnd XNOR2X1_78/B vdd NAND2X1
XAOI21X1_70 AOI21X1_68/Y NAND3X1_93/Y OAI21X1_89/B gnd OAI21X1_91/A vdd AOI21X1
XDFFPOSX1_238 INVX1_168/A CLKBUF1_20/Y INVX1_519/A gnd vdd DFFPOSX1
XOAI21X1_599 bloque_bytes[78] INVX2_87/Y OAI21X1_599/C gnd OR2X2_140/A vdd OAI21X1
XOR2X2_59 gnd OR2X2_59/B gnd OR2X2_59/Y vdd OR2X2
XMUX2X1_17 BUFX2_17/A INVX1_10/A MUX2X1_9/S gnd MUX2X1_17/Y vdd MUX2X1
XINVX1_420 INVX1_420/A gnd INVX1_420/Y vdd INVX1
XNAND2X1_713 AND2X2_197/B AND2X2_197/A gnd AOI21X1_400/C vdd NAND2X1
XXOR2X1_235 BUFX2_216/A gnd gnd NOR2X1_287/B vdd XOR2X1
XAOI21X1_372 INVX1_530/Y bloque_bytes[34] AOI21X1_372/C gnd NAND2X1_652/B vdd AOI21X1
XBUFX2_73 gnd gnd BUFX2_73/Y vdd BUFX2
XFILL_32_8_0 gnd vdd FILL
XNAND3X1_545 INVX1_594/A NAND3X1_545/B OR2X2_159/Y gnd OR2X2_162/B vdd NAND3X1
XNAND2X1_136 OAI21X1_110/Y OAI21X1_113/C gnd AOI21X1_93/C vdd NAND2X1
XAOI21X1_34 AOI21X1_32/Y NAND3X1_39/Y AOI21X1_34/C gnd AOI21X1_34/Y vdd AOI21X1
XOR2X2_23 OR2X2_23/A OR2X2_23/B gnd OR2X2_23/Y vdd OR2X2
XDFFPOSX1_202 INVX2_41/A CLKBUF1_50/Y bloque_bytes[0] gnd vdd DFFPOSX1
XINVX1_384 BUFX2_219/A gnd INVX1_384/Y vdd INVX1
XOAI21X1_563 NOR2X1_353/A NOR3X1_85/Y AOI21X1_321/Y gnd AOI21X1_322/B vdd OAI21X1
XBUFX2_37 gnd gnd BUFX2_37/Y vdd BUFX2
XNAND2X1_677 INVX2_88/Y INVX1_552/A gnd NAND2X1_677/Y vdd NAND2X1
XXOR2X1_199 BUFX2_200/A gnd gnd NOR2X1_239/B vdd XOR2X1
XNAND2X1_97 gnd OR2X2_33/B gnd NAND2X1_97/Y vdd NAND2X1
XNAND2X1_100 NAND3X1_80/Y OAI21X1_77/Y gnd XNOR2X1_43/A vdd NAND2X1
XNAND3X1_509 XNOR2X1_213/Y NAND3X1_509/B AND2X2_177/Y gnd AOI21X1_385/C vdd NAND3X1
XAOI21X1_336 AND2X2_166/B AND2X2_171/Y AOI21X1_336/C gnd DFFPOSX1_76/D vdd AOI21X1
XOAI21X1_82 AND2X2_28/Y NOR2X1_60/Y INVX1_57/A gnd AOI21X1_61/A vdd OAI21X1
XDFFPOSX1_166 INVX1_69/A CLKBUF1_44/Y bloque_bytes[44] gnd vdd DFFPOSX1
XXOR2X1_163 BUFX2_180/A gnd gnd NOR2X1_191/B vdd XOR2X1
XOAI21X1_527 gnd XOR2X1_270/Y INVX1_434/A gnd NAND2X1_572/A vdd OAI21X1
XINVX1_348 INVX1_348/A gnd INVX1_348/Y vdd INVX1
XNAND2X1_641 bloque_bytes[73] bloque_bytes[33] gnd AOI21X1_371/A vdd NAND2X1
XOAI21X1_46 OAI21X1_46/A OAI21X1_46/B INVX1_41/A gnd XOR2X1_30/A vdd OAI21X1
XNAND2X1_61 gnd OR2X2_18/B gnd NAND2X1_61/Y vdd NAND2X1
XDFFPOSX1_64 AND2X2_169/B CLKBUF1_38/Y NOR2X1_386/Y gnd vdd DFFPOSX1
XFILL_25_1 gnd vdd FILL
XNAND3X1_473 INVX1_451/Y INVX1_450/A AOI21X1_314/B gnd AND2X2_153/B vdd NAND3X1
XAOI21X1_300 AOI21X1_300/A AOI21X1_300/B INVX1_421/A gnd NOR2X1_328/A vdd AOI21X1
XDFFPOSX1_130 INVX2_14/A CLKBUF1_37/Y bloque_bytes[72] gnd vdd DFFPOSX1
XFILL_16_1_0 gnd vdd FILL
XOAI21X1_491 NOR3X1_80/C INVX2_70/Y NOR3X1_80/A gnd AND2X2_144/A vdd OAI21X1
XINVX1_312 INVX1_312/A gnd INVX1_312/Y vdd INVX1
XFILL_14_3_1 gnd vdd FILL
XXOR2X1_127 XOR2X1_127/A OR2X2_101/A gnd OR2X2_109/B vdd XOR2X1
XNOR2X1_8 NOR2X1_8/A NOR2X1_8/B gnd NOR2X1_8/Y vdd NOR2X1
XNAND2X1_605 INVX1_466/Y NOR2X1_356/B gnd NAND2X1_605/Y vdd NAND2X1
XAOI21X1_264 AOI21X1_264/A AOI21X1_264/B NAND2X1_469/Y gnd AOI21X1_264/Y vdd AOI21X1
XNAND2X1_25 INVX1_19/A NAND2X1_25/B gnd OAI21X1_17/A vdd NAND2X1
XOAI21X1_10 AND2X2_3/Y NOR3X1_26/B INVX1_12/Y gnd NAND3X1_8/A vdd OAI21X1
XDFFPOSX1_28 INVX1_513/A CLKBUF1_20/Y AND2X2_159/Y gnd vdd DFFPOSX1
XNAND3X1_437 INVX1_401/A NAND3X1_437/B INVX2_70/Y gnd NAND3X1_437/Y vdd NAND3X1
XINVX1_276 INVX1_276/A gnd INVX1_276/Y vdd INVX1
XOAI21X1_455 NOR3X1_75/A INVX1_361/A OAI21X1_461/B gnd NOR2X1_290/A vdd OAI21X1
XAOI21X1_4 AOI21X1_4/A AOI21X1_3/Y OAI21X1_5/Y gnd AOI21X1_5/A vdd AOI21X1
XXOR2X1_71 XOR2X1_71/A XOR2X1_71/B gnd XOR2X1_71/Y vdd XOR2X1
XOR2X2_154 OR2X2_149/A OR2X2_141/A gnd OR2X2_154/Y vdd OR2X2
XNAND2X1_569 NAND2X1_569/A AOI22X1_20/C gnd AOI21X1_305/C vdd NAND2X1
XAOI21X1_228 AOI21X1_228/A AOI21X1_228/B INVX1_250/A gnd NOR2X1_220/A vdd AOI21X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XNAND3X1_401 INVX1_346/Y INVX1_347/Y INVX1_348/Y gnd NAND3X1_401/Y vdd NAND3X1
XINVX1_240 INVX1_240/A gnd INVX1_240/Y vdd INVX1
XNAND3X1_66 INVX1_47/Y AOI21X1_52/A OR2X2_28/Y gnd NAND3X1_67/B vdd NAND3X1
XNOR2X1_452 NOR2X1_452/A INVX1_595/Y gnd NOR2X1_452/Y vdd NOR2X1
XXOR2X1_35 XOR2X1_30/Y gnd gnd OR2X2_35/B vdd XOR2X1
XAND2X2_171 INVX2_83/A INVX1_490/Y gnd AND2X2_171/Y vdd AND2X2
XOAI21X1_419 gnd NOR2X1_267/B INVX1_324/Y gnd OAI21X1_419/Y vdd OAI21X1
XNAND2X1_533 INVX1_396/Y NOR2X1_310/Y gnd NAND2X1_534/B vdd NAND2X1
XOR2X2_118 OR2X2_118/A OR2X2_118/B gnd INVX1_170/A vdd OR2X2
XINVX1_86 OR2X2_56/Y gnd INVX1_86/Y vdd INVX1
XFILL_11_8_1 gnd vdd FILL
XFILL_13_6_0 gnd vdd FILL
XAOI21X1_192 AOI21X1_192/A AOI21X1_192/B NAND3X1_279/A gnd NOR2X1_171/A vdd AOI21X1
XNAND3X1_365 INVX1_293/A NAND3X1_365/B NAND3X1_365/C gnd NAND3X1_365/Y vdd NAND3X1
XINVX1_204 INVX1_204/A gnd INVX1_204/Y vdd INVX1
XOAI21X1_383 INVX1_289/A INVX1_290/A INVX1_291/A gnd INVX1_293/A vdd OAI21X1
XAND2X2_135 NOR2X1_287/Y INVX1_359/Y gnd NOR3X1_76/C vdd AND2X2
XNAND3X1_30 INVX1_25/Y NAND3X1_30/B OR2X2_12/Y gnd NAND3X1_31/B vdd NAND3X1
XNOR2X1_416 bloque_bytes[32] OR2X2_142/B gnd NOR2X1_416/Y vdd NOR2X1
XNAND2X1_497 INVX1_359/Y NOR2X1_287/Y gnd NAND2X1_497/Y vdd NAND2X1
XAOI21X1_156 AOI21X1_156/A AOI21X1_156/B NAND3X1_224/C gnd NOR2X1_141/A vdd AOI21X1
XFILL_23_1_0 gnd vdd FILL
XINVX1_50 INVX1_50/A gnd OR2X2_31/B vdd INVX1
XFILL_1_4_1 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XNAND3X1_329 INVX1_231/A OAI21X1_327/Y NAND3X1_324/Y gnd NAND3X1_329/Y vdd NAND3X1
XFILL_21_3_1 gnd vdd FILL
XNOR2X1_380 INVX1_472/Y NOR2X1_383/B gnd NOR2X1_380/Y vdd NOR2X1
XINVX1_168 INVX1_168/A gnd INVX1_168/Y vdd INVX1
XOAI21X1_347 NOR3X1_63/C OAI21X1_347/B INVX1_256/A gnd NOR2X1_221/A vdd OAI21X1
XNAND2X1_461 INVX1_325/A NAND2X1_460/Y gnd NOR3X1_71/B vdd NAND2X1
XNAND3X1_293 INVX2_59/A NAND3X1_293/B NAND3X1_293/C gnd NOR3X1_57/A vdd NAND3X1
XAND2X2_72 AND2X2_72/A AND2X2_72/B gnd AND2X2_72/Y vdd AND2X2
XAOI21X1_120 NAND3X1_175/A AOI21X1_120/B AOI21X1_120/C gnd NOR2X1_111/A vdd AOI21X1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XOAI21X1_311 BUFX2_180/A NOR2X1_198/B INVX1_216/Y gnd NAND3X1_313/B vdd OAI21X1
XINVX1_132 INVX1_132/A gnd INVX1_132/Y vdd INVX1
XNAND2X1_425 INVX1_286/Y NOR2X1_243/Y gnd AOI21X1_245/B vdd NAND2X1
XNOR2X1_344 INVX1_447/Y NOR2X1_344/B gnd INVX1_449/A vdd NOR2X1
XBUFX2_258 XOR2X1_71/A gnd BUFX2_258/Y vdd BUFX2
XAND2X2_36 AND2X2_36/A AND2X2_36/B gnd AND2X2_36/Y vdd AND2X2
XNAND3X1_257 INVX1_165/A NAND3X1_257/B OR2X2_113/Y gnd NAND3X1_260/B vdd NAND3X1
XOAI21X1_275 AND2X2_97/Y NOR2X1_174/Y INVX1_180/Y gnd NAND3X1_289/A vdd OAI21X1
XFILL_20_6_0 gnd vdd FILL
XBUFX4_21 BUFX4_18/A gnd BUFX4_21/Y vdd BUFX4
XFILL_0_7_0 gnd vdd FILL
XFILL_18_8_1 gnd vdd FILL
XNAND2X1_389 INVX1_254/A NOR2X1_222/Y gnd NAND3X1_339/C vdd NAND2X1
XNOR2X1_308 INVX1_390/Y NOR2X1_308/B gnd INVX1_392/A vdd NOR2X1
XNAND3X1_221 INVX1_143/A NAND2X1_249/Y OR2X2_97/Y gnd NAND2X1_250/B vdd NAND3X1
XNOR2X1_75 NOR2X1_75/A INVX1_71/Y gnd NOR2X1_75/Y vdd NOR2X1
XBUFX2_222 BUFX2_222/A gnd BUFX2_222/Y vdd BUFX2
XINVX2_60 INVX2_60/A gnd INVX2_60/Y vdd INVX2
XOAI21X1_239 XNOR2X1_125/A OAI21X1_239/B AND2X2_84/B gnd XNOR2X1_126/A vdd OAI21X1
XNOR2X1_272 INVX1_333/Y NOR2X1_272/B gnd INVX1_335/A vdd NOR2X1
XFILL_30_1_0 gnd vdd FILL
XFILL_28_3_1 gnd vdd FILL
XFILL_8_4_1 gnd vdd FILL
XNAND2X1_353 AOI21X1_217/A AOI21X1_217/B gnd XOR2X1_179/B vdd NAND2X1
XBUFX2_186 BUFX2_186/A gnd BUFX2_186/Y vdd BUFX2
XNAND3X1_185 INVX1_121/A NAND3X1_185/B OR2X2_81/Y gnd NAND3X1_185/Y vdd NAND3X1
XNAND3X1_4 AND2X2_1/Y NAND3X1_4/B NAND3X1_4/C gnd NOR2X1_16/B vdd NAND3X1
XNOR2X1_39 gnd OR2X2_18/B gnd NOR3X1_30/B vdd NOR2X1
XXNOR2X1_224 bloque_bytes[30] INVX1_548/A gnd XNOR2X1_224/Y vdd XNOR2X1
XOAI21X1_203 AND2X2_71/Y NOR2X1_132/Y INVX1_135/Y gnd NAND3X1_213/A vdd OAI21X1
XINVX2_24 INVX2_24/A gnd INVX2_24/Y vdd INVX2
XNAND2X1_317 NAND3X1_289/A OR2X2_128/B gnd OR2X2_126/A vdd NAND2X1
XNOR2X1_236 INVX1_276/Y NOR2X1_236/B gnd INVX1_278/A vdd NOR2X1
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XNAND3X1_149 INVX1_99/A NAND2X1_173/Y OR2X2_65/Y gnd NAND3X1_152/B vdd NAND3X1
XCLKBUF1_27 BUFX4_1/Y gnd CLKBUF1_27/Y vdd CLKBUF1
XBUFX2_150 gnd gnd BUFX2_150/Y vdd BUFX2
XINVX1_565 INVX1_565/A gnd INVX1_565/Y vdd INVX1
XXNOR2X1_188 NOR2X1_302/A NAND2X1_521/Y gnd BUFX2_230/A vdd XNOR2X1
XNOR2X1_200 INVX1_219/Y NOR2X1_200/B gnd INVX1_221/A vdd NOR2X1
XOAI21X1_167 AND2X2_58/Y NOR2X1_110/Y INVX1_112/A gnd AOI21X1_121/A vdd OAI21X1
XNAND2X1_281 NAND2X1_281/A OR2X2_111/Y gnd OR2X2_112/A vdd NAND2X1
XNOR3X1_80 NOR3X1_80/A INVX2_70/Y NOR3X1_80/C gnd NOR3X1_80/Y vdd NOR3X1
XNAND3X1_113 INVX1_77/A NAND3X1_113/B OR2X2_49/Y gnd OAI21X1_113/C vdd NAND3X1
XINVX1_529 INVX1_529/A gnd INVX1_529/Y vdd INVX1
XFILL_25_8_1 gnd vdd FILL
XDFFPOSX1_347 INVX1_416/A CLKBUF1_8/Y OAI21X1_627/Y gnd vdd DFFPOSX1
XFILL_27_6_0 gnd vdd FILL
XBUFX2_114 gnd gnd BUFX2_114/Y vdd BUFX2
XFILL_5_9_1 gnd vdd FILL
XFILL_7_7_0 gnd vdd FILL
XXNOR2X1_74 XOR2X1_81/Y XOR2X1_69/Y gnd XNOR2X1_75/A vdd XNOR2X1
XXNOR2X1_152 NOR2X1_194/A XNOR2X1_152/B gnd BUFX2_190/A vdd XNOR2X1
XNOR2X1_164 OR2X2_117/A OR2X2_117/B gnd NOR2X1_164/Y vdd NOR2X1
XNAND2X1_245 NAND2X1_245/A OR2X2_96/Y gnd INVX1_139/A vdd NAND2X1
XOAI21X1_131 OAI21X1_131/A XNOR2X1_70/B INVX1_96/A gnd XOR2X1_80/A vdd OAI21X1
XNOR3X1_44 INVX1_111/Y NOR3X1_44/B AND2X2_57/Y gnd NOR3X1_44/Y vdd NOR3X1
XDFFPOSX1_311 INVX1_330/A CLKBUF1_34/Y INVX1_555/Y gnd vdd DFFPOSX1
XINVX1_493 bloque_bytes[24] gnd INVX1_493/Y vdd INVX1
XFILL_35_3_1 gnd vdd FILL
XXNOR2X1_38 XOR2X1_41/Y XOR2X1_29/Y gnd XNOR2X1_39/A vdd XNOR2X1
XXNOR2X1_116 XNOR2X1_116/A AND2X2_78/Y gnd XOR2X1_136/A vdd XNOR2X1
XXOR2X1_308 XOR2X1_308/A XOR2X1_295/Y gnd XOR2X1_308/Y vdd XOR2X1
XNOR2X1_128 gnd OR2X2_89/B gnd NOR3X1_47/B vdd NOR2X1
XNAND2X1_209 NAND2X1_209/A NAND2X1_209/B gnd XOR2X1_109/A vdd NAND2X1
XDFFPOSX1_275 INVX1_245/A CLKBUF1_27/Y NOR2X1_432/B gnd vdd DFFPOSX1
XOAI21X1_636 NOR3X1_98/Y NOR2X1_450/A NOR3X1_97/Y gnd NAND2X1_708/B vdd OAI21X1
XOR2X2_96 OR2X2_96/A OR2X2_96/B gnd OR2X2_96/Y vdd OR2X2
XINVX1_457 INVX1_457/A gnd INVX1_457/Y vdd INVX1
XXOR2X1_272 BUFX2_233/A gnd gnd NOR2X1_336/B vdd XOR2X1
XNAND2X1_173 gnd OR2X2_65/B gnd NAND2X1_173/Y vdd NAND2X1
XOAI21X1_600 bloque_bytes[79] INVX1_505/Y AND2X2_177/A gnd OR2X2_141/A vdd OAI21X1
XAOI21X1_71 NAND3X1_97/B OR2X2_42/Y INVX1_67/A gnd NOR2X1_73/A vdd AOI21X1
XDFFPOSX1_239 INVX1_169/A CLKBUF1_9/Y INVX1_522/A gnd vdd DFFPOSX1
XOR2X2_60 OR2X2_60/A OR2X2_60/B gnd OR2X2_60/Y vdd OR2X2
XMUX2X1_18 BUFX2_18/A MUX2X1_18/B MUX2X1_9/S gnd MUX2X1_18/Y vdd MUX2X1
XINVX1_421 INVX1_421/A gnd INVX1_421/Y vdd INVX1
XNAND2X1_714 gnd gnd gnd NAND3X1_545/B vdd NAND2X1
XBUFX2_74 gnd gnd BUFX2_74/Y vdd BUFX2
XXOR2X1_236 BUFX2_217/A gnd gnd XOR2X1_236/Y vdd XOR2X1
XFILL_34_6_0 gnd vdd FILL
XNAND2X1_137 gnd OR2X2_50/B gnd AOI21X1_83/A vdd NAND2X1
XAOI21X1_373 NAND2X1_644/Y OR2X2_133/Y INVX1_503/A gnd NAND2X1_653/B vdd AOI21X1
XFILL_32_8_1 gnd vdd FILL
XNAND3X1_546 NAND3X1_546/A OR2X2_162/B OR2X2_160/B gnd AOI21X1_400/B vdd NAND3X1
XAOI21X1_35 NAND2X1_61/Y OR2X2_18/Y INVX1_34/A gnd NOR2X1_43/A vdd AOI21X1
XDFFPOSX1_203 INVX1_121/A CLKBUF1_49/Y bloque_bytes[1] gnd vdd DFFPOSX1
XOR2X2_24 OR2X2_24/A OR2X2_24/B gnd OR2X2_24/Y vdd OR2X2
XXOR2X1_200 BUFX2_201/A gnd gnd XOR2X1_200/Y vdd XOR2X1
XINVX1_385 INVX1_385/A gnd INVX1_385/Y vdd INVX1
XOAI21X1_564 OAI21X1_564/A INVX1_468/A INVX1_471/A gnd NAND2X1_608/A vdd OAI21X1
XNAND2X1_678 INVX2_89/Y INVX1_553/A gnd NAND2X1_678/Y vdd NAND2X1
XBUFX2_38 gnd gnd BUFX2_38/Y vdd BUFX2
XOAI21X1_83 AND2X2_29/Y NOR2X1_62/Y INVX1_58/A gnd NAND3X1_85/C vdd OAI21X1
XNAND2X1_101 INVX1_63/A OAI21X1_79/Y gnd OAI21X1_85/A vdd NAND2X1
XNAND2X1_98 OAI21X1_76/Y NAND3X1_77/Y gnd NAND2X1_98/Y vdd NAND2X1
XNAND3X1_510 NAND2X1_657/A NAND3X1_510/B NOR2X1_410/Y gnd AOI21X1_386/C vdd NAND3X1
XAOI21X1_337 INVX1_479/Y NAND2X1_624/Y NAND2X1_627/Y gnd DFFPOSX1_77/D vdd AOI21X1
XDFFPOSX1_167 INVX1_70/A CLKBUF1_44/Y bloque_bytes[45] gnd vdd DFFPOSX1
XINVX1_349 INVX1_349/A gnd INVX1_349/Y vdd INVX1
XFILL_3_1 gnd vdd FILL
XXOR2X1_164 BUFX2_181/A gnd gnd NOR2X1_192/B vdd XOR2X1
XNAND2X1_642 AOI21X1_371/A OR2X2_132/Y gnd NAND2X1_642/Y vdd NAND2X1
XOAI21X1_528 gnd XOR2X1_271/Y INVX1_435/A gnd INVX2_72/A vdd OAI21X1
XAOI21X1_301 INVX1_421/A NAND3X1_452/B INVX1_420/Y gnd NOR3X1_81/C vdd AOI21X1
XOAI21X1_47 AND2X2_16/Y NOR2X1_40/Y INVX1_35/Y gnd AOI21X1_36/A vdd OAI21X1
XNAND2X1_62 NAND2X1_62/A NAND2X1_62/B gnd XNOR2X1_25/A vdd NAND2X1
XDFFPOSX1_65 INVX1_475/A CLKBUF1_38/Y DFFPOSX1_65/D gnd vdd DFFPOSX1
XFILL_25_2 gnd vdd FILL
XNAND3X1_474 INVX1_449/Y INVX1_452/Y AND2X2_153/A gnd NAND2X1_589/B vdd NAND3X1
XDFFPOSX1_131 INVX1_22/A CLKBUF1_1/Y bloque_bytes[73] gnd vdd DFFPOSX1
XFILL_16_1_1 gnd vdd FILL
XINVX1_313 INVX1_313/A gnd INVX1_313/Y vdd INVX1
XOAI21X1_492 gnd XOR2X1_254/Y INVX1_398/A gnd INVX1_401/A vdd OAI21X1
XXOR2X1_128 XOR2X1_128/A BUFX2_161/A gnd XOR2X1_128/Y vdd XOR2X1
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XNAND2X1_606 NAND2X1_605/Y INVX1_468/Y gnd INVX1_469/A vdd NAND2X1
XNAND2X1_26 gnd OR2X2_3/B gnd AOI21X1_14/A vdd NAND2X1
XAOI21X1_265 NAND3X1_391/Y AOI21X1_265/B NAND2X1_474/Y gnd AOI21X1_265/Y vdd AOI21X1
XNAND3X1_438 INVX1_401/A NAND3X1_438/B NAND3X1_438/C gnd NAND3X1_445/B vdd NAND3X1
XOAI21X1_11 OAI21X1_9/A OAI21X1_9/B NAND3X1_6/A gnd NAND2X1_25/B vdd OAI21X1
XDFFPOSX1_29 INVX1_516/A CLKBUF1_20/Y NOR2X1_359/Y gnd vdd DFFPOSX1
XXOR2X1_72 OR2X2_68/A gnd gnd XOR2X1_72/Y vdd XOR2X1
XINVX1_277 INVX1_277/A gnd INVX1_277/Y vdd INVX1
XOAI21X1_456 NOR3X1_76/A NOR3X1_76/C INVX2_68/A gnd NOR2X1_289/A vdd OAI21X1
XAOI21X1_5 AOI21X1_5/A AOI21X1_5/B AOI21X1_5/C gnd AOI21X1_5/Y vdd AOI21X1
XOR2X2_155 gnd gnd gnd OR2X2_155/Y vdd OR2X2
XNAND2X1_570 OAI21X1_526/Y NAND3X1_461/Y gnd XOR2X1_286/A vdd NAND2X1
XAOI21X1_229 INVX1_250/A NAND2X1_387/Y INVX1_249/Y gnd NOR3X1_63/C vdd AOI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XNAND3X1_402 INVX1_348/A INVX1_346/Y INVX1_347/Y gnd NAND3X1_402/Y vdd NAND3X1
XINVX1_241 INVX1_241/A gnd INVX1_241/Y vdd INVX1
XOAI21X1_420 gnd NOR2X1_267/B INVX1_324/A gnd INVX1_326/A vdd OAI21X1
XNOR2X1_453 INVX1_597/Y NOR2X1_453/B gnd NOR2X1_454/B vdd NOR2X1
XNAND3X1_67 NAND3X1_67/A NAND3X1_67/B NAND3X1_67/C gnd AND2X2_24/B vdd NAND3X1
XXOR2X1_36 XOR2X1_36/A OR2X2_28/A gnd OR2X2_36/B vdd XOR2X1
XAND2X2_172 INVX2_83/A AND2X2_172/B gnd AND2X2_172/Y vdd AND2X2
XOR2X2_119 OR2X2_119/A OR2X2_119/B gnd OR2X2_119/Y vdd OR2X2
XNAND2X1_534 OAI21X1_489/Y NAND2X1_534/B gnd BUFX2_231/A vdd NAND2X1
XFILL_15_4_0 gnd vdd FILL
XAOI21X1_193 AOI21X1_193/A AOI21X1_193/B NOR3X1_56/Y gnd INVX2_57/A vdd AOI21X1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XFILL_13_6_1 gnd vdd FILL
XNAND3X1_366 AOI22X1_13/B INVX1_295/A INVX1_293/Y gnd AOI21X1_249/B vdd NAND3X1
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XNOR2X1_417 bloque_bytes[33] OR2X2_143/B gnd NOR2X1_417/Y vdd NOR2X1
XOAI21X1_384 INVX1_289/A INVX1_290/A INVX1_291/Y gnd OAI21X1_384/Y vdd OAI21X1
XAND2X2_136 AND2X2_136/A NOR3X1_75/A gnd BUFX2_224/A vdd AND2X2
XNAND3X1_31 AOI21X1_24/A NAND3X1_31/B OAI21X1_32/Y gnd AND2X2_12/B vdd NAND3X1
XNAND2X1_498 INVX1_360/Y NOR2X1_288/Y gnd NAND2X1_499/B vdd NAND2X1
XFILL_5_0_0 gnd vdd FILL
XNAND3X1_330 INVX1_242/Y INVX1_241/A AOI21X1_226/B gnd AND2X2_109/B vdd NAND3X1
XAOI21X1_157 AOI21X1_157/A AOI21X1_157/B NOR3X1_50/Y gnd INVX2_48/A vdd AOI21X1
XFILL_23_1_1 gnd vdd FILL
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XFILL_3_2_1 gnd vdd FILL
XNOR2X1_381 MUX2X1_3/S INVX1_487/Y gnd NOR2X1_381/Y vdd NOR2X1
XAND2X2_100 AND2X2_100/A NOR3X1_57/A gnd BUFX2_184/A vdd AND2X2
XINVX1_169 INVX1_169/A gnd INVX1_169/Y vdd INVX1
XOAI21X1_348 NOR2X1_221/Y NOR2X1_220/B AOI22X1_11/C gnd XOR2X1_197/A vdd OAI21X1
XNAND2X1_462 INVX1_324/A NOR2X1_267/Y gnd NAND2X1_462/Y vdd NAND2X1
XNAND3X1_294 INVX1_192/A NAND2X1_328/B INVX2_59/Y gnd OAI21X1_284/C vdd NAND3X1
XAND2X2_73 OR2X2_93/A OR2X2_93/B gnd AND2X2_73/Y vdd AND2X2
XAOI21X1_121 AOI21X1_121/A AOI21X1_121/B NOR3X1_44/Y gnd INVX2_39/A vdd AOI21X1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XFILL_12_9_0 gnd vdd FILL
XOAI21X1_312 BUFX2_180/A NOR2X1_198/B INVX1_216/A gnd AOI22X1_9/B vdd OAI21X1
XINVX1_133 INVX1_133/A gnd INVX1_133/Y vdd INVX1
XNAND2X1_426 NAND3X1_360/Y INVX1_294/A gnd XNOR2X1_168/B vdd NAND2X1
XNOR2X1_345 BUFX2_234/A NOR2X1_345/B gnd NOR2X1_345/Y vdd NOR2X1
XAND2X2_37 OR2X2_45/A OR2X2_45/B gnd AND2X2_37/Y vdd AND2X2
XNAND3X1_258 NAND3X1_260/B OAI21X1_246/Y NAND3X1_258/C gnd NAND3X1_258/Y vdd NAND3X1
XBUFX2_259 OR2X2_60/A gnd BUFX2_259/Y vdd BUFX2
XFILL_2_5_0 gnd vdd FILL
XOAI21X1_276 XNOR2X1_143/A NAND2X1_322/Y NOR2X1_175/Y gnd NOR2X1_176/B vdd OAI21X1
XFILL_20_6_1 gnd vdd FILL
XFILL_22_4_0 gnd vdd FILL
XBUFX4_22 BUFX4_18/A gnd NOR3X1_2/C vdd BUFX4
XNOR2X1_309 BUFX2_222/A NOR2X1_309/B gnd NOR2X1_309/Y vdd NOR2X1
XFILL_0_7_1 gnd vdd FILL
XNAND2X1_390 INVX1_254/Y NOR2X1_222/Y gnd INVX1_257/A vdd NAND2X1
XNAND3X1_222 NAND2X1_250/B NAND2X1_250/A XNOR2X1_114/B gnd XNOR2X1_115/B vdd NAND3X1
XBUFX2_223 BUFX2_223/A gnd BUFX2_223/Y vdd BUFX2
XNOR2X1_76 INVX1_73/Y NOR2X1_76/B gnd NOR2X1_76/Y vdd NOR2X1
XOAI21X1_240 AND2X2_85/Y NOR2X1_154/Y INVX1_158/A gnd NAND3X1_251/B vdd OAI21X1
XFILL_30_1_1 gnd vdd FILL
XINVX2_61 INVX2_61/A gnd INVX2_61/Y vdd INVX2
XNAND2X1_354 INVX1_208/A NOR2X1_192/Y gnd AOI21X1_214/B vdd NAND2X1
XNOR2X1_273 BUFX2_210/A XOR2X1_223/Y gnd NOR2X1_273/Y vdd NOR2X1
XNAND3X1_5 INVX1_11/A NAND3X1_5/B OR2X2_1/Y gnd NAND3X1_6/A vdd NAND3X1
XNAND3X1_186 NAND3X1_185/Y OAI21X1_178/Y XNOR2X1_96/B gnd XNOR2X1_97/B vdd NAND3X1
XBUFX2_187 INVX1_251/A gnd BUFX2_187/Y vdd BUFX2
XNOR2X1_40 gnd OR2X2_19/B gnd NOR2X1_40/Y vdd NOR2X1
XXNOR2X1_225 bloque_bytes[31] OR2X2_149/B gnd NAND3X1_509/B vdd XNOR2X1
XOAI21X1_204 OAI21X1_199/A XNOR2X1_106/B OAI21X1_204/C gnd OAI21X1_204/Y vdd OAI21X1
XINVX2_25 INVX2_25/A gnd INVX2_25/Y vdd INVX2
XNOR2X1_237 BUFX2_194/A XOR2X1_196/Y gnd NOR2X1_237/Y vdd NOR2X1
XNAND2X1_318 OR2X2_127/B OR2X2_127/A gnd NAND2X1_319/A vdd NAND2X1
XNAND3X1_150 NAND3X1_152/B OAI21X1_144/Y XNOR2X1_78/B gnd XNOR2X1_79/B vdd NAND3X1
XFILL_19_9_0 gnd vdd FILL
XINVX1_566 INVX1_566/A gnd INVX1_566/Y vdd INVX1
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XBUFX2_151 XOR2X1_2/A gnd BUFX2_151/Y vdd BUFX2
XXNOR2X1_189 NOR2X1_305/Y NOR2X1_304/Y gnd XOR2X1_265/A vdd XNOR2X1
XCLKBUF1_28 BUFX4_2/Y gnd CLKBUF1_28/Y vdd CLKBUF1
XNOR2X1_201 BUFX2_182/A NOR2X1_201/B gnd NOR2X1_201/Y vdd NOR2X1
XFILL_16_1 gnd vdd FILL
XOAI21X1_168 AND2X2_59/Y NOR2X1_112/Y INVX1_113/A gnd NAND3X1_175/C vdd OAI21X1
XNAND2X1_282 OR2X2_112/B OR2X2_112/A gnd NAND2X1_283/A vdd NAND2X1
XFILL_29_4_0 gnd vdd FILL
XNOR3X1_81 NOR3X1_81/A INVX1_418/A NOR3X1_81/C gnd NOR3X1_81/Y vdd NOR3X1
XNAND3X1_114 OAI21X1_113/C OAI21X1_110/Y XNOR2X1_60/B gnd XNOR2X1_61/B vdd NAND3X1
XFILL_9_5_0 gnd vdd FILL
XINVX1_530 bloque_bytes[74] gnd INVX1_530/Y vdd INVX1
XDFFPOSX1_348 INVX1_417/A CLKBUF1_2/Y OAI21X1_628/Y gnd vdd DFFPOSX1
XFILL_27_6_1 gnd vdd FILL
XBUFX2_115 gnd gnd BUFX2_115/Y vdd BUFX2
XFILL_7_7_1 gnd vdd FILL
XXNOR2X1_75 XNOR2X1_75/A OR2X2_63/Y gnd INVX1_98/A vdd XNOR2X1
XXNOR2X1_153 NOR2X1_197/Y NOR2X1_196/Y gnd XOR2X1_184/A vdd XNOR2X1
XOAI21X1_132 AND2X2_46/Y NOR2X1_90/Y INVX1_90/Y gnd AOI21X1_96/A vdd OAI21X1
XNOR2X1_165 NOR2X1_165/A INVX1_170/Y gnd NOR2X1_165/Y vdd NOR2X1
XNAND2X1_246 INVX2_46/A AND2X2_72/Y gnd AOI21X1_154/C vdd NAND2X1
XNOR3X1_45 INVX1_121/Y NOR3X1_45/B AND2X2_62/Y gnd NOR3X1_45/Y vdd NOR3X1
XDFFPOSX1_312 INVX1_334/A CLKBUF1_23/Y INVX1_556/Y gnd vdd DFFPOSX1
XXOR2X1_309 gnd vdd gnd XNOR2X1_4/B vdd XOR2X1
XXNOR2X1_117 XNOR2X1_117/A INVX2_49/Y gnd XOR2X1_137/A vdd XNOR2X1
XINVX1_494 bloque_bytes[25] gnd INVX1_494/Y vdd INVX1
XXNOR2X1_39 XNOR2X1_39/A OR2X2_31/Y gnd INVX1_54/A vdd XNOR2X1
XNOR2X1_129 gnd OR2X2_90/B gnd NOR3X1_48/B vdd NOR2X1
XNAND2X1_210 INVX2_41/Y XNOR2X1_94/Y gnd XNOR2X1_96/B vdd NAND2X1
XOAI21X1_637 NOR3X1_98/C NOR3X1_98/B NOR3X1_98/A gnd NAND3X1_535/A vdd OAI21X1
XOR2X2_97 gnd OR2X2_97/B gnd OR2X2_97/Y vdd OR2X2
XDFFPOSX1_276 INVX1_246/A CLKBUF1_32/Y NOR2X1_433/B gnd vdd DFFPOSX1
XINVX1_458 INVX1_458/A gnd INVX1_458/Y vdd INVX1
XFILL_26_9_0 gnd vdd FILL
XXOR2X1_273 BUFX2_234/A gnd gnd NOR2X1_339/B vdd XOR2X1
XNAND2X1_174 OAI21X1_144/Y NAND3X1_152/B gnd XNOR2X1_78/A vdd NAND2X1
XDFFPOSX1_240 INVX1_171/A CLKBUF1_26/Y INVX1_525/A gnd vdd DFFPOSX1
XAOI21X1_72 OAI21X1_98/Y AOI21X1_72/B AOI21X1_72/C gnd NOR2X1_71/A vdd AOI21X1
XOAI21X1_601 INVX1_506/Y bloque_bytes[16] INVX1_507/Y gnd AOI21X1_362/C vdd OAI21X1
XOR2X2_61 OR2X2_61/A OR2X2_61/B gnd OR2X2_61/Y vdd OR2X2
XINVX1_422 INVX1_422/A gnd INVX1_422/Y vdd INVX1
XMUX2X1_19 BUFX2_19/A INVX1_9/A BUFX4_9/Y gnd MUX2X1_19/Y vdd MUX2X1
XNAND2X1_715 AOI21X1_400/A AOI21X1_400/B gnd INVX2_94/A vdd NAND2X1
XBUFX2_75 gnd gnd BUFX2_75/Y vdd BUFX2
XXOR2X1_237 BUFX2_218/A gnd gnd NOR2X1_291/B vdd XOR2X1
XFILL_36_4_0 gnd vdd FILL
XFILL_34_6_1 gnd vdd FILL
XNAND3X1_547 INVX2_93/Y NAND3X1_547/B NAND2X1_712/B gnd AOI21X1_402/B vdd NAND3X1
XNAND2X1_138 NAND2X1_138/A OAI21X1_111/Y gnd XNOR2X1_61/A vdd NAND2X1
XAOI21X1_374 NAND2X1_647/Y OR2X2_134/Y INVX1_504/A gnd AOI21X1_374/Y vdd AOI21X1
XAOI21X1_36 AOI21X1_36/A AOI21X1_36/B AOI21X1_36/C gnd NOR2X1_41/A vdd AOI21X1
XDFFPOSX1_204 INVX1_122/A CLKBUF1_49/Y bloque_bytes[2] gnd vdd DFFPOSX1
XOR2X2_25 gnd OR2X2_25/B gnd OR2X2_25/Y vdd OR2X2
XOAI21X1_565 NOR2X1_381/Y INVX1_472/A BUFX4_30/Y gnd NOR2X1_382/B vdd OAI21X1
XXOR2X1_201 BUFX2_202/A gnd gnd XOR2X1_201/Y vdd XOR2X1
XINVX1_386 INVX1_386/A gnd INVX1_386/Y vdd INVX1
XBUFX2_39 gnd gnd BUFX2_39/Y vdd BUFX2
XNAND2X1_679 OR2X2_144/B OR2X2_144/A gnd AOI21X1_389/A vdd NAND2X1
XOAI21X1_84 AND2X2_29/Y NOR2X1_62/Y INVX1_58/Y gnd OAI21X1_84/Y vdd OAI21X1
XNAND2X1_102 gnd OR2X2_35/B gnd NAND3X1_83/B vdd NAND2X1
XNAND2X1_99 gnd OR2X2_34/B gnd NAND2X1_99/Y vdd NAND2X1
XAOI21X1_338 INVX1_480/A AND2X2_172/Y OAI21X1_580/Y gnd AOI21X1_338/Y vdd AOI21X1
XNAND3X1_511 XNOR2X1_215/Y XNOR2X1_227/Y NOR2X1_411/Y gnd AOI21X1_387/C vdd NAND3X1
XDFFPOSX1_168 INVX1_72/A CLKBUF1_7/Y bloque_bytes[46] gnd vdd DFFPOSX1
XFILL_10_2_0 gnd vdd FILL
XINVX1_350 INVX1_350/A gnd INVX1_350/Y vdd INVX1
XOAI21X1_529 NOR3X1_84/C INVX2_72/Y NOR3X1_84/A gnd AND2X2_152/A vdd OAI21X1
XXOR2X1_165 BUFX2_182/A gnd gnd XOR2X1_165/Y vdd XOR2X1
XNAND2X1_643 INVX1_502/Y NAND2X1_642/Y gnd OR2X2_151/B vdd NAND2X1
XAOI21X1_302 AOI21X1_302/A NAND2X1_563/Y INVX2_71/A gnd AOI21X1_302/Y vdd AOI21X1
XOAI21X1_48 AND2X2_16/Y NOR2X1_40/Y INVX1_35/A gnd AOI21X1_37/A vdd OAI21X1
XNAND2X1_63 INVX1_41/A NAND2X1_63/B gnd OAI21X1_46/A vdd NAND2X1
XDFFPOSX1_132 INVX1_23/A CLKBUF1_37/Y bloque_bytes[74] gnd vdd DFFPOSX1
XDFFPOSX1_66 AND2X2_161/B CLKBUF1_26/Y DFFPOSX1_66/D gnd vdd DFFPOSX1
XFILL_33_9_0 gnd vdd FILL
XNAND3X1_475 INVX2_73/A NAND3X1_475/B NAND3X1_475/C gnd NOR3X1_85/A vdd NAND3X1
XXOR2X1_129 XOR2X1_129/A BUFX2_162/A gnd XOR2X1_129/Y vdd XOR2X1
XOAI21X1_493 NOR3X1_79/A INVX1_399/A NAND3X1_437/Y gnd NOR2X1_314/A vdd OAI21X1
XINVX1_314 INVX1_314/A gnd INVX1_314/Y vdd INVX1
XNAND2X1_607 NAND2X1_607/A AOI22X1_22/C gnd AOI21X1_321/C vdd NAND2X1
XOAI21X1_12 OAI21X1_17/A XNOR2X1_7/B INVX1_19/A gnd XOR2X1_10/A vdd OAI21X1
XNAND2X1_27 gnd OR2X2_4/B gnd NAND3X1_14/B vdd NAND2X1
XAOI21X1_266 INVX1_337/Y AOI21X1_266/B INVX1_336/A gnd OAI21X1_431/A vdd AOI21X1
XNAND3X1_439 INVX1_402/A NAND3X1_439/B INVX1_401/Y gnd INVX1_408/A vdd NAND3X1
XDFFPOSX1_30 INVX1_519/A CLKBUF1_20/Y NOR2X1_360/Y gnd vdd DFFPOSX1
XINVX1_278 INVX1_278/A gnd INVX1_278/Y vdd INVX1
XAOI21X1_6 AND2X2_1/A AND2X2_1/B AOI21X1_8/C gnd AOI21X1_6/Y vdd AOI21X1
XXOR2X1_73 OR2X2_69/A gnd gnd OR2X2_65/B vdd XOR2X1
XNAND2X1_571 INVX1_434/Y NOR2X1_334/Y gnd NAND3X1_462/B vdd NAND2X1
XOAI21X1_457 gnd NOR2X1_291/B INVX1_362/Y gnd OAI21X1_457/Y vdd OAI21X1
XOR2X2_156 gnd gnd gnd OR2X2_156/Y vdd OR2X2
XAOI21X1_230 AOI21X1_230/A AOI21X1_230/B INVX2_62/A gnd AOI21X1_231/B vdd AOI21X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XNAND3X1_403 INVX1_350/A NAND3X1_401/Y INVX1_345/Y gnd AOI22X1_16/C vdd NAND3X1
XAND2X2_173 INVX2_83/A INVX2_84/Y gnd AND2X2_173/Y vdd AND2X2
XINVX1_242 INVX1_242/A gnd INVX1_242/Y vdd INVX1
XOAI21X1_421 BUFX2_207/A INVX1_328/A INVX1_329/A gnd INVX1_331/A vdd OAI21X1
XNAND3X1_68 INVX1_47/A AOI21X1_52/A OR2X2_28/Y gnd NAND3X1_68/Y vdd NAND3X1
XNOR2X1_454 NOR2X1_454/A NOR2X1_454/B gnd XOR2X1_8/A vdd NOR2X1
XXOR2X1_37 XOR2X1_37/A OR2X2_29/A gnd OR2X2_37/B vdd XOR2X1
XOR2X2_120 OR2X2_120/A OR2X2_120/B gnd INVX1_174/A vdd OR2X2
XFILL_17_2_0 gnd vdd FILL
XNAND2X1_535 INVX1_397/Y NOR2X1_311/Y gnd NAND3X1_436/C vdd NAND2X1
XFILL_15_4_1 gnd vdd FILL
XAOI21X1_194 NAND3X1_281/B OR2X2_123/Y INVX1_178/A gnd AOI21X1_194/Y vdd AOI21X1
XNAND3X1_367 INVX1_285/Y NAND3X1_360/Y NOR3X1_68/Y gnd AOI21X1_248/B vdd NAND3X1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_206 INVX1_206/A gnd INVX1_206/Y vdd INVX1
XNOR2X1_418 INVX2_85/Y INVX1_544/Y gnd NOR2X1_418/Y vdd NOR2X1
XOAI21X1_385 NOR3X1_67/C OAI21X1_385/B INVX1_294/A gnd NOR2X1_245/A vdd OAI21X1
XAND2X2_137 AND2X2_137/A AND2X2_137/B gnd XOR2X1_258/A vdd AND2X2
XNAND3X1_32 INVX1_25/A NAND3X1_30/B OR2X2_12/Y gnd NAND3X1_33/B vdd NAND3X1
XNAND2X1_499 INVX1_363/A NAND2X1_499/B gnd INVX1_361/A vdd NAND2X1
XFILL_5_0_1 gnd vdd FILL
XNAND3X1_331 INVX1_240/Y INVX1_243/Y AND2X2_109/A gnd NAND3X1_331/Y vdd NAND3X1
XAOI21X1_158 NAND3X1_227/B OR2X2_99/Y INVX1_145/A gnd NAND3X1_231/C vdd AOI21X1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_170 INVX1_170/A gnd INVX1_170/Y vdd INVX1
XOAI21X1_349 BUFX2_188/A NOR2X1_222/B INVX1_254/Y gnd NAND3X1_339/B vdd OAI21X1
XNOR2X1_382 NOR2X1_380/Y NOR2X1_382/B gnd NOR2X1_382/Y vdd NOR2X1
XAND2X2_101 AND2X2_101/A AND2X2_101/B gnd AND2X2_101/Y vdd AND2X2
XNAND2X1_463 INVX1_324/Y NOR2X1_267/Y gnd AOI21X1_261/B vdd NAND2X1
XAOI21X1_122 NAND3X1_173/B OR2X2_75/Y INVX1_112/A gnd NAND3X1_177/C vdd AOI21X1
XINVX1_16 OR2X2_6/Y gnd INVX1_16/Y vdd INVX1
XNAND3X1_295 INVX1_192/A NAND3X1_295/B NAND2X1_329/Y gnd NAND2X1_331/A vdd NAND3X1
XAND2X2_74 gnd OR2X2_97/B gnd AND2X2_74/Y vdd AND2X2
XFILL_12_9_1 gnd vdd FILL
XFILL_14_7_0 gnd vdd FILL
XOAI21X1_313 gnd NOR2X1_192/B INVX1_208/Y gnd AOI21X1_214/A vdd OAI21X1
XINVX1_134 INVX1_134/A gnd INVX1_134/Y vdd INVX1
XNAND2X1_427 INVX1_292/A NOR2X1_246/Y gnd NAND3X1_365/C vdd NAND2X1
XNOR2X1_346 gnd XOR2X1_279/Y gnd NOR2X1_346/Y vdd NOR2X1
XAND2X2_38 gnd OR2X2_49/B gnd NOR3X1_37/C vdd AND2X2
XNAND3X1_259 INVX1_166/A NAND3X1_259/B OR2X2_114/Y gnd AOI21X1_180/C vdd NAND3X1
XFILL_22_4_1 gnd vdd FILL
XBUFX2_260 OR2X2_61/A gnd BUFX2_260/Y vdd BUFX2
XFILL_24_2_0 gnd vdd FILL
XFILL_2_5_1 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XOAI21X1_277 INVX2_58/Y AND2X2_96/B INVX1_181/A gnd OAI21X1_278/B vdd OAI21X1
XNOR2X1_310 gnd NOR2X1_310/B gnd NOR2X1_310/Y vdd NOR2X1
XBUFX4_23 INVX8_1/Y gnd NOR3X1_9/A vdd BUFX4
XNAND2X1_391 AOI21X1_233/A AOI21X1_233/B gnd XOR2X1_197/B vdd NAND2X1
XNAND3X1_223 INVX1_144/A AOI21X1_155/A OR2X2_98/Y gnd NAND3X1_224/C vdd NAND3X1
XBUFX2_224 BUFX2_224/A gnd BUFX2_224/Y vdd BUFX2
XNOR2X1_77 NOR2X1_77/A NOR2X1_76/Y gnd NOR2X1_77/Y vdd NOR2X1
XOAI21X1_241 AND2X2_85/Y NOR2X1_154/Y INVX1_158/Y gnd NAND3X1_253/A vdd OAI21X1
XNAND2X1_355 XOR2X1_179/B NOR2X1_196/Y gnd NAND2X1_355/Y vdd NAND2X1
XINVX2_62 INVX2_62/A gnd INVX2_62/Y vdd INVX2
XNOR2X1_274 gnd XOR2X1_225/Y gnd NOR2X1_274/Y vdd NOR2X1
XNOR2X1_41 NOR2X1_41/A INVX2_18/A gnd XOR2X1_30/B vdd NOR2X1
XNAND3X1_6 NAND3X1_6/A NAND3X1_6/B XNOR2X1_6/B gnd XNOR2X1_7/B vdd NAND3X1
XNAND3X1_187 INVX1_122/A NAND3X1_187/B OR2X2_82/Y gnd NAND3X1_187/Y vdd NAND3X1
XXNOR2X1_226 NOR2X1_410/A bloque_bytes[16] gnd NAND3X1_510/B vdd XNOR2X1
XBUFX2_188 BUFX2_188/A gnd BUFX2_188/Y vdd BUFX2
XINVX2_26 INVX2_26/A gnd INVX2_26/Y vdd INVX2
XOAI21X1_205 NAND2X1_237/Y OAI21X1_205/B AND2X2_72/B gnd XNOR2X1_108/A vdd OAI21X1
XNOR2X1_238 gnd XOR2X1_198/Y gnd NOR2X1_238/Y vdd NOR2X1
XNAND2X1_319 NAND2X1_319/A OR2X2_127/Y gnd OR2X2_128/A vdd NAND2X1
XFILL_21_7_0 gnd vdd FILL
XOR2X2_9 gnd OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XFILL_1_8_0 gnd vdd FILL
XBUFX2_152 XOR2X1_3/A gnd BUFX2_152/Y vdd BUFX2
XCLKBUF1_29 BUFX4_6/Y gnd CLKBUF1_29/Y vdd CLKBUF1
XNAND3X1_151 INVX1_100/A NAND2X1_175/Y OR2X2_66/Y gnd AOI21X1_108/C vdd NAND3X1
XFILL_19_9_1 gnd vdd FILL
XINVX1_567 INVX1_567/A gnd INVX1_567/Y vdd INVX1
XXNOR2X1_190 NOR2X1_309/Y XNOR2X1_190/B gnd XNOR2X1_190/Y vdd XNOR2X1
XFILL_16_2 gnd vdd FILL
XNOR2X1_202 gnd NOR2X1_202/B gnd NOR2X1_202/Y vdd NOR2X1
XNAND2X1_283 NAND2X1_283/A INVX1_163/A gnd INVX1_161/A vdd NAND2X1
XOAI21X1_169 AND2X2_59/Y NOR2X1_112/Y INVX1_113/Y gnd NAND3X1_179/A vdd OAI21X1
XFILL_31_2_0 gnd vdd FILL
XNOR3X1_82 NOR3X1_82/A INVX2_71/Y NOR3X1_82/C gnd NOR3X1_82/Y vdd NOR3X1
XDFFPOSX1_349 INVX1_419/A CLKBUF1_46/Y NAND3X1_516/Y gnd vdd DFFPOSX1
XFILL_29_4_1 gnd vdd FILL
XNAND3X1_115 INVX1_78/A AOI21X1_83/A OR2X2_50/Y gnd AOI21X1_84/C vdd NAND3X1
XFILL_9_5_1 gnd vdd FILL
XINVX1_531 INVX1_531/A gnd INVX1_531/Y vdd INVX1
XBUFX2_116 gnd gnd BUFX2_116/Y vdd BUFX2
XXNOR2X1_76 gnd XOR2X1_72/Y gnd XNOR2X1_77/A vdd XNOR2X1
XXNOR2X1_154 NOR2X1_201/Y XNOR2X1_154/B gnd XNOR2X1_155/A vdd XNOR2X1
XOAI21X1_133 AND2X2_46/Y NOR2X1_90/Y INVX1_90/A gnd AOI21X1_97/A vdd OAI21X1
XNOR2X1_166 INVX1_172/Y NOR2X1_166/B gnd NOR2X1_166/Y vdd NOR2X1
XNAND2X1_247 NAND2X1_247/A NAND2X1_247/B gnd XOR2X1_129/A vdd NAND2X1
XNOR3X1_46 NOR3X1_46/A NOR3X1_46/B NOR3X1_46/C gnd NOR3X1_46/Y vdd NOR3X1
XINVX1_495 bloque_bytes[26] gnd INVX1_495/Y vdd INVX1
XDFFPOSX1_313 XNOR2X1_178/B CLKBUF1_23/Y OR2X2_149/A gnd vdd DFFPOSX1
XXOR2X1_310 vdd gnd gnd OR2X2_1/B vdd XOR2X1
XXNOR2X1_118 BUFX2_161/A XOR2X1_118/Y gnd OR2X2_103/A vdd XNOR2X1
XXNOR2X1_40 gnd XOR2X1_32/Y gnd AOI21X1_69/B vdd XNOR2X1
XNOR2X1_130 gnd OR2X2_91/B gnd NOR2X1_130/Y vdd NOR2X1
XNAND2X1_211 gnd OR2X2_81/B gnd NAND3X1_185/B vdd NAND2X1
XNOR3X1_10 NOR3X1_9/A NOR3X1_10/B NOR3X1_9/C gnd NOR3X1_10/Y vdd NOR3X1
XOAI21X1_638 NOR3X1_98/Y NOR2X1_450/A NAND3X1_533/A gnd NAND2X1_709/B vdd OAI21X1
XOR2X2_98 gnd OR2X2_98/B gnd OR2X2_98/Y vdd OR2X2
XDFFPOSX1_277 INVX1_248/A CLKBUF1_27/Y INVX1_538/Y gnd vdd DFFPOSX1
XINVX1_459 INVX1_459/A gnd INVX1_459/Y vdd INVX1
XFILL_26_9_1 gnd vdd FILL
XXOR2X1_274 XOR2X1_274/A INVX1_422/A gnd INVX1_442/A vdd XOR2X1
XFILL_28_7_0 gnd vdd FILL
XNAND2X1_175 gnd OR2X2_66/B gnd NAND2X1_175/Y vdd NAND2X1
XFILL_8_8_0 gnd vdd FILL
XAOI21X1_73 OAI21X1_99/Y AOI21X1_73/B NOR2X1_73/B gnd INVX2_27/A vdd AOI21X1
XDFFPOSX1_241 XOR2X1_151/B CLKBUF1_26/Y INVX1_528/A gnd vdd DFFPOSX1
XMUX2X1_20 BUFX2_20/A INVX2_10/A MUX2X1_9/S gnd MUX2X1_20/Y vdd MUX2X1
XOR2X2_62 OR2X2_62/A OR2X2_62/B gnd OR2X2_62/Y vdd OR2X2
XOAI21X1_602 INVX1_509/Y bloque_bytes[17] INVX1_510/Y gnd AOI21X1_363/C vdd OAI21X1
XXOR2X1_238 XOR2X1_238/A INVX1_346/A gnd INVX1_366/A vdd XOR2X1
XFILL_36_4_1 gnd vdd FILL
XINVX1_423 INVX1_423/A gnd INVX1_423/Y vdd INVX1
XNAND2X1_716 NAND3X1_546/A OR2X2_162/B gnd OR2X2_160/A vdd NAND2X1
XBUFX2_76 gnd gnd BUFX2_76/Y vdd BUFX2
XNAND3X1_548 NAND3X1_548/A XNOR2X1_254/A XOR2X1_317/B gnd NAND3X1_548/Y vdd NAND3X1
XNAND2X1_139 INVX1_85/A OAI21X1_113/Y gnd OAI21X1_119/A vdd NAND2X1
XAOI21X1_375 INVX1_532/Y bloque_bytes[37] AOI21X1_375/C gnd OAI21X1_611/C vdd AOI21X1
XAOI21X1_37 AOI21X1_37/A AOI21X1_37/B NOR2X1_43/B gnd INVX2_18/A vdd AOI21X1
XOR2X2_26 gnd OR2X2_26/B gnd OR2X2_26/Y vdd OR2X2
XOAI21X1_566 NOR2X1_380/Y AND2X2_158/B BUFX4_33/Y gnd NOR2X1_384/B vdd OAI21X1
XDFFPOSX1_205 INVX1_123/A CLKBUF1_50/Y bloque_bytes[3] gnd vdd DFFPOSX1
XINVX1_387 INVX1_387/A gnd INVX1_387/Y vdd INVX1
XXOR2X1_202 XOR2X1_202/A BUFX2_191/A gnd INVX1_290/A vdd XOR2X1
XNAND2X1_680 INVX1_531/Y INVX1_554/A gnd NAND2X1_680/Y vdd NAND2X1
XAOI21X1_339 INVX2_77/Y NAND2X1_628/Y AOI21X1_339/C gnd AOI21X1_339/Y vdd AOI21X1
XBUFX2_40 gnd gnd BUFX2_40/Y vdd BUFX2
XNAND2X1_103 OR2X2_36/A OR2X2_36/B gnd NAND3X1_84/B vdd NAND2X1
XOAI21X1_85 OAI21X1_85/A OAI21X1_85/B OAI21X1_85/C gnd OAI21X1_85/Y vdd OAI21X1
XFILL_10_2_1 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XNAND3X1_512 XNOR2X1_216/Y NAND3X1_512/B NAND2X1_659/B gnd AOI21X1_388/C vdd NAND3X1
XDFFPOSX1_169 XOR2X1_61/B CLKBUF1_12/Y bloque_bytes[47] gnd vdd DFFPOSX1
XOAI21X1_530 gnd NOR2X1_336/B INVX1_436/A gnd INVX1_439/A vdd OAI21X1
XINVX1_351 INVX1_351/A gnd INVX1_351/Y vdd INVX1
XNAND2X1_644 bloque_bytes[75] bloque_bytes[35] gnd NAND2X1_644/Y vdd NAND2X1
XXOR2X1_166 XOR2X1_166/A INVX1_194/A gnd INVX1_214/A vdd XOR2X1
XNAND2X1_64 gnd OR2X2_19/B gnd NAND3X1_46/B vdd NAND2X1
XNAND3X1_476 INVX1_458/A NAND3X1_476/B INVX2_73/Y gnd OAI21X1_556/B vdd NAND3X1
XAOI21X1_303 AOI21X1_303/A AOI21X1_302/Y INVX1_427/Y gnd AOI21X1_304/A vdd AOI21X1
XFILL_35_7_0 gnd vdd FILL
XOAI21X1_49 AND2X2_17/Y NOR2X1_42/Y INVX1_36/A gnd NAND3X1_49/C vdd OAI21X1
XDFFPOSX1_133 INVX1_24/A CLKBUF1_37/Y bloque_bytes[75] gnd vdd DFFPOSX1
XDFFPOSX1_67 INVX1_476/A CLKBUF1_26/Y AOI21X1_329/Y gnd vdd DFFPOSX1
XFILL_33_9_1 gnd vdd FILL
XXOR2X1_130 XOR2X1_130/A XOR2X1_130/B gnd BUFX2_170/A vdd XOR2X1
XOAI21X1_494 NOR3X1_80/A NOR3X1_80/C INVX2_70/A gnd NOR2X1_313/A vdd OAI21X1
XINVX1_315 INVX1_315/A gnd INVX1_315/Y vdd INVX1
XNAND2X1_608 NAND2X1_608/A NAND2X1_608/B gnd NAND2X1_608/Y vdd NAND2X1
XNAND2X1_28 INVX2_12/Y NAND2X1_28/B gnd XNOR2X1_8/A vdd NAND2X1
XOAI21X1_13 AND2X2_4/Y NOR2X1_20/Y INVX1_13/Y gnd AOI21X1_12/A vdd OAI21X1
XDFFPOSX1_31 INVX1_522/A CLKBUF1_9/Y NOR2X1_361/Y gnd vdd DFFPOSX1
XNAND3X1_440 INVX1_403/Y INVX1_404/Y INVX1_405/Y gnd NAND3X1_440/Y vdd NAND3X1
XAOI21X1_267 INVX1_350/A NAND3X1_401/Y INVX1_345/Y gnd NOR2X1_280/B vdd AOI21X1
XINVX1_279 INVX1_279/A gnd INVX1_279/Y vdd INVX1
XAOI21X1_7 INVX1_7/A INVX4_1/Y AOI21X1_7/C gnd AOI22X1_7/D vdd AOI21X1
XOAI21X1_458 gnd NOR2X1_291/B INVX1_362/A gnd INVX1_364/A vdd OAI21X1
XOR2X2_157 vdd gnd gnd OR2X2_157/Y vdd OR2X2
XXOR2X1_74 XOR2X1_74/A gnd gnd OR2X2_66/B vdd XOR2X1
XNAND2X1_572 NAND2X1_572/A NAND3X1_462/B gnd BUFX2_243/A vdd NAND2X1
XAOI21X1_231 NAND3X1_334/Y AOI21X1_231/B INVX1_256/Y gnd AOI21X1_232/A vdd AOI21X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XNAND3X1_404 INVX1_350/A OAI21X1_444/Y NAND3X1_404/C gnd NAND2X1_486/A vdd NAND3X1
XAND2X2_174 INVX1_481/A INVX1_482/A gnd AND2X2_174/Y vdd AND2X2
XINVX1_243 INVX1_243/A gnd INVX1_243/Y vdd INVX1
XFILL_19_0_0 gnd vdd FILL
XOAI21X1_422 BUFX2_207/A INVX1_328/A INVX1_329/Y gnd NAND3X1_394/B vdd OAI21X1
XNAND3X1_69 NAND3X1_69/A NAND3X1_68/Y NAND3X1_69/C gnd AND2X2_24/A vdd NAND3X1
XXOR2X1_38 XOR2X1_38/A BUFX2_241/A gnd XOR2X1_38/Y vdd XOR2X1
XFILL_17_2_1 gnd vdd FILL
XOR2X2_121 gnd AND2X2_92/B gnd OR2X2_121/Y vdd OR2X2
XNAND2X1_536 INVX1_398/Y NOR2X1_312/Y gnd NAND3X1_437/B vdd NAND2X1
XAOI21X1_195 NOR3X1_55/Y NOR2X1_173/Y NOR2X1_171/A gnd OAI21X1_272/C vdd AOI21X1
XNAND3X1_368 INVX1_288/A OAI21X1_384/Y NAND3X1_363/Y gnd NAND2X1_436/A vdd NAND3X1
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XNAND3X1_33 NAND3X1_35/A NAND3X1_33/B AOI21X1_26/Y gnd AND2X2_12/A vdd NAND3X1
XNOR2X1_419 bloque_bytes[34] INVX1_544/A gnd NOR2X1_419/Y vdd NOR2X1
XOAI21X1_386 NOR2X1_245/Y NOR2X1_244/B AOI22X1_13/C gnd XOR2X1_215/A vdd OAI21X1
XNAND2X1_500 INVX1_362/A NOR2X1_291/Y gnd NAND3X1_412/C vdd NAND2X1
XAND2X2_138 NOR2X1_298/Y INVX1_377/Y gnd NOR3X1_78/A vdd AND2X2
XINVX1_53 OR2X2_32/Y gnd INVX1_53/Y vdd INVX1
XAOI21X1_159 NOR3X1_49/Y NOR2X1_143/Y NOR2X1_141/A gnd OAI21X1_221/C vdd AOI21X1
XNAND3X1_332 INVX2_62/A NAND2X1_382/B NAND3X1_332/C gnd NOR3X1_63/A vdd NAND3X1
XINVX1_171 INVX1_171/A gnd OR2X2_119/B vdd INVX1
XOAI21X1_350 BUFX2_188/A NOR2X1_222/B INVX1_254/A gnd AOI22X1_11/B vdd OAI21X1
XAND2X2_102 AND2X2_102/A INVX1_206/Y gnd NOR3X1_60/A vdd AND2X2
XNOR2X1_383 OR2X2_129/A NOR2X1_383/B gnd NOR2X1_384/A vdd NOR2X1
XNAND2X1_464 NAND3X1_386/Y INVX1_332/A gnd NAND2X1_464/Y vdd NAND2X1
XNAND3X1_296 INVX1_193/A NAND3X1_296/B INVX1_192/Y gnd INVX1_199/A vdd NAND3X1
XAND2X2_75 gnd OR2X2_98/B gnd NOR3X1_50/C vdd AND2X2
XAOI21X1_123 NOR3X1_43/Y NOR2X1_113/Y NOR2X1_111/A gnd OAI21X1_170/C vdd AOI21X1
XINVX1_17 INVX1_17/A gnd OR2X2_7/B vdd INVX1
XFILL_14_7_1 gnd vdd FILL
XFILL_16_5_0 gnd vdd FILL
XOAI21X1_314 BUFX2_181/A XOR2X1_168/Y INVX1_220/A gnd NAND2X1_357/A vdd OAI21X1
XINVX1_135 INVX1_135/A gnd INVX1_135/Y vdd INVX1
XNOR2X1_347 gnd NOR2X1_347/B gnd NOR2X1_347/Y vdd NOR2X1
XNAND2X1_428 INVX1_292/Y NOR2X1_246/Y gnd INVX1_295/A vdd NAND2X1
XAND2X2_39 gnd OR2X2_50/B gnd NOR3X1_38/C vdd AND2X2
XNAND3X1_260 NAND3X1_261/B NAND3X1_260/B AOI21X1_180/C gnd NAND3X1_260/Y vdd NAND3X1
XBUFX2_261 XOR2X1_78/B gnd BUFX2_261/Y vdd BUFX2
XFILL_26_0_0 gnd vdd FILL
XNOR3X1_1 NOR3X1_2/A MUX2X1_1/Y NOR3X1_2/C gnd NOR3X1_1/Y vdd NOR3X1
XFILL_4_3_1 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XOAI21X1_278 OAI21X1_278/A OAI21X1_278/B INVX1_183/Y gnd NAND3X1_292/C vdd OAI21X1
XFILL_24_2_1 gnd vdd FILL
XNAND2X1_392 INVX1_246/A NOR2X1_216/Y gnd AOI21X1_230/B vdd NAND2X1
XBUFX4_24 INVX8_1/Y gnd NOR3X1_2/A vdd BUFX4
XNOR2X1_311 gnd NOR2X1_311/B gnd NOR2X1_311/Y vdd NOR2X1
XNAND3X1_224 NAND3X1_224/A NAND2X1_250/B NAND3X1_224/C gnd NAND2X1_252/A vdd NAND3X1
XBUFX2_225 BUFX2_225/A gnd BUFX2_225/Y vdd BUFX2
XNOR2X1_78 gnd OR2X2_49/B gnd NOR3X1_37/B vdd NOR2X1
XOAI21X1_242 XNOR2X1_125/A NAND2X1_284/Y NOR2X1_155/Y gnd NOR2X1_156/B vdd OAI21X1
XNAND2X1_356 INVX1_220/Y NOR2X1_199/Y gnd NAND2X1_357/B vdd NAND2X1
XINVX2_63 INVX2_63/A gnd INVX2_63/Y vdd INVX2
XNOR2X1_275 gnd NOR2X1_275/B gnd NOR2X1_275/Y vdd NOR2X1
XNAND3X1_188 NAND3X1_189/B NAND3X1_185/Y NAND3X1_187/Y gnd NAND2X1_214/A vdd NAND3X1
XNOR2X1_42 OR2X2_20/A OR2X2_20/B gnd NOR2X1_42/Y vdd NOR2X1
XNAND3X1_7 INVX1_12/A NAND3X1_7/B OR2X2_2/Y gnd NAND3X1_8/C vdd NAND3X1
XBUFX2_189 BUFX2_189/A gnd BUFX2_189/Y vdd BUFX2
XXNOR2X1_227 NOR2X1_411/A bloque_bytes[17] gnd XNOR2X1_227/Y vdd XNOR2X1
XINVX2_27 INVX2_27/A gnd INVX2_27/Y vdd INVX2
XFILL_23_5_0 gnd vdd FILL
XOAI21X1_206 AND2X2_73/Y NOR2X1_134/Y INVX1_136/A gnd NAND3X1_215/B vdd OAI21X1
XNOR2X1_239 gnd NOR2X1_239/B gnd NOR2X1_239/Y vdd NOR2X1
XFILL_3_6_0 gnd vdd FILL
XNAND2X1_320 OR2X2_128/B OR2X2_128/A gnd NAND2X1_321/A vdd NAND2X1
XFILL_21_7_1 gnd vdd FILL
XFILL_1_8_1 gnd vdd FILL
XBUFX2_153 XOR2X1_4/A gnd BUFX2_153/Y vdd BUFX2
XNAND3X1_152 OAI21X1_146/Y NAND3X1_152/B AOI21X1_108/C gnd NAND2X1_176/A vdd NAND3X1
XCLKBUF1_30 BUFX4_3/Y gnd CLKBUF1_30/Y vdd CLKBUF1
XINVX1_568 INVX1_568/A gnd INVX1_568/Y vdd INVX1
XOAI21X1_170 OAI21X1_165/A XNOR2X1_88/B OAI21X1_170/C gnd OAI21X1_170/Y vdd OAI21X1
XXNOR2X1_191 XNOR2X1_190/Y XNOR2X1_191/B gnd INVX1_395/A vdd XNOR2X1
XNOR2X1_203 gnd NOR2X1_203/B gnd AND2X2_107/A vdd NOR2X1
XNAND2X1_284 INVX2_52/A AND2X2_84/Y gnd NAND2X1_284/Y vdd NAND2X1
XFILL_33_0_0 gnd vdd FILL
XFILL_31_2_1 gnd vdd FILL
XDFFPOSX1_350 INVX1_424/A CLKBUF1_19/Y NAND3X1_517/Y gnd vdd DFFPOSX1
XNOR3X1_83 NOR3X1_83/A INVX1_437/A NOR3X1_83/C gnd NOR3X1_83/Y vdd NOR3X1
XBUFX2_117 gnd gnd BUFX2_117/Y vdd BUFX2
XNAND3X1_116 OAI21X1_112/Y OAI21X1_113/C AOI21X1_84/C gnd NAND2X1_138/A vdd NAND3X1
XXNOR2X1_155 XNOR2X1_155/A NAND2X1_357/A gnd INVX1_224/A vdd XNOR2X1
XINVX1_532 bloque_bytes[77] gnd INVX1_532/Y vdd INVX1
XXNOR2X1_77 XNOR2X1_77/A INVX2_35/Y gnd OR2X2_84/A vdd XNOR2X1
XNOR2X1_167 NOR2X1_167/A NOR2X1_166/Y gnd XOR2X1_158/A vdd NOR2X1
XOAI21X1_134 AND2X2_47/Y NOR2X1_92/Y INVX1_91/A gnd OAI21X1_134/Y vdd OAI21X1
XNAND2X1_248 INVX2_47/Y NAND2X1_248/B gnd XNOR2X1_114/B vdd NAND2X1
XNOR3X1_47 INVX1_132/Y NOR3X1_47/B NOR3X1_47/C gnd NOR3X1_47/Y vdd NOR3X1
XINVX1_496 bloque_bytes[27] gnd INVX1_496/Y vdd INVX1
XDFFPOSX1_314 INVX1_339/A CLKBUF1_2/Y INVX1_558/Y gnd vdd DFFPOSX1
XXOR2X1_311 vdd gnd gnd OR2X2_2/B vdd XOR2X1
XXNOR2X1_41 AOI21X1_69/B INVX2_23/Y gnd OR2X2_52/A vdd XNOR2X1
XXNOR2X1_119 XOR2X1_131/Y XOR2X1_119/Y gnd XNOR2X1_120/A vdd XNOR2X1
XNAND2X1_212 OAI21X1_178/Y NAND3X1_185/Y gnd XNOR2X1_96/A vdd NAND2X1
XNOR2X1_131 NOR2X1_131/A INVX2_45/A gnd XOR2X1_120/B vdd NOR2X1
XDFFPOSX1_278 INVX1_253/A CLKBUF1_27/Y INVX1_539/Y gnd vdd DFFPOSX1
XNOR3X1_11 BUFX4_25/Y NOR3X1_11/B BUFX4_21/Y gnd NOR3X1_11/Y vdd NOR3X1
XOAI21X1_639 OAI21X1_639/A XNOR2X1_254/B INVX1_598/A gnd XOR2X1_317/A vdd OAI21X1
XOR2X2_99 gnd OR2X2_99/B gnd OR2X2_99/Y vdd OR2X2
XINVX1_460 INVX1_460/A gnd INVX1_460/Y vdd INVX1
XFILL_30_5_0 gnd vdd FILL
XFILL_28_7_1 gnd vdd FILL
XFILL_8_8_1 gnd vdd FILL
XXOR2X1_275 XOR2X1_275/A BUFX2_228/A gnd NOR2X1_342/B vdd XOR2X1
XNAND2X1_176 NAND2X1_176/A OAI21X1_145/Y gnd XNOR2X1_79/A vdd NAND2X1
XAOI21X1_74 AOI21X1_74/A OR2X2_43/Y INVX1_68/A gnd AOI21X1_74/Y vdd AOI21X1
XDFFPOSX1_242 INVX2_56/A CLKBUF1_21/Y OR2X2_150/B gnd vdd DFFPOSX1
XMUX2X1_21 BUFX2_21/A INVX1_8/A BUFX4_8/Y gnd MUX2X1_21/Y vdd MUX2X1
XOR2X2_63 OR2X2_63/A OR2X2_63/B gnd OR2X2_63/Y vdd OR2X2
XOAI21X1_603 INVX1_512/Y bloque_bytes[18] INVX1_513/Y gnd OAI21X1_603/Y vdd OAI21X1
XINVX1_424 INVX1_424/A gnd INVX1_424/Y vdd INVX1
XXOR2X1_239 XOR2X1_233/Y BUFX2_212/A gnd NOR2X1_294/B vdd XOR2X1
XNAND2X1_717 OR2X2_161/B OR2X2_161/A gnd NAND2X1_718/A vdd NAND2X1
XBUFX2_77 gnd gnd BUFX2_77/Y vdd BUFX2
XNAND3X1_549 INVX1_599/A INVX1_600/A NAND3X1_549/C gnd NAND2X1_722/A vdd NAND3X1
XNAND2X1_140 gnd OR2X2_51/B gnd AOI21X1_86/A vdd NAND2X1
XAOI21X1_376 INVX1_536/Y bloque_bytes[26] AOI21X1_376/C gnd NAND2X1_659/B vdd AOI21X1
XOR2X2_27 gnd OR2X2_27/B gnd OR2X2_27/Y vdd OR2X2
XAOI21X1_38 NAND3X1_46/B OR2X2_19/Y INVX1_35/A gnd NAND3X1_51/C vdd AOI21X1
XDFFPOSX1_206 INVX1_124/A CLKBUF1_50/Y bloque_bytes[4] gnd vdd DFFPOSX1
XOAI21X1_567 NOR2X1_384/A AND2X2_159/B BUFX4_33/Y gnd OAI21X1_567/Y vdd OAI21X1
XINVX1_388 INVX1_388/A gnd INVX1_388/Y vdd INVX1
XBUFX2_41 gnd gnd BUFX2_41/Y vdd BUFX2
XXOR2X1_203 XOR2X1_197/Y BUFX2_192/A gnd XOR2X1_203/Y vdd XOR2X1
XNAND2X1_681 INVX1_533/Y INVX1_555/A gnd NAND2X1_681/Y vdd NAND2X1
XNAND2X1_104 INVX2_24/Y OAI21X1_85/Y gnd OAI21X1_89/A vdd NAND2X1
XAOI21X1_340 INVX1_481/A AND2X2_173/Y OAI21X1_582/Y gnd DFFPOSX1_80/D vdd AOI21X1
XDFFPOSX1_170 INVX2_29/A CLKBUF1_37/Y bloque_bytes[32] gnd vdd DFFPOSX1
XOAI21X1_86 OAI21X1_89/A AOI21X1_65/C AND2X2_30/B gnd OAI21X1_86/Y vdd OAI21X1
XFILL_12_0_1 gnd vdd FILL
XNAND3X1_513 XNOR2X1_217/Y NAND3X1_513/B AOI21X1_393/B gnd NAND3X1_513/Y vdd NAND3X1
XXOR2X1_167 XOR2X1_167/A BUFX2_176/A gnd NOR2X1_198/B vdd XOR2X1
XINVX1_352 INVX1_352/A gnd INVX1_352/Y vdd INVX1
XOAI21X1_531 NOR3X1_83/A INVX1_437/A OAI21X1_537/B gnd NOR2X1_338/A vdd OAI21X1
XNAND2X1_645 NAND2X1_644/Y OR2X2_133/Y gnd NAND2X1_646/B vdd NAND2X1
XOAI21X1_50 AND2X2_17/Y NOR2X1_42/Y INVX1_36/Y gnd NAND3X1_51/A vdd OAI21X1
XNAND2X1_65 OR2X2_20/A OR2X2_20/B gnd NAND3X1_50/B vdd NAND2X1
XNAND3X1_477 INVX1_458/A OAI21X1_552/Y NAND2X1_595/Y gnd NAND3X1_477/Y vdd NAND3X1
XFILL_35_7_1 gnd vdd FILL
XAOI21X1_304 AOI21X1_304/A AOI21X1_304/B AOI21X1_304/C gnd AOI21X1_304/Y vdd AOI21X1
XDFFPOSX1_134 INVX1_25/A CLKBUF1_37/Y bloque_bytes[76] gnd vdd DFFPOSX1
XDFFPOSX1_68 AND2X2_162/B CLKBUF1_26/Y AOI21X1_330/Y gnd vdd DFFPOSX1
XINVX1_316 INVX1_316/A gnd INVX1_316/Y vdd INVX1
XNAND2X1_609 inicio INVX1_486/Y gnd NOR2X1_383/B vdd NAND2X1
XXOR2X1_131 BUFX2_162/A XOR2X1_131/B gnd XOR2X1_131/Y vdd XOR2X1
XOAI21X1_495 gnd XOR2X1_255/Y INVX1_400/Y gnd NAND3X1_438/B vdd OAI21X1
XAOI21X1_268 OAI21X1_441/Y NAND3X1_402/Y INVX1_345/A gnd NOR2X1_280/A vdd AOI21X1
XNAND2X1_29 AND2X2_6/B AND2X2_6/A gnd OAI21X1_18/B vdd NAND2X1
XOAI21X1_14 AND2X2_4/Y NOR2X1_20/Y INVX1_13/A gnd AOI21X1_13/A vdd OAI21X1
XDFFPOSX1_32 INVX1_525/A CLKBUF1_9/Y AND2X2_160/Y gnd vdd DFFPOSX1
XNAND3X1_441 INVX1_405/A INVX1_403/Y INVX1_404/Y gnd NAND3X1_441/Y vdd NAND3X1
XFILL_11_3_0 gnd vdd FILL
XINVX1_280 INVX1_280/A gnd INVX1_280/Y vdd INVX1
XOAI21X1_459 BUFX2_215/A INVX1_366/A INVX1_367/A gnd INVX1_369/A vdd OAI21X1
XAOI21X1_8 INVX1_10/Y target[0] AOI21X1_8/C gnd NAND3X1_4/B vdd AOI21X1
XOR2X2_158 gnd gnd gnd OR2X2_158/Y vdd OR2X2
XXOR2X1_75 XOR2X1_75/A gnd gnd OR2X2_67/B vdd XOR2X1
XNAND2X1_573 INVX1_435/Y NOR2X1_335/Y gnd NAND2X1_573/Y vdd NAND2X1
XAOI21X1_232 AOI21X1_232/A AOI21X1_232/B NAND2X1_393/Y gnd AOI21X1_232/Y vdd AOI21X1
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XNAND3X1_405 AOI22X1_16/B INVX1_352/A INVX1_350/Y gnd NAND2X1_486/B vdd NAND3X1
XAND2X2_1 AND2X2_1/A AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XXOR2X1_39 XOR2X1_39/A XOR2X1_39/B gnd XOR2X1_39/Y vdd XOR2X1
XNAND3X1_70 INVX1_48/Y NAND3X1_72/B OR2X2_29/Y gnd NAND3X1_71/C vdd NAND3X1
XAND2X2_175 AND2X2_175/A AND2X2_175/B gnd AND2X2_175/Y vdd AND2X2
XFILL_19_0_1 gnd vdd FILL
XINVX1_244 INVX1_244/A gnd INVX1_244/Y vdd INVX1
XOAI21X1_423 NOR3X1_71/C OAI21X1_423/B INVX1_332/A gnd NOR2X1_269/A vdd OAI21X1
XOR2X2_122 gnd OR2X2_122/B gnd OR2X2_122/Y vdd OR2X2
XNAND2X1_537 INVX1_401/A NAND3X1_437/B gnd INVX1_399/A vdd NAND2X1
XAOI21X1_196 AOI21X1_196/A OR2X2_124/Y INVX1_179/A gnd OR2X2_126/B vdd AOI21X1
XNAND3X1_369 INVX1_299/Y INVX1_298/A AOI21X1_250/B gnd AND2X2_121/B vdd NAND3X1
XINVX1_208 INVX1_208/A gnd INVX1_208/Y vdd INVX1
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XOAI21X1_387 BUFX2_200/A XOR2X1_203/Y INVX1_292/Y gnd NAND3X1_365/B vdd OAI21X1
XNAND3X1_34 INVX1_26/Y NAND3X1_34/B OR2X2_13/Y gnd NAND3X1_35/C vdd NAND3X1
XNOR2X1_420 bloque_bytes[35] INVX1_571/A gnd NOR2X1_420/Y vdd NOR2X1
XNAND2X1_501 INVX1_362/Y NOR2X1_291/Y gnd NAND2X1_501/Y vdd NAND2X1
XAND2X2_139 NOR2X1_299/Y INVX1_378/Y gnd NOR3X1_78/C vdd AND2X2
XAOI21X1_160 NAND3X1_228/B OR2X2_100/Y INVX1_146/A gnd OR2X2_102/B vdd AOI21X1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XFILL_7_1 gnd vdd FILL
XNAND3X1_333 INVX1_249/A NAND2X1_385/B INVX2_62/Y gnd OAI21X1_347/B vdd NAND3X1
XNOR2X1_384 NOR2X1_384/A NOR2X1_384/B gnd NOR2X1_384/Y vdd NOR2X1
XINVX1_172 INVX1_172/A gnd INVX1_172/Y vdd INVX1
XAND2X2_103 AND2X2_103/A INVX1_207/Y gnd NOR3X1_60/C vdd AND2X2
XOAI21X1_351 gnd XOR2X1_182/Y INVX1_246/Y gnd AOI21X1_230/A vdd OAI21X1
XNAND2X1_465 INVX1_330/A NOR2X1_270/Y gnd NAND3X1_391/C vdd NAND2X1
XNAND3X1_297 INVX1_194/Y INVX1_195/Y INVX1_196/Y gnd AOI21X1_203/B vdd NAND3X1
XFILL_18_3_0 gnd vdd FILL
XAND2X2_76 gnd OR2X2_99/B gnd AND2X2_76/Y vdd AND2X2
XAOI21X1_124 NAND3X1_176/B OR2X2_76/Y INVX1_113/A gnd OR2X2_78/B vdd AOI21X1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XFILL_16_5_1 gnd vdd FILL
XOAI21X1_315 OAI21X1_315/A INVX1_223/A INVX1_222/Y gnd AND2X2_105/A vdd OAI21X1
XINVX1_136 INVX1_136/A gnd INVX1_136/Y vdd INVX1
XNAND2X1_429 NAND3X1_365/Y AOI21X1_249/B gnd XOR2X1_215/B vdd NAND2X1
XNOR2X1_348 gnd NOR2X1_348/B gnd NOR2X1_348/Y vdd NOR2X1
XAND2X2_40 gnd OR2X2_51/B gnd AND2X2_40/Y vdd AND2X2
XBUFX2_262 BUFX2_262/A gnd BUFX2_262/Y vdd BUFX2
XNAND3X1_261 AOI21X1_180/C NAND3X1_261/B NOR3X1_53/Y gnd INVX1_173/A vdd NAND3X1
XFILL_26_0_1 gnd vdd FILL
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XFILL_6_1_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd NOR3X1_42/A vdd INVX1
XOAI21X1_279 NOR2X1_177/A INVX1_185/Y INVX1_186/Y gnd NAND2X1_323/B vdd OAI21X1
XBUFX4_25 INVX8_1/Y gnd BUFX4_25/Y vdd BUFX4
XNAND2X1_393 XOR2X1_197/B NOR2X1_220/Y gnd NAND2X1_393/Y vdd NAND2X1
XNOR2X1_312 gnd XOR2X1_254/Y gnd NOR2X1_312/Y vdd NOR2X1
XNOR2X1_79 gnd OR2X2_50/B gnd NOR2X1_79/Y vdd NOR2X1
XNAND3X1_225 NAND3X1_224/C NAND3X1_224/A NOR3X1_49/Y gnd INVX1_151/A vdd NAND3X1
XBUFX2_226 BUFX2_226/A gnd BUFX2_226/Y vdd BUFX2
XFILL_15_8_0 gnd vdd FILL
XOAI21X1_243 INVX2_52/Y AND2X2_84/B INVX1_159/A gnd OAI21X1_243/Y vdd OAI21X1
XINVX2_64 INVX2_64/A gnd INVX2_64/Y vdd INVX2
XNOR2X1_276 gnd NOR2X1_276/B gnd NOR2X1_276/Y vdd NOR2X1
XNAND2X1_357 NAND2X1_357/A NAND2X1_357/B gnd NOR2X1_200/B vdd NAND2X1
XNAND3X1_189 NAND3X1_187/Y NAND3X1_189/B NOR3X1_45/Y gnd INVX1_129/A vdd NAND3X1
XBUFX2_190 BUFX2_190/A gnd BUFX2_190/Y vdd BUFX2
XNOR2X1_43 NOR2X1_43/A NOR2X1_43/B gnd NOR2X1_43/Y vdd NOR2X1
XNAND3X1_8 NAND3X1_8/A NAND3X1_6/A NAND3X1_8/C gnd NAND3X1_8/Y vdd NAND3X1
XXNOR2X1_228 INVX1_537/A bloque_bytes[18] gnd NAND3X1_512/B vdd XNOR2X1
XOAI21X1_207 AND2X2_73/Y NOR2X1_134/Y INVX1_136/Y gnd NAND3X1_217/A vdd OAI21X1
XFILL_5_4_0 gnd vdd FILL
XINVX2_28 INVX2_28/A gnd INVX2_28/Y vdd INVX2
XNAND2X1_321 NAND2X1_321/A INVX1_185/A gnd INVX1_183/A vdd NAND2X1
XFILL_23_5_1 gnd vdd FILL
XNOR2X1_240 gnd XOR2X1_200/Y gnd NOR2X1_240/Y vdd NOR2X1
XFILL_25_3_0 gnd vdd FILL
XFILL_3_6_1 gnd vdd FILL
XBUFX2_154 XOR2X1_5/A gnd BUFX2_154/Y vdd BUFX2
XNAND3X1_153 AOI21X1_108/C OAI21X1_146/Y NOR3X1_41/Y gnd INVX1_107/A vdd NAND3X1
XCLKBUF1_31 BUFX4_1/Y gnd CLKBUF1_31/Y vdd CLKBUF1
XINVX1_569 INVX1_569/A gnd INVX1_569/Y vdd INVX1
XOAI21X1_171 XNOR2X1_89/A AOI21X1_125/C AND2X2_60/B gnd XNOR2X1_90/A vdd OAI21X1
XFILL_33_0_1 gnd vdd FILL
XXNOR2X1_192 NOR2X1_314/A XNOR2X1_192/B gnd BUFX2_234/A vdd XNOR2X1
XNOR2X1_204 gnd NOR2X1_204/B gnd NOR2X1_204/Y vdd NOR2X1
XNAND2X1_285 NAND2X1_285/A NAND2X1_285/B gnd XOR2X1_149/A vdd NAND2X1
XNAND3X1_117 AOI21X1_84/C OAI21X1_112/Y NOR3X1_37/Y gnd INVX1_85/A vdd NAND3X1
XINVX1_533 INVX1_533/A gnd INVX1_533/Y vdd INVX1
XDFFPOSX1_351 INVX1_425/A CLKBUF1_2/Y NAND3X1_518/Y gnd vdd DFFPOSX1
XNOR3X1_84 NOR3X1_84/A INVX2_72/Y NOR3X1_84/C gnd NOR3X1_84/Y vdd NOR3X1
XBUFX2_118 gnd gnd BUFX2_118/Y vdd BUFX2
XXNOR2X1_156 NOR2X1_206/A NAND2X1_369/Y gnd BUFX2_194/A vdd XNOR2X1
XXNOR2X1_78 XNOR2X1_78/A XNOR2X1_78/B gnd OR2X2_85/A vdd XNOR2X1
XNOR2X1_168 gnd AND2X2_92/B gnd NOR3X1_55/B vdd NOR2X1
XOAI21X1_135 AND2X2_47/Y NOR2X1_92/Y INVX1_91/Y gnd OAI21X1_135/Y vdd OAI21X1
XNAND2X1_249 gnd OR2X2_97/B gnd NAND2X1_249/Y vdd NAND2X1
XNOR3X1_48 INVX1_133/Y NOR3X1_48/B NOR3X1_48/C gnd NOR3X1_48/Y vdd NOR3X1
XINVX1_497 bloque_bytes[28] gnd INVX1_497/Y vdd INVX1
XFILL_22_8_0 gnd vdd FILL
XDFFPOSX1_315 INVX1_340/A CLKBUF1_8/Y INVX1_560/Y gnd vdd DFFPOSX1
XFILL_2_9_0 gnd vdd FILL
XXOR2X1_312 vdd vdd gnd OR2X2_3/B vdd XOR2X1
XXNOR2X1_42 NAND2X1_98/Y NAND3X1_78/C gnd OR2X2_53/A vdd XNOR2X1
XXNOR2X1_120 XNOR2X1_120/A OR2X2_103/Y gnd INVX1_153/A vdd XNOR2X1
XNAND2X1_213 gnd OR2X2_82/B gnd NAND3X1_187/B vdd NAND2X1
XNOR2X1_132 OR2X2_92/A OR2X2_92/B gnd NOR2X1_132/Y vdd NOR2X1
XDFFPOSX1_279 INVX1_254/A CLKBUF1_27/Y INVX1_540/Y gnd vdd DFFPOSX1
XNOR3X1_12 BUFX4_25/Y MUX2X1_12/Y BUFX4_21/Y gnd NOR3X1_12/Y vdd NOR3X1
XFILL_32_3_0 gnd vdd FILL
XOAI21X1_640 AND2X2_195/Y NOR2X1_447/Y INVX1_592/Y gnd AOI21X1_395/A vdd OAI21X1
XINVX1_461 INVX1_461/A gnd INVX1_461/Y vdd INVX1
XXOR2X1_276 XOR2X1_276/A BUFX2_229/A gnd NOR2X1_343/B vdd XOR2X1
XFILL_30_5_1 gnd vdd FILL
XNAND2X1_177 INVX1_107/A NAND2X1_177/B gnd OAI21X1_153/A vdd NAND2X1
XAOI21X1_75 NOR3X1_35/Y NOR2X1_73/Y NOR2X1_71/A gnd AOI21X1_75/Y vdd AOI21X1
XOAI21X1_604 INVX1_515/Y bloque_bytes[19] INVX1_516/Y gnd AOI21X1_365/C vdd OAI21X1
XOR2X2_64 OR2X2_64/A OR2X2_64/B gnd OR2X2_64/Y vdd OR2X2
XDFFPOSX1_243 INVX1_176/A CLKBUF1_2/Y OR2X2_151/B gnd vdd DFFPOSX1
XMUX2X1_22 BUFX2_22/A INVX1_7/A BUFX4_8/Y gnd NOR3X1_22/B vdd MUX2X1
XINVX1_425 INVX1_425/A gnd INVX1_425/Y vdd INVX1
XNAND2X1_718 NAND2X1_718/A OR2X2_161/Y gnd OR2X2_162/A vdd NAND2X1
XXOR2X1_240 XOR2X1_240/A BUFX2_213/A gnd XOR2X1_240/Y vdd XOR2X1
XNAND2X1_141 OR2X2_52/A OR2X2_52/B gnd AOI21X1_88/A vdd NAND2X1
XAOI21X1_377 INVX1_542/Y bloque_bytes[31] AOI21X1_377/C gnd AOI21X1_393/B vdd AOI21X1
XBUFX2_78 gnd gnd BUFX2_78/Y vdd BUFX2
XDFFPOSX1_207 INVX1_125/A CLKBUF1_50/Y bloque_bytes[5] gnd vdd DFFPOSX1
XOR2X2_28 OR2X2_28/A OR2X2_28/B gnd OR2X2_28/Y vdd OR2X2
XAOI21X1_39 NOR3X1_29/Y NOR2X1_43/Y NOR2X1_41/A gnd OAI21X1_51/C vdd AOI21X1
XOAI21X1_568 NAND2X1_611/Y INVX2_74/Y INVX8_2/A gnd OAI21X1_568/Y vdd OAI21X1
XFILL_20_1 gnd vdd FILL
XINVX1_389 INVX1_389/A gnd INVX1_389/Y vdd INVX1
XBUFX2_42 gnd gnd BUFX2_42/Y vdd BUFX2
XXOR2X1_204 AND2X2_113/Y BUFX2_193/A gnd XOR2X1_204/Y vdd XOR2X1
XNAND2X1_682 INVX1_548/Y INVX1_556/A gnd NAND2X1_682/Y vdd NAND2X1
XFILL_29_8_0 gnd vdd FILL
XNAND2X1_105 AND2X2_30/B AND2X2_30/A gnd AOI21X1_65/C vdd NAND2X1
XAOI21X1_341 OAI21X1_583/Y AOI21X1_341/B BUFX4_17/Y gnd DFFPOSX1_81/D vdd AOI21X1
XFILL_9_9_0 gnd vdd FILL
XNAND3X1_514 INVX1_574/Y XNOR2X1_234/Y INVX1_546/A gnd NAND3X1_514/Y vdd NAND3X1
XDFFPOSX1_171 INVX1_77/A CLKBUF1_1/Y bloque_bytes[33] gnd vdd DFFPOSX1
XOAI21X1_87 AND2X2_31/Y NOR2X1_64/Y INVX1_59/A gnd OAI21X1_87/Y vdd OAI21X1
XXOR2X1_168 XOR2X1_168/A BUFX2_177/A gnd XOR2X1_168/Y vdd XOR2X1
XINVX1_353 INVX1_353/A gnd INVX1_353/Y vdd INVX1
XOAI21X1_532 NOR3X1_84/A NOR3X1_84/C INVX2_72/A gnd NOR2X1_337/A vdd OAI21X1
XNAND2X1_646 INVX1_503/Y NAND2X1_646/B gnd OR2X2_152/B vdd NAND2X1
XNAND2X1_66 INVX2_18/Y OAI21X1_51/Y gnd OAI21X1_55/A vdd NAND2X1
XOAI21X1_51 OAI21X1_46/A OAI21X1_46/B OAI21X1_51/C gnd OAI21X1_51/Y vdd OAI21X1
XDFFPOSX1_69 AND2X2_163/B CLKBUF1_30/Y NOR2X1_392/Y gnd vdd DFFPOSX1
XNAND3X1_478 INVX1_459/A AOI21X1_317/B INVX1_458/Y gnd INVX1_465/A vdd NAND3X1
XAOI21X1_305 NAND2X1_562/A NAND2X1_562/B AOI21X1_305/C gnd OAI21X1_525/C vdd AOI21X1
XDFFPOSX1_135 INVX1_26/A CLKBUF1_5/Y bloque_bytes[77] gnd vdd DFFPOSX1
XOAI21X1_496 gnd XOR2X1_255/Y INVX1_400/A gnd INVX1_402/A vdd OAI21X1
XINVX1_317 INVX1_317/A gnd INVX1_317/Y vdd INVX1
XNAND2X1_610 INVX1_472/A AND2X2_158/B gnd OR2X2_129/A vdd NAND2X1
XXOR2X1_132 AND2X2_89/A gnd gnd XOR2X1_132/Y vdd XOR2X1
XAOI21X1_269 INVX1_345/A NAND2X1_482/Y INVX1_344/Y gnd NOR3X1_73/C vdd AOI21X1
XNAND2X1_30 vdd OR2X2_5/B gnd NAND3X1_16/B vdd NAND2X1
XOAI21X1_15 AND2X2_5/Y NOR2X1_22/Y INVX1_14/A gnd OAI21X1_15/Y vdd OAI21X1
XDFFPOSX1_33 INVX1_528/A CLKBUF1_20/Y NOR2X1_362/Y gnd vdd DFFPOSX1
XNAND3X1_442 INVX1_407/A NAND3X1_440/Y INVX1_402/Y gnd AOI22X1_19/C vdd NAND3X1
XXOR2X1_76 XOR2X1_76/A OR2X2_60/A gnd OR2X2_68/B vdd XOR2X1
XFILL_11_3_1 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XINVX1_281 INVX1_281/A gnd INVX1_281/Y vdd INVX1
XOAI21X1_460 BUFX2_215/A INVX1_366/A INVX1_367/Y gnd NAND3X1_420/B vdd OAI21X1
XAOI21X1_9 AOI21X1_9/A AOI22X1_7/Y NOR2X1_16/Y gnd AOI21X1_9/Y vdd AOI21X1
XOR2X2_159 gnd gnd gnd OR2X2_159/Y vdd OR2X2
XNAND2X1_574 INVX1_436/Y NOR2X1_336/Y gnd NAND2X1_574/Y vdd NAND2X1
XAOI21X1_233 AOI21X1_233/A AOI21X1_233/B NAND2X1_398/Y gnd AOI21X1_233/Y vdd AOI21X1
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XNAND3X1_406 INVX1_342/Y NAND3X1_399/Y NOR3X1_74/Y gnd AOI21X1_272/B vdd NAND3X1
XAND2X2_2 gnd OR2X2_1/B gnd AND2X2_2/Y vdd AND2X2
XINVX1_245 INVX1_245/A gnd INVX1_245/Y vdd INVX1
XFILL_36_8_0 gnd vdd FILL
XNAND3X1_71 NAND3X1_69/A NAND3X1_71/B NAND3X1_71/C gnd AOI21X1_53/A vdd NAND3X1
XXOR2X1_40 XOR2X1_40/A XOR2X1_40/B gnd XOR2X1_61/A vdd XOR2X1
XAND2X2_176 bloque_bytes[53] bloque_bytes[13] gnd AND2X2_176/Y vdd AND2X2
XNAND2X1_538 INVX1_400/A NOR2X1_315/Y gnd NAND3X1_438/C vdd NAND2X1
XOAI21X1_424 NOR2X1_269/Y NOR2X1_268/B AOI22X1_15/C gnd XOR2X1_233/A vdd OAI21X1
XAOI21X1_197 AOI21X1_197/A AOI21X1_197/B OAI21X1_273/B gnd NAND3X1_290/B vdd AOI21X1
XOR2X2_123 gnd OR2X2_123/B gnd OR2X2_123/Y vdd OR2X2
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XNAND3X1_370 INVX1_297/Y INVX1_300/Y AND2X2_121/A gnd NAND3X1_370/Y vdd NAND3X1
XINVX1_209 NOR3X1_59/B gnd INVX1_209/Y vdd INVX1
XOAI21X1_388 BUFX2_200/A XOR2X1_203/Y INVX1_292/A gnd AOI22X1_13/B vdd OAI21X1
XAND2X2_140 AND2X2_140/A NOR3X1_77/A gnd BUFX2_228/A vdd AND2X2
XNAND3X1_35 NAND3X1_35/A NAND3X1_35/B NAND3X1_35/C gnd AOI21X1_29/A vdd NAND3X1
XNOR2X1_421 bloque_bytes[36] INVX1_572/A gnd NOR2X1_421/Y vdd NOR2X1
XNAND2X1_502 NAND3X1_419/B INVX1_370/A gnd XNOR2X1_184/B vdd NAND2X1
XFILL_10_6_0 gnd vdd FILL
XAOI21X1_161 AOI21X1_161/A AOI21X1_161/B OAI21X1_222/B gnd NAND3X1_236/B vdd AOI21X1
XNAND3X1_334 INVX1_249/A OAI21X1_343/Y NAND3X1_334/C gnd NAND3X1_334/Y vdd NAND3X1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XFILL_7_2 gnd vdd FILL
XNOR2X1_385 INVX4_2/Y NOR2X1_385/B gnd NOR2X1_385/Y vdd NOR2X1
XINVX1_173 INVX1_173/A gnd INVX1_173/Y vdd INVX1
XOAI21X1_352 BUFX2_189/A NOR2X1_223/B INVX1_258/A gnd XNOR2X1_163/B vdd OAI21X1
XAND2X2_104 AND2X2_104/A NOR3X1_59/A gnd BUFX2_188/A vdd AND2X2
XFILL_20_1_0 gnd vdd FILL
XNAND2X1_466 INVX1_330/Y NOR2X1_270/Y gnd INVX1_333/A vdd NAND2X1
XFILL_0_2_0 gnd vdd FILL
XNAND3X1_298 INVX1_196/A INVX1_194/Y INVX1_195/Y gnd AOI21X1_204/B vdd NAND3X1
XAND2X2_77 AND2X2_77/A AND2X2_77/B gnd AND2X2_77/Y vdd AND2X2
XFILL_18_3_1 gnd vdd FILL
XAOI21X1_125 NAND3X1_179/Y NAND3X1_181/Y AOI21X1_125/C gnd NAND3X1_182/B vdd AOI21X1
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XOAI21X1_316 NOR2X1_197/A NOR3X1_59/Y OAI21X1_316/C gnd AOI21X1_218/B vdd OAI21X1
XINVX1_137 OR2X2_94/Y gnd INVX1_137/Y vdd INVX1
XNAND2X1_430 INVX1_284/A NOR2X1_240/Y gnd AOI21X1_246/B vdd NAND2X1
XNOR2X1_349 NOR2X1_349/A INVX1_456/Y gnd NOR2X1_349/Y vdd NOR2X1
XAND2X2_41 OR2X2_52/A OR2X2_52/B gnd AND2X2_41/Y vdd AND2X2
XNOR3X1_3 NOR3X1_3/A MUX2X1_3/Y NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XNAND3X1_262 INVX1_167/A NAND3X1_262/B OR2X2_115/Y gnd AOI21X1_180/B vdd NAND3X1
XBUFX2_263 OR2X2_68/A gnd BUFX2_263/Y vdd BUFX2
XINVX1_101 INVX1_101/A gnd INVX1_101/Y vdd INVX1
XOAI21X1_280 gnd NOR2X1_178/B INVX1_187/A gnd NAND2X1_325/A vdd OAI21X1
XBUFX4_26 INVX8_1/Y gnd NOR3X1_3/A vdd BUFX4
XNAND2X1_394 INVX1_258/Y NOR2X1_223/Y gnd NAND2X1_395/B vdd NAND2X1
XNOR2X1_313 NOR2X1_313/A INVX1_399/Y gnd NOR2X1_314/B vdd NOR2X1
XNAND3X1_226 INVX1_145/A NAND3X1_227/B OR2X2_99/Y gnd AOI21X1_156/B vdd NAND3X1
XNOR2X1_80 gnd OR2X2_51/B gnd NOR2X1_80/Y vdd NOR2X1
XFILL_17_6_0 gnd vdd FILL
XBUFX2_227 INVX1_422/A gnd BUFX2_227/Y vdd BUFX2
XFILL_15_8_1 gnd vdd FILL
XOAI21X1_244 OAI21X1_244/A OAI21X1_243/Y INVX1_161/Y gnd NAND3X1_256/C vdd OAI21X1
XINVX2_65 INVX2_65/A gnd INVX2_65/Y vdd INVX2
XNOR2X1_277 NOR2X1_277/A INVX1_342/Y gnd NOR2X1_278/B vdd NOR2X1
XNAND2X1_358 INVX1_219/Y NOR2X1_200/B gnd NAND2X1_359/A vdd NAND2X1
XNAND3X1_190 INVX1_123/A NAND2X1_216/Y OR2X2_83/Y gnd NAND3X1_190/Y vdd NAND3X1
XNAND3X1_9 NAND3X1_8/C NAND3X1_8/A NOR3X1_25/Y gnd INVX1_19/A vdd NAND3X1
XBUFX2_191 BUFX2_191/A gnd BUFX2_191/Y vdd BUFX2
XNOR2X1_44 OR2X2_21/A OR2X2_21/B gnd NOR2X1_44/Y vdd NOR2X1
XXNOR2X1_229 AOI21X1_353/C bloque_bytes[19] gnd AND2X2_183/B vdd XNOR2X1
XOAI21X1_208 NAND2X1_237/Y AOI21X1_154/C NOR2X1_135/Y gnd NOR2X1_136/B vdd OAI21X1
XFILL_25_3_1 gnd vdd FILL
XFILL_27_1_0 gnd vdd FILL
XINVX2_29 INVX2_29/A gnd INVX2_29/Y vdd INVX2
XFILL_5_4_1 gnd vdd FILL
XFILL_7_2_0 gnd vdd FILL
XNAND2X1_322 INVX2_58/A AND2X2_96/Y gnd NAND2X1_322/Y vdd NAND2X1
XNOR2X1_241 NOR2X1_241/A INVX1_285/Y gnd NOR2X1_242/B vdd NOR2X1
XNAND3X1_154 INVX1_101/A AOI21X1_110/A OR2X2_67/Y gnd NAND3X1_154/Y vdd NAND3X1
XINVX1_570 INVX1_570/A gnd INVX1_570/Y vdd INVX1
XCLKBUF1_32 BUFX4_5/Y gnd CLKBUF1_32/Y vdd CLKBUF1
XBUFX2_155 OR2X2_92/A gnd BUFX2_155/Y vdd BUFX2
XXNOR2X1_193 NOR2X1_317/Y NOR2X1_316/Y gnd XOR2X1_274/A vdd XNOR2X1
XNOR2X1_205 NOR2X1_205/A INVX1_228/Y gnd NOR2X1_206/B vdd NOR2X1
XOAI21X1_172 AND2X2_61/Y NOR2X1_114/Y INVX1_114/A gnd OAI21X1_172/Y vdd OAI21X1
XNAND2X1_286 INVX2_53/Y XNOR2X1_131/A gnd NAND3X1_258/C vdd NAND2X1
XNOR3X1_85 NOR3X1_85/A INVX1_456/A NOR3X1_85/C gnd NOR3X1_85/Y vdd NOR3X1
XNAND3X1_118 INVX1_79/A AOI21X1_86/A OR2X2_51/Y gnd AOI21X1_84/B vdd NAND3X1
XBUFX2_119 gnd gnd BUFX2_119/Y vdd BUFX2
XINVX1_534 INVX1_534/A gnd INVX1_534/Y vdd INVX1
XDFFPOSX1_352 INVX1_429/A CLKBUF1_22/Y NAND3X1_519/Y gnd vdd DFFPOSX1
XXNOR2X1_79 XNOR2X1_79/A XNOR2X1_79/B gnd XOR2X1_94/A vdd XNOR2X1
XBUFX4_1 clk gnd BUFX4_1/Y vdd BUFX4
XXNOR2X1_157 NOR2X1_209/Y NOR2X1_208/Y gnd XOR2X1_193/A vdd XNOR2X1
XNAND2X1_250 NAND2X1_250/A NAND2X1_250/B gnd XNOR2X1_114/A vdd NAND2X1
XNOR2X1_169 gnd OR2X2_122/B gnd NOR3X1_56/B vdd NOR2X1
XOAI21X1_136 OAI21X1_131/A XNOR2X1_70/B AOI21X1_99/Y gnd NAND3X1_146/C vdd OAI21X1
XNOR3X1_49 INVX1_143/Y NOR3X1_49/B AND2X2_74/Y gnd NOR3X1_49/Y vdd NOR3X1
XFILL_24_6_0 gnd vdd FILL
XDFFPOSX1_316 INVX1_341/A CLKBUF1_39/Y INVX1_561/Y gnd vdd DFFPOSX1
XFILL_4_7_0 gnd vdd FILL
XINVX1_498 bloque_bytes[29] gnd INVX1_498/Y vdd INVX1
XFILL_22_8_1 gnd vdd FILL
XFILL_2_9_1 gnd vdd FILL
XXOR2X1_313 vdd gnd gnd OR2X2_4/B vdd XOR2X1
XXNOR2X1_43 XNOR2X1_43/A OAI21X1_85/B gnd XOR2X1_54/A vdd XNOR2X1
XOAI21X1_100 AND2X2_35/Y NOR2X1_72/Y INVX1_69/A gnd OAI21X1_100/Y vdd OAI21X1
XXNOR2X1_121 gnd XOR2X1_122/Y gnd XNOR2X1_122/A vdd XNOR2X1
XNAND2X1_214 NAND2X1_214/A OAI21X1_179/Y gnd XNOR2X1_97/A vdd NAND2X1
XNOR2X1_133 NOR2X1_133/A NOR3X1_48/Y gnd NOR2X1_133/Y vdd NOR2X1
XFILL_34_1_0 gnd vdd FILL
XDFFPOSX1_280 INVX1_258/A CLKBUF1_31/Y INVX1_541/Y gnd vdd DFFPOSX1
XINVX1_462 INVX1_462/A gnd INVX1_462/Y vdd INVX1
XNOR3X1_13 BUFX4_27/Y NOR3X1_13/B BUFX4_20/Y gnd NOR3X1_13/Y vdd NOR3X1
XFILL_32_3_1 gnd vdd FILL
XOAI21X1_641 AND2X2_195/Y NOR2X1_447/Y INVX1_592/A gnd AOI21X1_396/A vdd OAI21X1
XXOR2X1_277 XOR2X1_277/A BUFX2_230/A gnd NOR2X1_345/B vdd XOR2X1
XNAND2X1_178 gnd OR2X2_67/B gnd AOI21X1_110/A vdd NAND2X1
XAOI21X1_76 AOI21X1_76/A OR2X2_44/Y INVX1_69/A gnd OR2X2_46/B vdd AOI21X1
XOAI21X1_605 INVX1_518/Y bloque_bytes[20] INVX1_519/Y gnd AOI21X1_366/C vdd OAI21X1
XDFFPOSX1_244 INVX1_177/A CLKBUF1_21/Y OR2X2_139/A gnd vdd DFFPOSX1
XOR2X2_65 gnd OR2X2_65/B gnd OR2X2_65/Y vdd OR2X2
XMUX2X1_23 BUFX2_23/A INVX1_6/A BUFX4_8/Y gnd NOR3X1_23/B vdd MUX2X1
XINVX1_426 INVX1_426/A gnd INVX1_426/Y vdd INVX1
XNAND2X1_719 OR2X2_162/B OR2X2_162/A gnd NAND2X1_720/A vdd NAND2X1
XBUFX2_79 gnd gnd BUFX2_79/Y vdd BUFX2
XXOR2X1_241 XOR2X1_241/A BUFX2_214/A gnd XOR2X1_241/Y vdd XOR2X1
XNAND2X1_142 INVX2_30/Y NAND3X1_128/C gnd XNOR2X1_62/A vdd NAND2X1
XAOI21X1_378 INVX1_547/Y bloque_bytes[38] OAI21X1_621/Y gnd AOI21X1_378/Y vdd AOI21X1
XAOI21X1_40 NAND3X1_50/B OR2X2_20/Y INVX1_36/A gnd OR2X2_22/B vdd AOI21X1
XDFFPOSX1_208 INVX1_127/A CLKBUF1_47/Y bloque_bytes[6] gnd vdd DFFPOSX1
XOR2X2_29 OR2X2_29/A OR2X2_29/B gnd OR2X2_29/Y vdd OR2X2
XOAI21X1_569 NAND2X1_611/Y INVX2_74/Y INVX1_473/Y gnd NAND2X1_612/B vdd OAI21X1
XFILL_20_2 gnd vdd FILL
XXOR2X1_205 XOR2X1_205/A BUFX2_194/A gnd XOR2X1_205/Y vdd XOR2X1
XINVX1_390 INVX1_390/A gnd INVX1_390/Y vdd INVX1
XNAND2X1_683 INVX1_558/A XNOR2X1_235/Y gnd NAND2X1_683/Y vdd NAND2X1
XFILL_31_6_0 gnd vdd FILL
XBUFX2_43 gnd gnd BUFX2_43/Y vdd BUFX2
XFILL_29_8_1 gnd vdd FILL
XNAND2X1_106 OR2X2_37/A OR2X2_37/B gnd NAND3X1_88/B vdd NAND2X1
XOAI21X1_88 AND2X2_31/Y NOR2X1_64/Y INVX1_59/Y gnd NAND3X1_91/A vdd OAI21X1
XFILL_9_9_1 gnd vdd FILL
XAOI21X1_342 INVX2_78/A NOR3X1_90/Y AOI21X1_342/C gnd AOI21X1_342/Y vdd AOI21X1
XNAND3X1_515 INVX1_575/Y INVX1_549/Y AOI21X1_378/Y gnd NAND2X1_688/B vdd NAND3X1
XDFFPOSX1_172 INVX1_78/A CLKBUF1_1/Y bloque_bytes[34] gnd vdd DFFPOSX1
XOAI21X1_533 gnd NOR2X1_339/B INVX1_438/Y gnd OAI21X1_533/Y vdd OAI21X1
XINVX1_354 INVX1_354/A gnd INVX1_354/Y vdd INVX1
XXOR2X1_169 XOR2X1_169/A BUFX2_178/A gnd NOR2X1_201/B vdd XOR2X1
XNAND2X1_647 bloque_bytes[76] bloque_bytes[36] gnd NAND2X1_647/Y vdd NAND2X1
XAOI21X1_306 INVX1_432/Y OAI21X1_525/Y INVX1_431/A gnd AOI21X1_306/Y vdd AOI21X1
XOAI21X1_52 OAI21X1_55/A OAI21X1_52/B AND2X2_18/B gnd OAI21X1_52/Y vdd OAI21X1
XNAND2X1_67 AND2X2_18/B AND2X2_18/A gnd OAI21X1_52/B vdd NAND2X1
XDFFPOSX1_70 INVX1_477/A CLKBUF1_26/Y NOR3X1_87/Y gnd vdd DFFPOSX1
XNAND3X1_479 INVX1_460/Y INVX1_461/Y INVX1_462/Y gnd AOI21X1_315/B vdd NAND3X1
XDFFPOSX1_136 INVX1_28/A CLKBUF1_5/Y bloque_bytes[78] gnd vdd DFFPOSX1
XOAI21X1_497 BUFX2_223/A INVX1_404/A INVX1_405/A gnd INVX1_407/A vdd OAI21X1
XINVX1_318 INVX1_318/A gnd INVX1_318/Y vdd INVX1
XNAND2X1_611 AND2X2_159/B NOR2X1_384/A gnd NAND2X1_611/Y vdd NAND2X1
XXOR2X1_133 OR2X2_117/A gnd gnd OR2X2_113/B vdd XOR2X1
XNAND2X1_31 AOI21X1_17/A AOI21X1_17/B gnd INVX2_13/A vdd NAND2X1
XNAND3X1_443 INVX1_407/A OAI21X1_501/Y NAND2X1_541/Y gnd NAND3X1_443/Y vdd NAND3X1
XAOI21X1_270 OAI21X1_446/Y NAND2X1_487/Y INVX2_67/A gnd AOI21X1_271/B vdd AOI21X1
XOAI21X1_16 AND2X2_5/Y NOR2X1_22/Y INVX1_14/Y gnd NAND3X1_17/A vdd OAI21X1
XFILL_13_1_1 gnd vdd FILL
XDFFPOSX1_34 NOR2X1_410/A CLKBUF1_18/Y AND2X2_161/Y gnd vdd DFFPOSX1
XDFFPOSX1_100 NOR2X1_5/A CLKBUF1_48/Y XNOR2X1_243/Y gnd vdd DFFPOSX1
XXOR2X1_77 XOR2X1_77/A OR2X2_61/A gnd OR2X2_69/B vdd XOR2X1
XINVX1_282 INVX1_282/A gnd INVX1_282/Y vdd INVX1
XOAI21X1_461 NOR3X1_75/C OAI21X1_461/B INVX1_370/A gnd NOR2X1_293/A vdd OAI21X1
XOR2X2_160 OR2X2_160/A OR2X2_160/B gnd INVX1_595/A vdd OR2X2
XNAND2X1_575 INVX1_439/A NAND2X1_574/Y gnd INVX1_437/A vdd NAND2X1
XAOI21X1_234 INVX1_261/Y NAND3X1_343/C INVX1_260/A gnd AOI21X1_234/Y vdd AOI21X1
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XNAND3X1_407 INVX1_345/A OAI21X1_441/Y NAND3X1_402/Y gnd NAND3X1_407/Y vdd NAND3X1
XAND2X2_3 gnd OR2X2_2/B gnd AND2X2_3/Y vdd AND2X2
XAND2X2_177 AND2X2_177/A AND2X2_177/B gnd AND2X2_177/Y vdd AND2X2
XINVX1_246 INVX1_246/A gnd INVX1_246/Y vdd INVX1
XFILL_36_8_1 gnd vdd FILL
XOAI21X1_425 BUFX2_208/A XOR2X1_221/Y INVX1_330/Y gnd NAND3X1_391/B vdd OAI21X1
XXOR2X1_41 XOR2X1_39/B XOR2X1_41/B gnd XOR2X1_41/Y vdd XOR2X1
XNAND3X1_72 INVX1_48/A NAND3X1_72/B OR2X2_29/Y gnd OR2X2_32/B vdd NAND3X1
XOR2X2_124 BUFX2_171/A OR2X2_124/B gnd OR2X2_124/Y vdd OR2X2
XNAND2X1_539 INVX1_400/Y NOR2X1_315/Y gnd NAND3X1_439/B vdd NAND2X1
XAOI21X1_198 OR2X2_126/B OR2X2_126/A AND2X2_96/B gnd NOR2X1_175/A vdd AOI21X1
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XNAND3X1_371 INVX2_65/A NAND2X1_439/B NAND3X1_371/C gnd NOR3X1_69/A vdd NAND3X1
XNOR2X1_422 INVX2_86/Y INVX2_88/Y gnd NOR2X1_422/Y vdd NOR2X1
XINVX1_210 INVX1_210/A gnd INVX1_210/Y vdd INVX1
XOAI21X1_389 gnd XOR2X1_200/Y INVX1_284/Y gnd OAI21X1_389/Y vdd OAI21X1
XAND2X2_141 AND2X2_141/A AND2X2_141/B gnd XOR2X1_267/A vdd AND2X2
XNAND3X1_36 INVX1_26/A NAND3X1_34/B OR2X2_13/Y gnd OR2X2_16/B vdd NAND3X1
XFILL_12_4_0 gnd vdd FILL
XNAND2X1_503 INVX1_368/A NOR2X1_294/Y gnd NAND3X1_417/C vdd NAND2X1
XFILL_7_3 gnd vdd FILL
XFILL_10_6_1 gnd vdd FILL
XAOI21X1_162 OR2X2_102/B OR2X2_102/A AND2X2_78/B gnd NOR2X1_145/A vdd AOI21X1
XNAND3X1_335 INVX1_250/A NAND2X1_387/Y INVX1_249/Y gnd INVX1_256/A vdd NAND3X1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_174 INVX1_174/A gnd INVX1_174/Y vdd INVX1
XNOR2X1_386 NOR2X1_386/A NOR2X1_386/B gnd NOR2X1_386/Y vdd NOR2X1
XAND2X2_105 AND2X2_105/A AND2X2_105/B gnd XOR2X1_186/A vdd AND2X2
XOAI21X1_353 AOI21X1_232/Y INVX1_261/A INVX1_260/Y gnd AND2X2_113/A vdd OAI21X1
XNAND2X1_467 NAND3X1_391/Y AOI21X1_265/B gnd XOR2X1_233/B vdd NAND2X1
XFILL_2_0_0 gnd vdd FILL
XFILL_20_1_1 gnd vdd FILL
XFILL_0_2_1 gnd vdd FILL
XINVX1_20 OR2X2_8/Y gnd INVX1_20/Y vdd INVX1
XNAND3X1_299 AOI22X1_8/D AOI21X1_203/B INVX1_193/Y gnd AOI22X1_8/C vdd NAND3X1
XAND2X2_78 AND2X2_78/A AND2X2_78/B gnd AND2X2_78/Y vdd AND2X2
XAOI21X1_126 OR2X2_78/B OR2X2_78/A AND2X2_60/B gnd NOR2X1_115/A vdd AOI21X1
XOAI21X1_317 OAI21X1_317/A INVX1_221/A INVX1_224/A gnd NAND2X1_361/A vdd OAI21X1
XINVX1_138 INVX1_138/A gnd OR2X2_95/B vdd INVX1
XNAND2X1_431 XOR2X1_215/B NOR2X1_244/Y gnd NAND2X1_431/Y vdd NAND2X1
XNOR2X1_350 NOR2X1_350/A NOR2X1_349/Y gnd NOR2X1_350/Y vdd NOR2X1
XAND2X2_42 AND2X2_42/A AND2X2_42/B gnd AND2X2_42/Y vdd AND2X2
XNAND3X1_263 INVX1_167/Y NAND3X1_262/B OR2X2_115/Y gnd NAND3X1_263/Y vdd NAND3X1
XNOR3X1_4 NOR3X1_2/A MUX2X1_4/Y NOR3X1_2/C gnd NOR3X1_4/Y vdd NOR3X1
XBUFX2_264 OR2X2_69/A gnd BUFX2_264/Y vdd BUFX2
XINVX1_102 INVX1_102/A gnd INVX1_102/Y vdd INVX1
XOAI21X1_281 gnd NOR2X1_179/B INVX1_188/A gnd INVX2_59/A vdd OAI21X1
XBUFX4_27 INVX8_1/Y gnd BUFX4_27/Y vdd BUFX4
XNOR2X1_314 NOR2X1_314/A NOR2X1_314/B gnd BUFX2_233/A vdd NOR2X1
XNAND2X1_395 XNOR2X1_163/B NAND2X1_395/B gnd NOR2X1_224/B vdd NAND2X1
XNAND3X1_227 INVX1_145/Y NAND3X1_227/B OR2X2_99/Y gnd AOI21X1_157/B vdd NAND3X1
XBUFX2_228 BUFX2_228/A gnd BUFX2_228/Y vdd BUFX2
XNOR2X1_81 NOR2X1_81/A INVX2_30/A gnd NOR2X1_81/Y vdd NOR2X1
XFILL_17_6_1 gnd vdd FILL
XFILL_19_4_0 gnd vdd FILL
XOAI21X1_245 NOR2X1_157/A INVX1_163/Y INVX1_164/Y gnd NAND2X1_285/B vdd OAI21X1
XNAND2X1_359 NAND2X1_359/A INVX1_221/Y gnd INVX1_222/A vdd NAND2X1
XINVX2_66 INVX2_66/A gnd INVX2_66/Y vdd INVX2
XNOR2X1_278 NOR2X1_278/A NOR2X1_278/B gnd BUFX2_221/A vdd NOR2X1
XFILL_11_1 gnd vdd FILL
XXNOR2X1_230 AOI21X1_354/C bloque_bytes[20] gnd AND2X2_184/B vdd XNOR2X1
XBUFX2_192 BUFX2_192/A gnd BUFX2_192/Y vdd BUFX2
XNAND3X1_191 INVX1_123/Y NAND2X1_216/Y OR2X2_83/Y gnd AOI21X1_133/B vdd NAND3X1
XNOR2X1_45 NOR2X1_45/A INVX1_38/Y gnd NOR2X1_45/Y vdd NOR2X1
XFILL_7_2_1 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XOAI21X1_209 INVX2_46/Y AND2X2_72/B OR2X2_94/Y gnd OAI21X1_210/B vdd OAI21X1
XFILL_27_1_1 gnd vdd FILL
XINVX2_30 INVX2_30/A gnd INVX2_30/Y vdd INVX2
XNAND2X1_323 NAND2X1_323/A NAND2X1_323/B gnd XOR2X1_169/A vdd NAND2X1
XNOR2X1_242 NOR2X1_242/A NOR2X1_242/B gnd BUFX2_209/A vdd NOR2X1
XNAND3X1_155 INVX1_101/Y AOI21X1_110/A OR2X2_67/Y gnd AOI21X1_109/B vdd NAND3X1
XCLKBUF1_33 BUFX4_1/Y gnd CLKBUF1_33/Y vdd CLKBUF1
XINVX1_571 INVX1_571/A gnd INVX1_571/Y vdd INVX1
XBUFX2_156 OR2X2_93/A gnd BUFX2_156/Y vdd BUFX2
XXNOR2X1_194 NOR2X1_321/Y XNOR2X1_194/B gnd XNOR2X1_195/A vdd XNOR2X1
XNOR2X1_206 NOR2X1_206/A NOR2X1_206/B gnd BUFX2_193/A vdd NOR2X1
XOAI21X1_173 AND2X2_61/Y NOR2X1_114/Y INVX1_114/Y gnd OAI21X1_173/Y vdd OAI21X1
XFILL_33_1 gnd vdd FILL
XNAND2X1_287 gnd OR2X2_113/B gnd NAND3X1_257/B vdd NAND2X1
XFILL_16_9_0 gnd vdd FILL
XNOR3X1_86 NOR3X1_86/A INVX2_73/Y NOR3X1_86/C gnd NOR3X1_86/Y vdd NOR3X1
XNAND3X1_119 INVX1_79/Y AOI21X1_86/A OR2X2_51/Y gnd AOI21X1_85/B vdd NAND3X1
XINVX1_535 bloque_bytes[79] gnd INVX1_535/Y vdd INVX1
XBUFX2_120 gnd gnd BUFX2_120/Y vdd BUFX2
XDFFPOSX1_353 XNOR2X1_198/B CLKBUF1_46/Y OAI21X1_629/Y gnd vdd DFFPOSX1
XXNOR2X1_80 XNOR2X1_80/A AND2X2_54/Y gnd XOR2X1_96/A vdd XNOR2X1
XXNOR2X1_158 NOR2X1_213/Y XNOR2X1_158/B gnd XNOR2X1_159/A vdd XNOR2X1
XOAI21X1_137 XNOR2X1_71/A AOI21X1_101/C AND2X2_48/B gnd XNOR2X1_72/A vdd OAI21X1
XBUFX4_2 clk gnd BUFX4_2/Y vdd BUFX4
XNAND2X1_251 gnd OR2X2_98/B gnd AOI21X1_155/A vdd NAND2X1
XNOR2X1_170 gnd OR2X2_123/B gnd NOR2X1_170/Y vdd NOR2X1
XFILL_26_4_0 gnd vdd FILL
XFILL_6_5_0 gnd vdd FILL
XNOR3X1_50 INVX1_144/Y NOR3X1_50/B NOR3X1_50/C gnd NOR3X1_50/Y vdd NOR3X1
XFILL_24_6_1 gnd vdd FILL
XDFFPOSX1_317 INVX1_343/A CLKBUF1_39/Y INVX1_563/Y gnd vdd DFFPOSX1
XFILL_4_7_1 gnd vdd FILL
XXOR2X1_314 vdd gnd gnd OR2X2_5/B vdd XOR2X1
XINVX1_499 bloque_bytes[30] gnd INVX1_499/Y vdd INVX1
XXNOR2X1_122 XNOR2X1_122/A INVX2_50/Y gnd BUFX2_171/A vdd XNOR2X1
XXNOR2X1_44 OAI21X1_89/A AND2X2_30/Y gnd XOR2X1_56/A vdd XNOR2X1
XOAI21X1_101 AND2X2_35/Y NOR2X1_72/Y INVX1_69/Y gnd NAND3X1_107/A vdd OAI21X1
XNOR2X1_134 OR2X2_93/A OR2X2_93/B gnd NOR2X1_134/Y vdd NOR2X1
XNAND2X1_215 INVX1_129/A NAND2X1_215/B gnd OAI21X1_182/A vdd NAND2X1
XFILL_34_1_1 gnd vdd FILL
XNOR3X1_14 BUFX4_25/Y MUX2X1_14/Y BUFX4_21/Y gnd NOR3X1_14/Y vdd NOR3X1
XOAI21X1_642 AND2X2_196/Y NOR2X1_449/Y INVX1_593/A gnd NAND3X1_540/C vdd OAI21X1
XDFFPOSX1_281 XNOR2X1_162/B CLKBUF1_31/Y NOR2X1_434/B gnd vdd DFFPOSX1
XINVX1_463 INVX1_463/A gnd INVX1_463/Y vdd INVX1
XXOR2X1_278 XOR2X1_278/A XOR2X1_278/B gnd XOR2X1_278/Y vdd XOR2X1
XNAND2X1_179 OR2X2_68/A OR2X2_68/B gnd NAND2X1_179/Y vdd NAND2X1
XDFFPOSX1_245 INVX1_178/A CLKBUF1_21/Y OR2X2_152/B gnd vdd DFFPOSX1
XMUX2X1_24 BUFX2_24/A INVX1_5/A MUX2X1_8/S gnd MUX2X1_24/Y vdd MUX2X1
XOR2X2_66 gnd OR2X2_66/B gnd OR2X2_66/Y vdd OR2X2
XAOI21X1_77 AOI21X1_77/A AOI21X1_77/B AOI21X1_77/C gnd AOI21X1_77/Y vdd AOI21X1
XOAI21X1_606 INVX1_521/Y bloque_bytes[21] INVX1_522/Y gnd AOI21X1_367/C vdd OAI21X1
XINVX1_427 INVX1_427/A gnd INVX1_427/Y vdd INVX1
XNAND2X1_720 NAND2X1_720/A INVX1_599/A gnd INVX1_597/A vdd NAND2X1
XFILL_23_9_0 gnd vdd FILL
XBUFX2_80 gnd gnd BUFX2_80/Y vdd BUFX2
XXOR2X1_242 XOR2X1_242/A XOR2X1_242/B gnd XOR2X1_242/Y vdd XOR2X1
XNAND2X1_143 AND2X2_42/B AND2X2_42/A gnd AOI21X1_89/C vdd NAND2X1
XAOI21X1_379 AOI21X1_379/A AOI21X1_379/B AOI21X1_379/C gnd INVX1_558/A vdd AOI21X1
XOR2X2_30 OR2X2_30/A OR2X2_30/B gnd INVX1_49/A vdd OR2X2
XAOI21X1_41 AOI21X1_41/A AOI21X1_41/B OAI21X1_52/B gnd NAND3X1_56/B vdd AOI21X1
XDFFPOSX1_209 XOR2X1_111/B CLKBUF1_49/Y bloque_bytes[7] gnd vdd DFFPOSX1
XOAI21X1_570 INVX4_2/Y INVX1_474/A BUFX4_33/Y gnd OAI21X1_570/Y vdd OAI21X1
XFILL_20_3 gnd vdd FILL
XXOR2X1_206 XOR2X1_206/A XOR2X1_206/B gnd XOR2X1_206/Y vdd XOR2X1
XFILL_33_4_0 gnd vdd FILL
XINVX1_391 INVX1_391/A gnd INVX1_391/Y vdd INVX1
XFILL_31_6_1 gnd vdd FILL
XNAND2X1_684 INVX1_560/A XNOR2X1_236/Y gnd NAND2X1_684/Y vdd NAND2X1
XBUFX2_44 gnd gnd BUFX2_44/Y vdd BUFX2
XOAI21X1_89 OAI21X1_89/A OAI21X1_89/B NOR2X1_65/Y gnd NOR2X1_66/B vdd OAI21X1
XNAND2X1_107 NAND3X1_89/Y AOI21X1_65/B gnd INVX2_25/A vdd NAND2X1
XAOI21X1_343 NOR2X1_404/Y NOR3X1_90/Y BUFX4_15/Y gnd AND2X2_175/B vdd AOI21X1
XNAND3X1_516 INVX1_516/Y INVX1_571/Y INVX1_550/A gnd NAND3X1_516/Y vdd NAND3X1
XDFFPOSX1_173 INVX1_79/A CLKBUF1_1/Y bloque_bytes[35] gnd vdd DFFPOSX1
XOAI21X1_534 gnd NOR2X1_339/B INVX1_438/A gnd INVX1_440/A vdd OAI21X1
XINVX1_355 INVX1_355/A gnd INVX1_355/Y vdd INVX1
XXOR2X1_170 XOR2X1_170/A XOR2X1_170/B gnd XOR2X1_176/A vdd XOR2X1
XNAND2X1_648 NAND2X1_647/Y OR2X2_134/Y gnd NAND2X1_648/Y vdd NAND2X1
XAOI21X1_307 INVX1_445/A NAND3X1_466/Y INVX1_440/Y gnd NOR2X1_340/B vdd AOI21X1
XDFFPOSX1_137 XOR2X1_21/B CLKBUF1_16/Y bloque_bytes[79] gnd vdd DFFPOSX1
XNAND2X1_68 OR2X2_21/A OR2X2_21/B gnd NAND3X1_52/B vdd NAND2X1
XOAI21X1_53 AND2X2_19/Y NOR2X1_44/Y INVX1_37/A gnd NAND3X1_53/B vdd OAI21X1
XDFFPOSX1_71 AND2X2_164/B CLKBUF1_15/Y NOR2X1_396/Y gnd vdd DFFPOSX1
XNAND3X1_480 INVX1_462/A INVX1_460/Y INVX1_461/Y gnd NAND3X1_480/Y vdd NAND3X1
XXOR2X1_134 BUFX2_169/A gnd gnd OR2X2_114/B vdd XOR2X1
XOAI21X1_498 BUFX2_223/A INVX1_404/A INVX1_405/Y gnd NAND3X1_446/B vdd OAI21X1
XINVX1_319 INVX1_319/A gnd INVX1_319/Y vdd INVX1
XNAND2X1_612 INVX8_2/A NAND2X1_612/B gnd NOR2X1_385/B vdd NAND2X1
XOAI21X1_17 OAI21X1_17/A XNOR2X1_7/B OAI21X1_17/C gnd NAND2X1_28/B vdd OAI21X1
XNAND2X1_32 NAND3X1_19/A OR2X2_8/B gnd OR2X2_6/A vdd NAND2X1
XNAND3X1_444 AOI22X1_19/B INVX1_409/A INVX1_407/Y gnd NAND3X1_444/Y vdd NAND3X1
XAOI21X1_271 NAND3X1_399/Y AOI21X1_271/B INVX1_351/Y gnd AOI21X1_272/A vdd AOI21X1
XFILL_30_9_0 gnd vdd FILL
XDFFPOSX1_35 NOR2X1_411/A CLKBUF1_18/Y NOR2X1_363/Y gnd vdd DFFPOSX1
XINVX1_283 INVX1_283/A gnd INVX1_283/Y vdd INVX1
XOAI21X1_462 NOR2X1_293/Y NOR2X1_292/B AOI22X1_17/C gnd XOR2X1_251/A vdd OAI21X1
XDFFPOSX1_101 NOR2X1_4/A CLKBUF1_42/Y XNOR2X1_244/Y gnd vdd DFFPOSX1
XXOR2X1_78 NOR2X1_87/Y XOR2X1_78/B gnd XOR2X1_78/Y vdd XOR2X1
XNAND2X1_576 INVX1_438/A NOR2X1_339/Y gnd NAND2X1_576/Y vdd NAND2X1
XOR2X2_161 OR2X2_161/A OR2X2_161/B gnd OR2X2_161/Y vdd OR2X2
XAOI22X1_10 INVX1_238/A AOI22X1_10/B AOI22X1_10/C INVX1_236/A gnd INVX1_242/A vdd
+ AOI22X1
XAOI21X1_235 INVX1_274/A AOI21X1_235/B INVX1_269/Y gnd NOR2X1_232/B vdd AOI21X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XNAND3X1_408 INVX1_356/Y INVX1_355/A OAI21X1_449/Y gnd AND2X2_133/B vdd NAND3X1
XAND2X2_4 gnd OR2X2_3/B gnd AND2X2_4/Y vdd AND2X2
XAND2X2_178 bloque_bytes[32] OR2X2_142/B gnd AND2X2_178/Y vdd AND2X2
XINVX1_247 INVX1_247/A gnd INVX1_247/Y vdd INVX1
XOAI21X1_426 BUFX2_208/A XOR2X1_221/Y INVX1_330/A gnd AOI22X1_15/B vdd OAI21X1
XNAND3X1_73 NAND3X1_73/A OR2X2_32/B OR2X2_30/B gnd AOI21X1_53/B vdd NAND3X1
XXOR2X1_42 OR2X2_44/A gnd gnd XOR2X1_42/Y vdd XOR2X1
XOR2X2_125 OR2X2_125/A OR2X2_125/B gnd OR2X2_125/Y vdd OR2X2
XNAND2X1_540 NAND3X1_445/B INVX1_408/A gnd XNOR2X1_192/B vdd NAND2X1
XAOI21X1_199 NOR2X1_175/Y AOI21X1_199/B INVX1_183/A gnd NOR2X1_177/A vdd AOI21X1
XNAND3X1_372 INVX1_306/A NAND2X1_442/B INVX2_65/Y gnd OAI21X1_404/B vdd NAND3X1
XINVX1_93 OR2X2_62/Y gnd INVX1_93/Y vdd INVX1
XNAND3X1_37 NAND3X1_37/A OR2X2_16/B OR2X2_14/B gnd AOI21X1_29/B vdd NAND3X1
XFILL_14_2_0 gnd vdd FILL
XNOR2X1_423 bloque_bytes[37] INVX2_88/A gnd NOR2X1_423/Y vdd NOR2X1
XINVX1_211 INVX1_211/A gnd INVX1_211/Y vdd INVX1
XOAI21X1_390 BUFX2_201/A XOR2X1_204/Y INVX1_296/A gnd OAI21X1_390/Y vdd OAI21X1
XAND2X2_142 NOR2X1_310/Y INVX1_396/Y gnd NOR3X1_80/A vdd AND2X2
XFILL_12_4_1 gnd vdd FILL
XNAND2X1_504 INVX1_368/Y NOR2X1_294/Y gnd INVX1_371/A vdd NAND2X1
XAOI21X1_163 NOR2X1_145/Y AOI21X1_163/B INVX1_150/A gnd NOR2X1_147/A vdd AOI21X1
XNAND3X1_336 INVX1_251/Y INVX1_252/Y INVX1_253/Y gnd NAND3X1_336/Y vdd NAND3X1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XINVX1_175 INVX1_175/A gnd INVX1_175/Y vdd INVX1
XOAI21X1_354 NOR2X1_221/A NOR3X1_63/Y AOI21X1_233/Y gnd NAND3X1_343/C vdd OAI21X1
XNOR2X1_387 OR2X2_129/A OR2X2_129/B gnd NOR2X1_387/Y vdd NOR2X1
XAND2X2_106 NOR2X1_202/Y INVX1_225/Y gnd NOR3X1_62/A vdd AND2X2
XNAND2X1_468 INVX1_322/A NOR2X1_264/Y gnd NAND2X1_468/Y vdd NAND2X1
XFILL_2_0_1 gnd vdd FILL
XAND2X2_79 OR2X2_101/A OR2X2_101/B gnd AND2X2_79/Y vdd AND2X2
XAOI21X1_127 NOR2X1_115/Y AOI21X1_127/B INVX1_117/A gnd NOR2X1_117/A vdd AOI21X1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XNAND3X1_300 AOI22X1_8/D NAND3X1_300/B NAND3X1_300/C gnd NAND2X1_334/A vdd NAND3X1
XOAI21X1_318 gnd NOR2X1_202/B INVX1_225/A gnd NAND2X1_363/A vdd OAI21X1
XINVX1_139 INVX1_139/A gnd INVX1_139/Y vdd INVX1
XNOR2X1_351 gnd XOR2X1_282/Y gnd NOR2X1_351/Y vdd NOR2X1
XNAND2X1_432 INVX1_296/Y NOR2X1_247/Y gnd NAND2X1_433/B vdd NAND2X1
XAND2X2_43 OR2X2_53/A OR2X2_53/B gnd AND2X2_43/Y vdd AND2X2
XBUFX2_265 XOR2X1_74/A gnd BUFX2_265/Y vdd BUFX2
XNAND3X1_264 INVX1_168/Y NAND3X1_264/B OR2X2_116/Y gnd NAND3X1_265/B vdd NAND3X1
XNOR3X1_5 NOR3X1_3/A MUX2X1_5/Y NOR3X1_3/C gnd NOR3X1_5/Y vdd NOR3X1
XINVX1_103 INVX1_103/A gnd INVX1_103/Y vdd INVX1
XFILL_11_7_0 gnd vdd FILL
XOAI21X1_282 NOR3X1_58/C INVX2_59/Y NOR3X1_58/A gnd AND2X2_100/A vdd OAI21X1
XBUFX4_28 reset gnd INVX8_2/A vdd BUFX4
XNAND2X1_396 INVX1_257/Y NOR2X1_224/B gnd NAND2X1_397/A vdd NAND2X1
XAOI22X1_1 INVX2_1/Y target[5] target[4] INVX2_2/Y gnd NAND2X1_2/A vdd AOI22X1
XNOR2X1_315 gnd XOR2X1_255/Y gnd NOR2X1_315/Y vdd NOR2X1
XNAND3X1_228 INVX1_146/Y NAND3X1_228/B OR2X2_100/Y gnd NAND3X1_229/B vdd NAND3X1
XFILL_19_4_1 gnd vdd FILL
XFILL_21_2_0 gnd vdd FILL
XBUFX2_229 BUFX2_229/A gnd BUFX2_229/Y vdd BUFX2
XFILL_1_3_0 gnd vdd FILL
XNOR2X1_82 OR2X2_52/A OR2X2_52/B gnd NOR2X1_82/Y vdd NOR2X1
XOAI21X1_246 NOR3X1_53/C NOR3X1_53/B INVX1_165/Y gnd OAI21X1_246/Y vdd OAI21X1
XFILL_11_2 gnd vdd FILL
XNAND2X1_360 NAND2X1_360/A AOI22X1_9/C gnd NAND2X1_360/Y vdd NAND2X1
XINVX2_67 INVX2_67/A gnd INVX2_67/Y vdd INVX2
XNOR2X1_279 gnd NOR2X1_279/B gnd NOR2X1_279/Y vdd NOR2X1
XNOR2X1_46 INVX1_40/Y NOR2X1_46/B gnd NOR2X1_46/Y vdd NOR2X1
XXNOR2X1_231 INVX1_574/A bloque_bytes[21] gnd AND2X2_185/B vdd XNOR2X1
XNAND3X1_192 INVX1_124/Y AOI21X1_136/A OR2X2_84/Y gnd NAND3X1_193/B vdd NAND3X1
XBUFX2_193 BUFX2_193/A gnd BUFX2_193/Y vdd BUFX2
XINVX2_31 INVX2_31/A gnd INVX2_31/Y vdd INVX2
XFILL_9_0_1 gnd vdd FILL
XOAI21X1_210 OAI21X1_210/A OAI21X1_210/B INVX1_139/Y gnd OAI21X1_210/Y vdd OAI21X1
XNOR2X1_243 gnd XOR2X1_201/Y gnd NOR2X1_243/Y vdd NOR2X1
XNAND2X1_324 AND2X2_98/B AND2X2_98/A gnd NAND3X1_293/B vdd NAND2X1
XNAND3X1_156 INVX1_102/Y NAND2X1_179/Y OR2X2_68/Y gnd NAND3X1_157/B vdd NAND3X1
XBUFX2_157 BUFX2_157/A gnd BUFX2_157/Y vdd BUFX2
XINVX1_572 INVX1_572/A gnd INVX1_572/Y vdd INVX1
XCLKBUF1_34 BUFX4_5/Y gnd CLKBUF1_34/Y vdd CLKBUF1
XOAI21X1_174 XNOR2X1_89/A OAI21X1_174/B NOR2X1_115/Y gnd NOR2X1_116/B vdd OAI21X1
XNOR2X1_10 NOR2X1_10/A NOR2X1_10/B gnd AOI21X1_5/C vdd NOR2X1
XXNOR2X1_1 target[6] XOR2X1_1/B gnd XNOR2X1_1/Y vdd XNOR2X1
XXNOR2X1_195 XNOR2X1_195/A OAI21X1_504/Y gnd INVX1_414/A vdd XNOR2X1
XNAND2X1_288 OAI21X1_246/Y NAND3X1_260/B gnd NAND2X1_288/Y vdd NAND2X1
XNOR2X1_207 gnd NOR2X1_207/B gnd NOR2X1_207/Y vdd NOR2X1
XFILL_18_7_0 gnd vdd FILL
XFILL_33_2 gnd vdd FILL
XNOR3X1_87 BUFX4_14/Y NOR3X1_87/B NOR3X1_87/C gnd NOR3X1_87/Y vdd NOR3X1
XFILL_16_9_1 gnd vdd FILL
XDFFPOSX1_354 INVX1_434/A CLKBUF1_13/Y OR2X2_150/Y gnd vdd DFFPOSX1
XNAND3X1_120 INVX1_80/Y AOI21X1_88/A OR2X2_52/Y gnd NAND3X1_120/Y vdd NAND3X1
XBUFX4_3 clk gnd BUFX4_3/Y vdd BUFX4
XINVX1_536 bloque_bytes[66] gnd INVX1_536/Y vdd INVX1
XBUFX2_121 gnd gnd BUFX2_121/Y vdd BUFX2
XXNOR2X1_81 XNOR2X1_81/A INVX2_37/Y gnd XOR2X1_97/A vdd XNOR2X1
XXNOR2X1_159 XNOR2X1_159/A NAND2X1_376/A gnd INVX1_243/A vdd XNOR2X1
XOAI21X1_138 AND2X2_49/Y NOR2X1_94/Y INVX1_92/A gnd OAI21X1_138/Y vdd OAI21X1
XFILL_28_2_0 gnd vdd FILL
XFILL_8_3_0 gnd vdd FILL
XNAND2X1_252 NAND2X1_252/A NAND2X1_252/B gnd XNOR2X1_115/A vdd NAND2X1
XNOR2X1_171 NOR2X1_171/A INVX2_57/A gnd XOR2X1_160/B vdd NOR2X1
XFILL_26_4_1 gnd vdd FILL
XFILL_6_5_1 gnd vdd FILL
XINVX1_500 bloque_bytes[31] gnd INVX1_500/Y vdd INVX1
XNOR3X1_51 INVX1_154/Y NOR3X1_51/B NOR3X1_51/C gnd NOR3X1_51/Y vdd NOR3X1
XDFFPOSX1_318 INVX1_348/A CLKBUF1_39/Y INVX1_565/Y gnd vdd DFFPOSX1
XXOR2X1_315 vdd gnd gnd XOR2X1_315/Y vdd XOR2X1
XXNOR2X1_123 XNOR2X1_123/A XNOR2X1_123/B gnd OR2X2_125/A vdd XNOR2X1
XXNOR2X1_45 OAI21X1_86/Y INVX2_25/Y gnd XOR2X1_57/A vdd XNOR2X1
XOAI21X1_102 OAI21X1_97/A XNOR2X1_52/B AOI21X1_75/Y gnd NAND3X1_110/C vdd OAI21X1
XNOR2X1_135 NOR2X1_135/A INVX1_137/Y gnd NOR2X1_135/Y vdd NOR2X1
XNAND2X1_216 gnd OR2X2_83/B gnd NAND2X1_216/Y vdd NAND2X1
XNOR3X1_15 BUFX4_27/Y MUX2X1_15/Y BUFX4_20/Y gnd NOR3X1_15/Y vdd NOR3X1
XOAI21X1_643 AND2X2_196/Y NOR2X1_449/Y INVX1_593/Y gnd NAND3X1_544/A vdd OAI21X1
XDFFPOSX1_282 INVX1_263/A CLKBUF1_19/Y OR2X2_135/A gnd vdd DFFPOSX1
XINVX1_464 INVX1_464/A gnd INVX1_464/Y vdd INVX1
XXOR2X1_279 INVX1_460/A gnd gnd XOR2X1_279/Y vdd XOR2X1
XNAND2X1_180 INVX2_36/Y NAND3X1_164/C gnd XNOR2X1_80/A vdd NAND2X1
XAOI21X1_78 OR2X2_46/B OR2X2_46/A AND2X2_36/B gnd NOR2X1_75/A vdd AOI21X1
XDFFPOSX1_246 INVX1_179/A CLKBUF1_51/Y OR2X2_153/B gnd vdd DFFPOSX1
XOR2X2_67 gnd OR2X2_67/B gnd OR2X2_67/Y vdd OR2X2
XOAI21X1_607 INVX1_524/Y bloque_bytes[22] INVX1_525/Y gnd AOI21X1_368/C vdd OAI21X1
XFILL_23_9_1 gnd vdd FILL
XFILL_25_7_0 gnd vdd FILL
XINVX1_428 INVX1_428/A gnd INVX1_428/Y vdd INVX1
XXOR2X1_243 BUFX2_219/A gnd gnd XOR2X1_243/Y vdd XOR2X1
XNAND2X1_721 INVX2_94/A AND2X2_197/Y gnd OAI21X1_648/B vdd NAND2X1
XFILL_5_8_0 gnd vdd FILL
XBUFX2_81 gnd gnd BUFX2_81/Y vdd BUFX2
XNAND2X1_144 OR2X2_53/A OR2X2_53/B gnd NAND3X1_126/B vdd NAND2X1
XAOI21X1_380 NAND2X1_664/Y AOI21X1_380/B NAND3X1_504/Y gnd INVX1_560/A vdd AOI21X1
XOR2X2_31 OR2X2_31/A OR2X2_31/B gnd OR2X2_31/Y vdd OR2X2
XAOI21X1_42 OR2X2_22/B OR2X2_22/A AND2X2_18/B gnd NOR2X1_45/A vdd AOI21X1
XOAI21X1_571 INVX4_2/A NOR2X1_388/B BUFX4_33/Y gnd NOR2X1_386/A vdd OAI21X1
XDFFPOSX1_210 INVX2_44/A CLKBUF1_36/Y OR2X2_142/B gnd vdd DFFPOSX1
XFILL_35_2_0 gnd vdd FILL
XINVX1_392 INVX1_392/A gnd INVX1_392/Y vdd INVX1
XNAND2X1_685 INVX1_537/Y INVX1_561/A gnd NAND2X1_685/Y vdd NAND2X1
XFILL_33_4_1 gnd vdd FILL
XXOR2X1_207 BUFX2_203/A gnd gnd XOR2X1_207/Y vdd XOR2X1
XNAND2X1_108 NAND3X1_91/A OR2X2_40/B gnd OR2X2_38/A vdd NAND2X1
XBUFX2_45 gnd gnd BUFX2_45/Y vdd BUFX2
XAOI21X1_344 NOR2X1_404/Y NOR3X1_90/Y AND2X2_167/B gnd NOR2X1_405/A vdd AOI21X1
XDFFPOSX1_174 INVX1_80/A CLKBUF1_1/Y bloque_bytes[36] gnd vdd DFFPOSX1
XOAI21X1_90 INVX2_25/Y AND2X2_30/B OR2X2_38/Y gnd OAI21X1_90/Y vdd OAI21X1
XNAND3X1_517 INVX1_519/Y INVX1_572/Y INVX1_551/A gnd NAND3X1_517/Y vdd NAND3X1
XINVX1_356 INVX1_356/A gnd INVX1_356/Y vdd INVX1
XOAI21X1_535 BUFX2_231/A INVX1_442/A INVX1_443/A gnd INVX1_445/A vdd OAI21X1
XXOR2X1_171 BUFX2_183/A gnd gnd NOR2X1_202/B vdd XOR2X1
XNAND2X1_649 INVX1_504/Y NAND2X1_648/Y gnd OR2X2_153/B vdd NAND2X1
XNAND2X1_69 AOI21X1_41/A AOI21X1_41/B gnd INVX2_19/A vdd NAND2X1
XNAND3X1_481 INVX1_464/A AOI21X1_315/B INVX1_459/Y gnd AOI22X1_22/C vdd NAND3X1
XAOI21X1_308 OAI21X1_536/Y NAND3X1_467/Y INVX1_440/A gnd NOR2X1_340/A vdd AOI21X1
XOAI21X1_54 AND2X2_19/Y NOR2X1_44/Y INVX1_37/Y gnd NAND3X1_55/A vdd OAI21X1
XDFFPOSX1_138 INVX2_17/A CLKBUF1_33/Y bloque_bytes[64] gnd vdd DFFPOSX1
XDFFPOSX1_72 INVX1_478/A CLKBUF1_15/Y NOR3X1_88/Y gnd vdd DFFPOSX1
XXOR2X1_135 BUFX2_170/A gnd gnd OR2X2_115/B vdd XOR2X1
XINVX1_320 INVX1_320/A gnd INVX1_320/Y vdd INVX1
XOAI21X1_499 NOR3X1_79/C NAND3X1_437/Y INVX1_408/A gnd NOR2X1_317/A vdd OAI21X1
XNAND2X1_613 INVX1_474/A AND2X2_169/B gnd NOR2X1_388/B vdd NAND2X1
XFILL_32_7_0 gnd vdd FILL
XNAND2X1_33 OR2X2_7/B OR2X2_7/A gnd NAND2X1_34/A vdd NAND2X1
XOAI21X1_18 XNOR2X1_8/A OAI21X1_18/B AND2X2_6/B gnd XNOR2X1_9/A vdd OAI21X1
XDFFPOSX1_36 INVX1_537/A CLKBUF1_18/Y AND2X2_162/Y gnd vdd DFFPOSX1
XNAND3X1_445 INVX1_399/Y NAND3X1_445/B NOR3X1_80/Y gnd AOI21X1_296/B vdd NAND3X1
XAOI21X1_272 AOI21X1_272/A AOI21X1_272/B AOI21X1_272/C gnd OAI21X1_448/A vdd AOI21X1
XFILL_30_9_1 gnd vdd FILL
XINVX1_284 INVX1_284/A gnd INVX1_284/Y vdd INVX1
XOAI21X1_463 BUFX2_216/A NOR2X1_294/B INVX1_368/Y gnd OAI21X1_463/Y vdd OAI21X1
XDFFPOSX1_102 INVX2_2/A CLKBUF1_42/Y XOR2X1_305/Y gnd vdd DFFPOSX1
XOR2X2_162 OR2X2_162/A OR2X2_162/B gnd INVX1_599/A vdd OR2X2
XXOR2X1_79 XOR2X1_79/A BUFX2_262/A gnd XOR2X1_79/Y vdd XOR2X1
XNAND2X1_577 INVX1_438/Y NOR2X1_339/Y gnd AOI21X1_309/B vdd NAND2X1
XAOI22X1_11 INVX1_257/A AOI22X1_11/B AOI22X1_11/C INVX1_255/A gnd INVX1_261/A vdd
+ AOI22X1
XAOI21X1_236 AOI21X1_236/A AOI21X1_236/B INVX1_269/A gnd NOR2X1_232/A vdd AOI21X1
XNAND3X1_409 INVX1_354/Y INVX1_357/Y AND2X2_133/A gnd NAND3X1_409/Y vdd NAND3X1
XAND2X2_5 gnd OR2X2_4/B gnd AND2X2_5/Y vdd AND2X2
XXOR2X1_43 OR2X2_45/A gnd gnd OR2X2_41/B vdd XOR2X1
XAND2X2_179 bloque_bytes[33] OR2X2_143/B gnd AND2X2_179/Y vdd AND2X2
XINVX1_248 INVX1_248/A gnd INVX1_248/Y vdd INVX1
XOAI21X1_427 gnd NOR2X1_264/B INVX1_322/Y gnd OAI21X1_427/Y vdd OAI21X1
XNAND3X1_74 INVX2_21/Y AOI21X1_53/Y NAND3X1_74/C gnd AOI21X1_55/B vdd NAND3X1
XOR2X2_126 OR2X2_126/A OR2X2_126/B gnd INVX1_181/A vdd OR2X2
XNAND2X1_541 INVX1_406/A NOR2X1_318/Y gnd NAND2X1_541/Y vdd NAND2X1
XAOI21X1_200 INVX2_57/Y INVX1_184/Y NOR2X1_171/A gnd AOI21X1_202/A vdd AOI21X1
XFILL_24_1 gnd vdd FILL
XNAND3X1_373 INVX1_306/A OAI21X1_400/Y NAND3X1_373/C gnd AOI21X1_255/A vdd NAND3X1
XINVX1_94 INVX1_94/A gnd OR2X2_63/B vdd INVX1
XINVX1_212 INVX1_212/A gnd INVX1_212/Y vdd INVX1
XNAND3X1_38 INVX2_15/Y NAND3X1_38/B OAI21X1_34/Y gnd NAND3X1_38/Y vdd NAND3X1
XNOR2X1_424 INVX2_87/Y INVX2_89/Y gnd NOR2X1_424/Y vdd NOR2X1
XFILL_14_2_1 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XOAI21X1_391 OAI21X1_391/A INVX1_299/A INVX1_298/Y gnd AND2X2_121/A vdd OAI21X1
XNAND2X1_505 NAND3X1_417/Y AOI21X1_281/B gnd XOR2X1_251/B vdd NAND2X1
XAND2X2_143 NOR2X1_311/Y INVX1_397/Y gnd NOR3X1_80/C vdd AND2X2
XAOI21X1_164 INVX2_48/Y INVX1_151/Y NOR2X1_141/A gnd AOI21X1_166/A vdd AOI21X1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XNAND3X1_337 INVX1_253/A INVX1_251/Y INVX1_252/Y gnd AOI21X1_228/B vdd NAND3X1
XAND2X2_107 AND2X2_107/A INVX1_226/Y gnd NOR3X1_62/C vdd AND2X2
XOAI21X1_355 AOI21X1_234/Y INVX1_259/A INVX1_262/A gnd OAI21X1_355/Y vdd OAI21X1
XINVX1_176 INVX1_176/A gnd NOR3X1_55/A vdd INVX1
XNOR2X1_388 NOR2X1_388/A NOR2X1_388/B gnd NOR2X1_388/Y vdd NOR2X1
XNAND2X1_469 XOR2X1_233/B NOR2X1_268/Y gnd NAND2X1_469/Y vdd NAND2X1
XNAND3X1_301 AOI22X1_8/B INVX1_200/A INVX1_198/Y gnd NAND2X1_334/B vdd NAND3X1
XAND2X2_80 gnd OR2X2_105/B gnd NOR3X1_51/C vdd AND2X2
XAOI21X1_128 INVX2_39/Y INVX1_118/Y NOR2X1_111/A gnd AOI21X1_130/A vdd AOI21X1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XOAI21X1_319 gnd NOR2X1_203/B INVX1_226/A gnd INVX2_61/A vdd OAI21X1
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XNOR2X1_352 NOR2X1_352/A NOR2X1_352/B gnd NOR2X1_352/Y vdd NOR2X1
XNAND2X1_433 OAI21X1_390/Y NAND2X1_433/B gnd NOR2X1_248/B vdd NAND2X1
XNAND3X1_265 AOI21X1_180/A NAND3X1_265/B NAND3X1_265/C gnd AND2X2_90/B vdd NAND3X1
XFILL_11_7_1 gnd vdd FILL
XFILL_13_5_0 gnd vdd FILL
XBUFX2_266 XOR2X1_75/A gnd BUFX2_266/Y vdd BUFX2
XAND2X2_44 gnd OR2X2_57/B gnd NOR3X1_39/C vdd AND2X2
XNOR3X1_6 NOR3X1_2/A NOR3X1_6/B NOR3X1_2/C gnd NOR3X1_6/Y vdd NOR3X1
XOAI21X1_283 gnd NOR2X1_180/B INVX1_189/A gnd INVX1_192/A vdd OAI21X1
XINVX1_104 OR2X2_70/Y gnd INVX1_104/Y vdd INVX1
XBUFX4_29 reset gnd INVX8_1/A vdd BUFX4
XNAND2X1_397 NAND2X1_397/A INVX1_259/Y gnd INVX1_260/A vdd NAND2X1
XAOI22X1_2 INVX4_1/Y INVX2_1/A INVX2_3/Y INVX2_2/A gnd NAND2X1_2/B vdd AOI22X1
XNOR2X1_316 NOR2X1_316/A NOR2X1_316/B gnd NOR2X1_316/Y vdd NOR2X1
XFILL_23_0_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XNOR2X1_83 NOR2X1_83/A NOR3X1_38/Y gnd NOR2X1_83/Y vdd NOR2X1
XNAND3X1_229 AOI21X1_156/A NAND3X1_229/B NAND3X1_229/C gnd AND2X2_78/B vdd NAND3X1
XFILL_21_2_1 gnd vdd FILL
XBUFX2_230 BUFX2_230/A gnd BUFX2_230/Y vdd BUFX2
XFILL_1_3_1 gnd vdd FILL
XOAI21X1_247 NOR3X1_54/Y NOR2X1_163/A NOR3X1_53/Y gnd NAND2X1_290/B vdd OAI21X1
XNOR2X1_280 NOR2X1_280/A NOR2X1_280/B gnd NOR2X1_280/Y vdd NOR2X1
XFILL_11_3 gnd vdd FILL
XNAND2X1_361 NAND2X1_361/A NAND2X1_361/B gnd XOR2X1_187/A vdd NAND2X1
XINVX2_68 INVX2_68/A gnd INVX2_68/Y vdd INVX2
XNAND3X1_193 OAI21X1_183/Y NAND3X1_193/B NAND3X1_193/C gnd AND2X2_66/B vdd NAND3X1
XBUFX2_194 BUFX2_194/A gnd BUFX2_194/Y vdd BUFX2
XNOR2X1_47 NOR2X1_47/A NOR2X1_46/Y gnd XOR2X1_38/A vdd NOR2X1
XXNOR2X1_232 INVX1_575/A bloque_bytes[22] gnd AND2X2_186/B vdd XNOR2X1
XOAI21X1_211 NOR2X1_137/A INVX1_141/Y INVX1_142/Y gnd NAND2X1_247/B vdd OAI21X1
XINVX2_32 INVX2_32/A gnd INVX2_32/Y vdd INVX2
XNOR2X1_244 NOR2X1_244/A NOR2X1_244/B gnd NOR2X1_244/Y vdd NOR2X1
XNAND2X1_325 NAND2X1_325/A NAND3X1_293/B gnd BUFX2_183/A vdd NAND2X1
XNAND3X1_157 NAND3X1_157/A NAND3X1_157/B OAI21X1_151/Y gnd AND2X2_54/B vdd NAND3X1
XBUFX2_158 BUFX2_158/A gnd BUFX2_158/Y vdd BUFX2
XINVX1_573 INVX1_573/A gnd INVX1_573/Y vdd INVX1
XCLKBUF1_35 BUFX4_2/Y gnd CLKBUF1_35/Y vdd CLKBUF1
XFILL_20_5_0 gnd vdd FILL
XOAI21X1_175 INVX2_40/Y AND2X2_60/B OR2X2_78/Y gnd OAI21X1_176/B vdd OAI21X1
XXNOR2X1_196 NOR2X1_326/A NAND2X1_559/Y gnd BUFX2_238/A vdd XNOR2X1
XNOR2X1_11 NAND3X1_2/Y NOR2X1_11/B gnd NOR2X1_11/Y vdd NOR2X1
XXNOR2X1_2 target[3] NOR2X1_4/A gnd NAND2X1_3/A vdd XNOR2X1
XFILL_33_3 gnd vdd FILL
XFILL_0_6_0 gnd vdd FILL
XNAND2X1_289 gnd OR2X2_114/B gnd NAND3X1_259/B vdd NAND2X1
XNOR2X1_208 NOR2X1_208/A NOR2X1_208/B gnd NOR2X1_208/Y vdd NOR2X1
XFILL_18_7_1 gnd vdd FILL
XNOR3X1_88 BUFX4_14/Y NOR3X1_88/B NOR3X1_88/C gnd NOR3X1_88/Y vdd NOR3X1
XDFFPOSX1_355 INVX1_435/A CLKBUF1_40/Y OR2X2_151/Y gnd vdd DFFPOSX1
XBUFX2_122 gnd gnd BUFX2_122/Y vdd BUFX2
XNAND3X1_121 AOI21X1_84/A NAND3X1_120/Y OAI21X1_117/Y gnd AND2X2_42/B vdd NAND3X1
XXNOR2X1_160 NOR2X1_218/A NAND2X1_388/Y gnd BUFX2_202/A vdd XNOR2X1
XBUFX4_4 clk gnd BUFX4_4/Y vdd BUFX4
XINVX1_537 INVX1_537/A gnd INVX1_537/Y vdd INVX1
XXNOR2X1_82 XOR2X1_74/A XOR2X1_78/Y gnd OR2X2_71/A vdd XNOR2X1
XOAI21X1_139 AND2X2_49/Y NOR2X1_94/Y INVX1_92/Y gnd OAI21X1_139/Y vdd OAI21X1
XNOR2X1_172 BUFX2_171/A OR2X2_124/B gnd NOR2X1_172/Y vdd NOR2X1
XFILL_30_0_0 gnd vdd FILL
XFILL_28_2_1 gnd vdd FILL
XFILL_8_3_1 gnd vdd FILL
XNAND2X1_253 INVX1_151/A NAND2X1_253/B gnd OAI21X1_216/A vdd NAND2X1
XNOR3X1_52 INVX1_155/Y NOR3X1_52/B NOR3X1_52/C gnd NOR3X1_52/Y vdd NOR3X1
XINVX1_501 INVX1_501/A gnd INVX1_501/Y vdd INVX1
XDFFPOSX1_319 INVX1_349/A CLKBUF1_39/Y NAND2X1_670/Y gnd vdd DFFPOSX1
XXOR2X1_316 vdd vdd gnd XOR2X1_316/Y vdd XOR2X1
XXNOR2X1_46 BUFX2_249/A XOR2X1_38/Y gnd OR2X2_39/A vdd XNOR2X1
XXNOR2X1_124 XNOR2X1_124/A NAND3X1_240/Y gnd BUFX2_173/A vdd XNOR2X1
XOAI21X1_103 XNOR2X1_53/A AOI21X1_77/C AND2X2_36/B gnd XNOR2X1_54/A vdd OAI21X1
XNAND2X1_217 OR2X2_84/A OR2X2_84/B gnd AOI21X1_136/A vdd NAND2X1
XNOR2X1_136 INVX1_139/Y NOR2X1_136/B gnd NOR2X1_137/B vdd NOR2X1
XDFFPOSX1_283 INVX1_264/A CLKBUF1_32/Y OR2X2_136/A gnd vdd DFFPOSX1
XNOR3X1_16 BUFX4_25/Y MUX2X1_16/Y BUFX4_21/Y gnd NOR3X1_16/Y vdd NOR3X1
XOAI21X1_644 OAI21X1_639/A XNOR2X1_254/B OAI21X1_644/C gnd NAND2X1_712/B vdd OAI21X1
XINVX1_465 INVX1_465/A gnd INVX1_465/Y vdd INVX1
XXNOR2X1_10 vdd XOR2X1_315/Y gnd OR2X2_7/A vdd XNOR2X1
XXOR2X1_280 BUFX2_236/A gnd gnd NOR2X1_347/B vdd XOR2X1
XNOR2X1_100 gnd OR2X2_67/B gnd NOR2X1_100/Y vdd NOR2X1
XNAND2X1_181 AND2X2_54/B AND2X2_54/A gnd AOI21X1_113/C vdd NAND2X1
XAOI21X1_79 NOR2X1_75/Y AOI21X1_79/B INVX1_73/A gnd NOR2X1_77/A vdd AOI21X1
XOR2X2_68 OR2X2_68/A OR2X2_68/B gnd OR2X2_68/Y vdd OR2X2
XDFFPOSX1_247 INVX1_180/A CLKBUF1_21/Y XNOR2X1_234/A gnd vdd DFFPOSX1
XFILL_27_5_0 gnd vdd FILL
XINVX1_429 INVX1_429/A gnd INVX1_429/Y vdd INVX1
XNAND2X1_722 NAND2X1_722/A NAND2X1_722/B gnd XOR2X1_9/A vdd NAND2X1
XFILL_7_6_0 gnd vdd FILL
XOAI21X1_608 INVX1_527/Y bloque_bytes[23] INVX1_528/Y gnd OAI21X1_608/Y vdd OAI21X1
XFILL_25_7_1 gnd vdd FILL
XXOR2X1_244 BUFX2_220/A gnd gnd XOR2X1_244/Y vdd XOR2X1
XFILL_5_8_1 gnd vdd FILL
XBUFX2_82 gnd gnd BUFX2_82/Y vdd BUFX2
XNAND2X1_145 AOI21X1_89/A AOI21X1_89/B gnd INVX2_31/A vdd NAND2X1
XAOI21X1_381 AOI21X1_381/A OR2X2_139/Y AOI21X1_381/C gnd INVX1_561/A vdd AOI21X1
XAOI21X1_43 NOR2X1_45/Y NAND3X1_56/Y INVX1_40/A gnd NOR2X1_47/A vdd AOI21X1
XOR2X2_32 OR2X2_32/A OR2X2_32/B gnd OR2X2_32/Y vdd OR2X2
XOAI21X1_572 INVX4_2/A NOR2X1_388/B INVX1_475/A gnd AOI21X1_327/A vdd OAI21X1
XDFFPOSX1_211 INVX1_132/A CLKBUF1_3/Y OR2X2_143/B gnd vdd DFFPOSX1
XFILL_35_2_1 gnd vdd FILL
XINVX1_393 INVX1_393/A gnd INVX1_393/Y vdd INVX1
XBUFX2_46 gnd gnd BUFX2_46/Y vdd BUFX2
XNAND2X1_686 INVX1_563/A NAND3X1_523/B gnd NAND2X1_686/Y vdd NAND2X1
XXOR2X1_208 BUFX2_204/A gnd gnd XOR2X1_208/Y vdd XOR2X1
XNAND2X1_109 INVX1_61/Y OR2X2_39/A gnd NAND2X1_110/A vdd NAND2X1
XAOI21X1_345 INVX1_492/Y NOR3X1_90/Y INVX1_483/A gnd NOR3X1_93/B vdd AOI21X1
XNAND3X1_518 INVX1_522/Y INVX2_88/Y INVX1_552/A gnd NAND3X1_518/Y vdd NAND3X1
XDFFPOSX1_175 INVX1_81/A CLKBUF1_12/Y bloque_bytes[37] gnd vdd DFFPOSX1
XOAI21X1_91 OAI21X1_91/A OAI21X1_90/Y INVX1_62/Y gnd NAND3X1_94/C vdd OAI21X1
XXOR2X1_172 BUFX2_184/A gnd gnd NOR2X1_203/B vdd XOR2X1
XINVX1_357 INVX1_357/A gnd INVX1_357/Y vdd INVX1
XOAI21X1_536 BUFX2_231/A INVX1_442/A INVX1_443/Y gnd OAI21X1_536/Y vdd OAI21X1
XNAND2X1_650 XNOR2X1_208/Y AOI21X1_370/Y gnd XNOR2X1_235/A vdd NAND2X1
XBUFX2_10 BUFX2_10/A gnd hash[9] vdd BUFX2
XOAI21X1_55 OAI21X1_55/A AOI21X1_46/C NOR2X1_45/Y gnd NOR2X1_46/B vdd OAI21X1
XNAND2X1_70 NAND3X1_55/A OR2X2_24/B gnd OR2X2_22/A vdd NAND2X1
XAOI21X1_309 INVX1_440/A AOI21X1_309/B INVX1_439/Y gnd NOR3X1_83/C vdd AOI21X1
XNAND3X1_482 INVX1_464/A OAI21X1_558/Y NAND2X1_598/Y gnd NAND3X1_482/Y vdd NAND3X1
XDFFPOSX1_139 INVX1_33/A CLKBUF1_33/Y bloque_bytes[65] gnd vdd DFFPOSX1
XDFFPOSX1_73 INVX2_75/A CLKBUF1_24/Y AOI21X1_333/Y gnd vdd DFFPOSX1
XINVX1_321 INVX1_321/A gnd INVX1_321/Y vdd INVX1
XOAI21X1_500 NOR2X1_317/Y NOR2X1_316/B AOI22X1_19/C gnd XOR2X1_269/A vdd OAI21X1
XNAND2X1_614 INVX1_473/A INVX1_475/A gnd OR2X2_129/B vdd NAND2X1
XXOR2X1_136 XOR2X1_136/A OR2X2_108/A gnd AND2X2_89/B vdd XOR2X1
XFILL_34_5_0 gnd vdd FILL
XAOI21X1_273 NAND2X1_486/A NAND2X1_486/B AOI21X1_273/C gnd AOI21X1_273/Y vdd AOI21X1
XFILL_32_7_1 gnd vdd FILL
XNAND2X1_34 NAND2X1_34/A OR2X2_7/Y gnd OR2X2_8/A vdd NAND2X1
XOAI21X1_19 AND2X2_7/Y NOR2X1_24/Y INVX1_15/A gnd NAND3X1_17/B vdd OAI21X1
XDFFPOSX1_37 AOI21X1_353/C CLKBUF1_24/Y AND2X2_163/Y gnd vdd DFFPOSX1
XNAND3X1_446 INVX1_402/A NAND3X1_446/B NAND3X1_441/Y gnd NAND2X1_550/A vdd NAND3X1
XDFFPOSX1_103 INVX2_1/A CLKBUF1_42/Y NOR2X1_438/Y gnd vdd DFFPOSX1
XINVX1_285 NOR3X1_67/B gnd INVX1_285/Y vdd INVX1
XOAI21X1_464 BUFX2_216/A NOR2X1_294/B INVX1_368/A gnd AOI22X1_17/B vdd OAI21X1
XXOR2X1_80 XOR2X1_80/A NOR2X1_91/Y gnd XOR2X1_99/B vdd XOR2X1
XXOR2X1_100 XOR2X1_100/A XOR2X1_100/B gnd BUFX2_158/A vdd XOR2X1
XNAND2X1_578 NAND3X1_464/Y INVX1_446/A gnd NAND2X1_578/Y vdd NAND2X1
XAOI22X1_12 INVX1_276/A AOI22X1_12/B AOI22X1_12/C INVX1_274/A gnd INVX1_280/A vdd
+ AOI22X1
XNAND3X1_410 INVX2_68/A NAND3X1_410/B NAND2X1_497/Y gnd NOR3X1_75/A vdd NAND3X1
XAOI21X1_237 INVX1_269/A AOI21X1_237/B INVX1_268/Y gnd NOR3X1_65/C vdd AOI21X1
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNAND3X1_75 NAND3X1_75/A NAND3X1_75/B XOR2X1_40/B gnd AOI21X1_58/B vdd NAND3X1
XXOR2X1_44 BUFX2_253/A gnd gnd OR2X2_42/B vdd XOR2X1
XAND2X2_180 bloque_bytes[35] INVX1_571/A gnd AND2X2_180/Y vdd AND2X2
XINVX1_249 INVX1_249/A gnd INVX1_249/Y vdd INVX1
XOAI21X1_428 BUFX2_209/A NOR2X1_271/B INVX1_334/A gnd OAI21X1_428/Y vdd OAI21X1
XOR2X2_127 OR2X2_127/A OR2X2_127/B gnd OR2X2_127/Y vdd OR2X2
XNAND2X1_542 INVX1_406/Y NOR2X1_318/Y gnd INVX1_409/A vdd NAND2X1
XAOI21X1_201 INVX2_56/Y XNOR2X1_140/A XNOR2X1_141/A gnd AOI21X1_201/Y vdd AOI21X1
XNAND3X1_374 INVX1_307/A AOI21X1_253/B INVX1_306/Y gnd INVX1_313/A vdd NAND3X1
XINVX1_213 BUFX2_179/A gnd INVX1_213/Y vdd INVX1
XFILL_16_0_1 gnd vdd FILL
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XOAI21X1_392 NOR2X1_245/A NOR3X1_67/Y AOI21X1_249/Y gnd AOI21X1_250/B vdd OAI21X1
XAND2X2_144 AND2X2_144/A NOR3X1_79/A gnd BUFX2_232/A vdd AND2X2
XNAND3X1_39 NAND3X1_39/A XNOR2X1_16/A XOR2X1_20/B gnd NAND3X1_39/Y vdd NAND3X1
XNOR2X1_425 bloque_bytes[38] INVX2_89/A gnd NOR2X1_425/Y vdd NOR2X1
XNAND2X1_506 INVX1_360/A NOR2X1_288/Y gnd NAND2X1_506/Y vdd NAND2X1
XAOI21X1_165 INVX2_47/Y NAND2X1_248/B XNOR2X1_114/A gnd NAND3X1_237/A vdd AOI21X1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XNAND3X1_338 INVX1_255/A NAND3X1_336/Y INVX1_250/Y gnd AOI22X1_11/C vdd NAND3X1
XNOR2X1_389 NOR2X1_398/A INVX2_82/A gnd NOR2X1_389/Y vdd NOR2X1
XAND2X2_108 AND2X2_108/A NOR3X1_61/A gnd BUFX2_192/A vdd AND2X2
XINVX1_177 INVX1_177/A gnd NOR3X1_56/A vdd INVX1
XOAI21X1_356 gnd XOR2X1_189/Y INVX1_263/A gnd OAI21X1_356/Y vdd OAI21X1
XNAND2X1_470 INVX1_334/Y NOR2X1_271/Y gnd NAND2X1_471/B vdd NAND2X1
XNAND3X1_302 INVX1_190/Y NAND2X1_331/A NOR3X1_58/Y gnd NAND3X1_302/Y vdd NAND3X1
XAOI21X1_129 INVX2_38/Y XNOR2X1_85/Y XNOR2X1_87/A gnd AOI21X1_129/Y vdd AOI21X1
XAND2X2_81 gnd AND2X2_81/B gnd NOR3X1_52/C vdd AND2X2
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_141 OR2X2_96/Y gnd INVX1_141/Y vdd INVX1
XOAI21X1_320 NOR3X1_62/C INVX2_61/Y NOR3X1_62/A gnd AND2X2_108/A vdd OAI21X1
XNAND2X1_434 INVX1_295/Y NOR2X1_248/B gnd NAND2X1_435/A vdd NAND2X1
XNOR2X1_353 NOR2X1_353/A NOR3X1_85/Y gnd NOR2X1_353/Y vdd NOR2X1
XFILL_15_3_0 gnd vdd FILL
XNAND3X1_266 INVX1_168/A NAND3X1_264/B OR2X2_116/Y gnd NAND3X1_267/B vdd NAND3X1
XFILL_13_5_1 gnd vdd FILL
XAND2X2_45 gnd OR2X2_58/B gnd AND2X2_45/Y vdd AND2X2
XBUFX2_267 OR2X2_76/A gnd BUFX2_267/Y vdd BUFX2
XNOR3X1_7 BUFX4_27/Y MUX2X1_7/Y BUFX4_20/Y gnd NOR3X1_7/Y vdd NOR3X1
XINVX1_105 INVX1_105/A gnd OR2X2_71/B vdd INVX1
XBUFX4_30 reset gnd BUFX4_30/Y vdd BUFX4
XOAI21X1_284 NOR3X1_57/A NOR3X1_57/B OAI21X1_284/C gnd NOR2X1_182/A vdd OAI21X1
XNAND2X1_398 NAND3X1_342/Y AOI22X1_11/C gnd NAND2X1_398/Y vdd NAND2X1
XAOI22X1_3 INVX1_5/Y target[7] INVX1_6/Y target[6] gnd NAND3X1_2/C vdd AOI22X1
XNOR2X1_317 NOR2X1_317/A NOR3X1_79/Y gnd NOR2X1_317/Y vdd NOR2X1
XNAND3X1_230 INVX1_146/A NAND3X1_228/B OR2X2_100/Y gnd NAND3X1_231/B vdd NAND3X1
XFILL_23_0_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XNOR2X1_84 OR2X2_53/A OR2X2_53/B gnd NOR2X1_84/Y vdd NOR2X1
XBUFX2_231 BUFX2_231/A gnd BUFX2_231/Y vdd BUFX2
XOAI21X1_248 AND2X2_87/Y NOR3X1_54/B INVX1_166/Y gnd NAND3X1_261/B vdd OAI21X1
XNOR2X1_281 NOR2X1_281/A NOR3X1_73/Y gnd NOR2X1_281/Y vdd NOR2X1
XINVX2_69 INVX2_69/A gnd INVX2_69/Y vdd INVX2
XNAND2X1_362 INVX1_225/Y NOR2X1_202/Y gnd NAND3X1_319/B vdd NAND2X1
XBUFX2_195 OR2X2_20/A gnd BUFX2_195/Y vdd BUFX2
XNAND3X1_194 INVX1_124/A AOI21X1_136/A OR2X2_84/Y gnd NAND3X1_194/Y vdd NAND3X1
XNOR2X1_48 gnd OR2X2_25/B gnd NOR3X1_31/B vdd NOR2X1
XFILL_12_8_0 gnd vdd FILL
XXNOR2X1_233 INVX1_543/A bloque_bytes[23] gnd NAND3X1_513/B vdd XNOR2X1
XOAI21X1_212 AND2X2_74/Y NOR3X1_49/B INVX1_143/Y gnd NAND2X1_250/A vdd OAI21X1
XNAND2X1_326 AND2X2_99/B AND2X2_99/A gnd NAND3X1_293/C vdd NAND2X1
XINVX2_33 INVX2_33/A gnd INVX2_33/Y vdd INVX2
XNOR2X1_245 NOR2X1_245/A NOR3X1_67/Y gnd NOR2X1_245/Y vdd NOR2X1
XNAND3X1_158 INVX1_102/A NAND2X1_179/Y OR2X2_68/Y gnd NAND3X1_159/B vdd NAND3X1
XBUFX2_159 AND2X2_77/A gnd BUFX2_159/Y vdd BUFX2
XCLKBUF1_36 BUFX4_3/Y gnd CLKBUF1_36/Y vdd CLKBUF1
XINVX1_574 INVX1_574/A gnd INVX1_574/Y vdd INVX1
XXNOR2X1_3 target[2] NOR2X1_5/A gnd NAND2X1_3/B vdd XNOR2X1
XXNOR2X1_197 NOR2X1_329/Y NOR2X1_328/Y gnd XOR2X1_283/A vdd XNOR2X1
XFILL_20_5_1 gnd vdd FILL
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_176 OAI21X1_176/A OAI21X1_176/B INVX1_117/Y gnd NAND3X1_184/C vdd OAI21X1
XNOR2X1_12 MUX2X1_18/B INVX2_4/Y gnd AOI21X1_8/C vdd NOR2X1
XFILL_0_6_1 gnd vdd FILL
XFILL_2_4_0 gnd vdd FILL
XNAND2X1_290 NAND3X1_260/Y NAND2X1_290/B gnd NAND3X1_273/B vdd NAND2X1
XNOR2X1_209 NOR2X1_209/A NOR3X1_61/Y gnd NOR2X1_209/Y vdd NOR2X1
XNAND3X1_122 INVX1_80/A AOI21X1_88/A OR2X2_52/Y gnd NAND3X1_122/Y vdd NAND3X1
XNOR3X1_89 INVX1_487/Y MUX2X1_3/S NOR3X1_89/C gnd NOR3X1_89/Y vdd NOR3X1
XINVX1_538 INVX1_538/A gnd INVX1_538/Y vdd INVX1
XDFFPOSX1_356 INVX1_436/A CLKBUF1_13/Y NAND2X1_691/Y gnd vdd DFFPOSX1
XXNOR2X1_161 NOR2X1_221/Y NOR2X1_220/Y gnd XOR2X1_202/A vdd XNOR2X1
XBUFX4_5 clk gnd BUFX4_5/Y vdd BUFX4
XBUFX2_123 gnd gnd BUFX2_123/Y vdd BUFX2
XXNOR2X1_83 XOR2X1_91/Y XOR2X1_79/Y gnd XNOR2X1_83/Y vdd XNOR2X1
XNOR2X1_173 NOR2X1_173/A NOR3X1_56/Y gnd NOR2X1_173/Y vdd NOR2X1
XOAI21X1_140 XNOR2X1_71/A OAI21X1_140/B NOR2X1_95/Y gnd NOR2X1_96/B vdd OAI21X1
XFILL_30_0_1 gnd vdd FILL
XNOR3X1_53 INVX1_165/Y NOR3X1_53/B NOR3X1_53/C gnd NOR3X1_53/Y vdd NOR3X1
XNAND2X1_254 gnd OR2X2_99/B gnd NAND3X1_227/B vdd NAND2X1
XINVX1_502 INVX1_502/A gnd INVX1_502/Y vdd INVX1
XDFFPOSX1_320 INVX1_353/A CLKBUF1_32/Y INVX1_566/Y gnd vdd DFFPOSX1
XXNOR2X1_47 XOR2X1_51/Y XOR2X1_39/Y gnd XNOR2X1_47/Y vdd XNOR2X1
XXOR2X1_317 XOR2X1_317/A XOR2X1_317/B gnd XOR2X1_5/A vdd XOR2X1
XOAI21X1_104 AND2X2_37/Y NOR2X1_74/Y INVX1_70/A gnd NAND3X1_107/B vdd OAI21X1
XXNOR2X1_125 XNOR2X1_125/A AND2X2_84/Y gnd XOR2X1_146/A vdd XNOR2X1
XNAND2X1_218 INVX2_42/Y NAND3X1_200/C gnd XNOR2X1_98/A vdd NAND2X1
XNOR2X1_137 NOR2X1_137/A NOR2X1_137/B gnd XOR2X1_128/A vdd NOR2X1
XFILL_19_8_0 gnd vdd FILL
XDFFPOSX1_284 INVX1_265/A CLKBUF1_23/Y NOR2X1_427/B gnd vdd DFFPOSX1
XNOR3X1_17 NOR3X1_9/A MUX2X1_17/Y NOR3X1_9/C gnd NOR3X1_17/Y vdd NOR3X1
XOAI21X1_645 XNOR2X1_255/A AOI21X1_400/C AND2X2_197/B gnd XNOR2X1_256/A vdd OAI21X1
XXOR2X1_281 BUFX2_237/A gnd gnd NOR2X1_348/B vdd XOR2X1
XINVX1_466 INVX1_466/A gnd INVX1_466/Y vdd INVX1
XXNOR2X1_11 XOR2X1_11/Y XOR2X1_316/Y gnd XNOR2X1_12/A vdd XNOR2X1
XNOR2X1_101 NOR2X1_101/A INVX2_36/A gnd XOR2X1_90/B vdd NOR2X1
XFILL_15_1 gnd vdd FILL
XNAND2X1_182 OR2X2_69/A OR2X2_69/B gnd NAND3X1_162/B vdd NAND2X1
XFILL_29_3_0 gnd vdd FILL
XOR2X2_69 OR2X2_69/A OR2X2_69/B gnd OR2X2_69/Y vdd OR2X2
XFILL_9_4_0 gnd vdd FILL
XAOI21X1_80 INVX2_27/Y INVX1_74/Y NOR2X1_71/A gnd AOI21X1_82/A vdd AOI21X1
XDFFPOSX1_248 INVX1_182/A CLKBUF1_21/Y OR2X2_140/A gnd vdd DFFPOSX1
XOAI21X1_609 INVX1_530/Y bloque_bytes[34] INVX1_531/Y gnd AOI21X1_372/C vdd OAI21X1
XFILL_27_5_1 gnd vdd FILL
XINVX1_430 INVX1_430/A gnd INVX1_430/Y vdd INVX1
XFILL_7_6_1 gnd vdd FILL
XBUFX2_83 gnd gnd BUFX2_83/Y vdd BUFX2
XXOR2X1_245 BUFX2_221/A gnd gnd NOR2X1_300/B vdd XOR2X1
XNAND2X1_146 OAI21X1_122/Y OR2X2_56/B gnd OR2X2_54/A vdd NAND2X1
XAOI21X1_382 AOI21X1_382/A AOI21X1_382/B AOI21X1_382/C gnd INVX1_563/A vdd AOI21X1
XDFFPOSX1_212 INVX1_133/A CLKBUF1_10/Y INVX1_544/A gnd vdd DFFPOSX1
XAOI21X1_44 INVX2_18/Y INVX1_41/Y NOR2X1_41/A gnd AOI21X1_44/Y vdd AOI21X1
XOR2X2_33 gnd OR2X2_33/B gnd OR2X2_33/Y vdd OR2X2
XOAI21X1_573 INVX2_82/Y AND2X2_161/B BUFX4_31/Y gnd AOI21X1_328/C vdd OAI21X1
XFILL_37_1 gnd vdd FILL
XINVX1_394 INVX1_394/A gnd INVX1_394/Y vdd INVX1
XBUFX2_47 gnd gnd BUFX2_47/Y vdd BUFX2
XNAND2X1_687 INVX1_565/A XNOR2X1_238/Y gnd NAND2X1_687/Y vdd NAND2X1
XXOR2X1_209 BUFX2_205/A gnd gnd NOR2X1_252/B vdd XOR2X1
XNAND2X1_110 NAND2X1_110/A OR2X2_39/Y gnd OR2X2_40/A vdd NAND2X1
XAOI21X1_346 INVX1_484/Y AOI21X1_346/B NAND2X1_635/Y gnd DFFPOSX1_86/D vdd AOI21X1
XNAND3X1_519 INVX1_525/Y INVX2_89/Y INVX1_553/A gnd NAND3X1_519/Y vdd NAND3X1
XOAI21X1_92 NOR2X1_67/A INVX1_64/Y INVX1_65/Y gnd OAI21X1_92/Y vdd OAI21X1
XDFFPOSX1_176 INVX1_83/A CLKBUF1_12/Y bloque_bytes[38] gnd vdd DFFPOSX1
XXOR2X1_173 BUFX2_185/A gnd gnd NOR2X1_204/B vdd XOR2X1
XNAND2X1_651 XNOR2X1_209/Y AOI21X1_371/Y gnd XNOR2X1_236/A vdd NAND2X1
XINVX1_358 INVX1_358/A gnd INVX1_358/Y vdd INVX1
XOAI21X1_537 NOR3X1_83/C OAI21X1_537/B INVX1_446/A gnd NOR2X1_341/A vdd OAI21X1
XFILL_26_8_0 gnd vdd FILL
XBUFX2_11 BUFX2_11/A gnd hash[10] vdd BUFX2
XOAI21X1_56 INVX2_19/Y AND2X2_18/B INVX1_38/A gnd OAI21X1_56/Y vdd OAI21X1
XNAND2X1_71 OR2X2_23/B OR2X2_23/A gnd NAND2X1_72/A vdd NAND2X1
XFILL_6_9_0 gnd vdd FILL
XDFFPOSX1_74 INVX2_76/A CLKBUF1_3/Y AND2X2_170/Y gnd vdd DFFPOSX1
XAOI21X1_310 AOI21X1_310/A AOI21X1_310/B INVX2_72/A gnd AOI21X1_311/B vdd AOI21X1
XNAND3X1_483 AOI22X1_22/B INVX1_466/A INVX1_464/Y gnd NAND3X1_483/Y vdd NAND3X1
XDFFPOSX1_140 INVX1_34/A CLKBUF1_7/Y bloque_bytes[66] gnd vdd DFFPOSX1
XINVX1_322 INVX1_322/A gnd INVX1_322/Y vdd INVX1
XOAI21X1_501 BUFX2_224/A XOR2X1_257/Y INVX1_406/Y gnd OAI21X1_501/Y vdd OAI21X1
XNAND2X1_615 AND2X2_159/B INVX2_74/A gnd NOR2X1_388/A vdd NAND2X1
XXOR2X1_137 XOR2X1_137/A BUFX2_164/A gnd OR2X2_117/B vdd XOR2X1
XFILL_36_3_0 gnd vdd FILL
XFILL_34_5_1 gnd vdd FILL
XNAND2X1_35 OR2X2_8/B OR2X2_8/A gnd NAND2X1_36/A vdd NAND2X1
XAOI21X1_274 INVX1_356/Y OAI21X1_449/Y INVX1_355/A gnd OAI21X1_450/A vdd AOI21X1
XOAI21X1_20 AND2X2_7/Y NOR2X1_24/Y INVX1_15/Y gnd NAND3X1_19/A vdd OAI21X1
XDFFPOSX1_38 AOI21X1_354/C CLKBUF1_14/Y NOR2X1_364/Y gnd vdd DFFPOSX1
XNAND3X1_447 INVX1_413/Y INVX1_412/A NAND3X1_447/C gnd AND2X2_145/B vdd NAND3X1
XDFFPOSX1_104 XOR2X1_1/B CLKBUF1_28/Y XOR2X1_306/Y gnd vdd DFFPOSX1
XXOR2X1_81 BUFX2_262/A XOR2X1_81/B gnd XOR2X1_81/Y vdd XOR2X1
XXOR2X1_101 XOR2X1_99/B XOR2X1_101/B gnd XOR2X1_101/Y vdd XOR2X1
XINVX1_286 INVX1_286/A gnd INVX1_286/Y vdd INVX1
XOAI21X1_465 gnd XOR2X1_236/Y INVX1_360/Y gnd OAI21X1_465/Y vdd OAI21X1
XNAND2X1_579 INVX1_444/A NOR2X1_342/Y gnd NAND2X1_579/Y vdd NAND2X1
XAOI22X1_13 INVX1_295/A AOI22X1_13/B AOI22X1_13/C INVX1_293/A gnd INVX1_299/A vdd
+ AOI22X1
XAOI21X1_238 AOI21X1_238/A AOI21X1_238/B INVX2_63/A gnd AOI21X1_239/B vdd AOI21X1
XNAND3X1_411 INVX1_363/A NAND2X1_499/B INVX2_68/Y gnd OAI21X1_461/B vdd NAND3X1
XAND2X2_7 vdd OR2X2_5/B gnd AND2X2_7/Y vdd AND2X2
XFILL_10_1_0 gnd vdd FILL
XINVX1_250 INVX1_250/A gnd INVX1_250/Y vdd INVX1
XOAI21X1_429 AOI21X1_264/Y INVX1_337/A INVX1_336/Y gnd AND2X2_129/A vdd OAI21X1
XFILL_2_2 gnd vdd FILL
XNAND3X1_76 OR2X2_32/Y INVX1_54/A OAI21X1_74/Y gnd NAND2X1_95/A vdd NAND3X1
XXOR2X1_45 XOR2X1_61/A gnd gnd OR2X2_43/B vdd XOR2X1
XAND2X2_181 bloque_bytes[36] INVX1_572/A gnd AND2X2_181/Y vdd AND2X2
XNAND2X1_543 NAND3X1_443/Y NAND3X1_444/Y gnd XOR2X1_269/B vdd NAND2X1
XOR2X2_128 OR2X2_128/A OR2X2_128/B gnd INVX1_185/A vdd OR2X2
XAOI21X1_202 AOI21X1_202/A AOI21X1_202/B NAND2X1_322/Y gnd OAI21X1_278/A vdd AOI21X1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XFILL_33_8_0 gnd vdd FILL
XNAND3X1_375 INVX1_308/Y INVX1_309/Y INVX1_310/Y gnd NAND3X1_375/Y vdd NAND3X1
XINVX1_214 INVX1_214/A gnd INVX1_214/Y vdd INVX1
XOAI21X1_393 OAI21X1_393/A INVX1_297/A INVX1_300/A gnd NAND2X1_437/A vdd OAI21X1
XAND2X2_145 AND2X2_145/A AND2X2_145/B gnd XOR2X1_276/A vdd AND2X2
XNAND3X1_40 INVX1_31/A INVX1_32/A OAI21X1_40/Y gnd NAND2X1_57/A vdd NAND3X1
XNOR2X1_426 NOR2X1_426/A NOR2X1_426/B gnd INVX1_546/A vdd NOR2X1
XNAND2X1_507 XOR2X1_251/B NOR2X1_292/Y gnd NAND2X1_507/Y vdd NAND2X1
XAOI21X1_166 AOI21X1_166/A AOI21X1_166/B AOI21X1_166/C gnd OAI21X1_227/A vdd AOI21X1
XNAND3X1_339 INVX1_255/A NAND3X1_339/B NAND3X1_339/C gnd AOI21X1_233/A vdd NAND3X1
XINVX1_60 OR2X2_38/Y gnd INVX1_60/Y vdd INVX1
XAND2X2_109 AND2X2_109/A AND2X2_109/B gnd AND2X2_109/Y vdd AND2X2
XNOR2X1_390 INVX1_488/A INVX2_82/A gnd NOR2X1_390/Y vdd NOR2X1
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XOAI21X1_357 gnd XOR2X1_190/Y INVX1_264/A gnd INVX2_63/A vdd OAI21X1
XNAND2X1_471 OAI21X1_428/Y NAND2X1_471/B gnd NOR2X1_272/B vdd NAND2X1
XNAND3X1_303 INVX1_193/A AOI21X1_204/A AOI21X1_204/B gnd NAND2X1_341/A vdd NAND3X1
XAND2X2_82 gnd AND2X2_82/B gnd AND2X2_82/Y vdd AND2X2
XAOI21X1_130 AOI21X1_130/A AOI21X1_130/B OAI21X1_174/B gnd OAI21X1_176/A vdd AOI21X1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XOAI21X1_321 gnd NOR2X1_204/B INVX1_227/A gnd INVX1_230/A vdd OAI21X1
XINVX1_142 INVX1_142/A gnd INVX1_142/Y vdd INVX1
XFILL_17_1_0 gnd vdd FILL
XNAND2X1_435 NAND2X1_435/A INVX1_297/Y gnd INVX1_298/A vdd NAND2X1
XNOR2X1_354 BUFX2_236/A XOR2X1_284/Y gnd NOR2X1_354/Y vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XAND2X2_46 gnd OR2X2_59/B gnd AND2X2_46/Y vdd AND2X2
XNOR3X1_8 NOR3X1_2/A NOR3X1_8/B NOR3X1_2/C gnd NOR3X1_8/Y vdd NOR3X1
XNAND3X1_267 NAND3X1_267/A NAND3X1_267/B AOI21X1_182/Y gnd AND2X2_90/A vdd NAND3X1
XBUFX2_268 OR2X2_77/A gnd BUFX2_268/Y vdd BUFX2
XINVX1_106 INVX1_106/A gnd INVX1_106/Y vdd INVX1
XOAI21X1_285 NOR3X1_58/A NOR3X1_58/C INVX2_59/A gnd NOR2X1_181/A vdd OAI21X1
XBUFX4_31 reset gnd BUFX4_31/Y vdd BUFX4
XNOR2X1_318 BUFX2_224/A XOR2X1_257/Y gnd NOR2X1_318/Y vdd NOR2X1
XNAND2X1_399 OAI21X1_355/Y NAND3X1_344/Y gnd XOR2X1_205/A vdd NAND2X1
XAOI22X1_4 INVX1_7/Y target[5] INVX1_8/Y target[4] gnd AOI21X1_7/C vdd AOI22X1
XAND2X2_10 gnd OR2X2_11/B gnd AND2X2_10/Y vdd AND2X2
XNAND3X1_231 NAND3X1_233/A NAND3X1_231/B NAND3X1_231/C gnd AND2X2_78/A vdd NAND3X1
XBUFX2_232 BUFX2_232/A gnd BUFX2_232/Y vdd BUFX2
XNOR2X1_85 NOR2X1_85/A INVX1_82/Y gnd NOR2X1_85/Y vdd NOR2X1
XOAI21X1_249 NOR3X1_54/Y NOR2X1_163/A NAND3X1_260/B gnd OAI21X1_249/Y vdd OAI21X1
XNAND2X1_363 NAND2X1_363/A NAND3X1_319/B gnd BUFX2_191/A vdd NAND2X1
XINVX2_70 INVX2_70/A gnd INVX2_70/Y vdd INVX2
XNOR2X1_282 BUFX2_212/A XOR2X1_230/Y gnd NOR2X1_282/Y vdd NOR2X1
XBUFX2_196 OR2X2_21/A gnd BUFX2_196/Y vdd BUFX2
XNAND3X1_195 NAND3X1_197/A NAND3X1_194/Y AOI21X1_134/Y gnd AND2X2_66/A vdd NAND3X1
XNOR2X1_49 gnd OR2X2_26/B gnd NOR2X1_49/Y vdd NOR2X1
XFILL_12_8_1 gnd vdd FILL
XFILL_14_6_0 gnd vdd FILL
XXNOR2X1_234 XNOR2X1_234/A bloque_bytes[5] gnd XNOR2X1_234/Y vdd XNOR2X1
XOAI21X1_213 NOR3X1_50/Y NOR2X1_143/A NOR3X1_49/Y gnd NAND2X1_252/B vdd OAI21X1
XNAND2X1_327 INVX1_189/Y NOR2X1_180/Y gnd NAND2X1_328/B vdd NAND2X1
XINVX2_34 INVX2_34/A gnd INVX2_34/Y vdd INVX2
XNOR2X1_246 BUFX2_200/A XOR2X1_203/Y gnd NOR2X1_246/Y vdd NOR2X1
XNAND3X1_159 NAND3X1_161/A NAND3X1_159/B NAND3X1_159/C gnd AND2X2_54/A vdd NAND3X1
XXNOR2X1_4 gnd XNOR2X1_4/B gnd XNOR2X1_5/A vdd XNOR2X1
XCLKBUF1_37 BUFX4_6/Y gnd CLKBUF1_37/Y vdd CLKBUF1
XINVX1_575 INVX1_575/A gnd INVX1_575/Y vdd INVX1
XBUFX2_160 OR2X2_101/A gnd BUFX2_160/Y vdd BUFX2
XFILL_22_3_1 gnd vdd FILL
XFILL_24_1_0 gnd vdd FILL
XNOR2X1_13 OAI22X1_6/Y NOR2X1_13/B gnd NOR2X1_13/Y vdd NOR2X1
XXNOR2X1_198 NOR2X1_333/Y XNOR2X1_198/B gnd XNOR2X1_199/A vdd XNOR2X1
XFILL_2_4_1 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XNOR2X1_210 BUFX2_184/A NOR2X1_210/B gnd NOR2X1_210/Y vdd NOR2X1
XOAI21X1_177 NOR2X1_117/A INVX1_119/Y INVX1_120/Y gnd NAND2X1_209/B vdd OAI21X1
XNOR3X1_90 INVX2_84/A INVX1_491/A NOR3X1_90/C gnd NOR3X1_90/Y vdd NOR3X1
XNAND2X1_291 INVX1_173/A OAI21X1_249/Y gnd OAI21X1_250/A vdd NAND2X1
XINVX4_1 target[5] gnd INVX4_1/Y vdd INVX4
XNAND3X1_123 NAND3X1_123/A NAND3X1_122/Y AOI21X1_86/Y gnd AND2X2_42/A vdd NAND3X1
XBUFX2_124 gnd gnd BUFX2_124/Y vdd BUFX2
XINVX1_539 INVX1_539/A gnd INVX1_539/Y vdd INVX1
XDFFPOSX1_357 INVX1_438/A CLKBUF1_40/Y OR2X2_152/Y gnd vdd DFFPOSX1
XXNOR2X1_84 XNOR2X1_83/Y OR2X2_71/Y gnd INVX1_109/A vdd XNOR2X1
XBUFX4_6 clk gnd BUFX4_6/Y vdd BUFX4
XXNOR2X1_162 NOR2X1_225/Y XNOR2X1_162/B gnd XNOR2X1_163/A vdd XNOR2X1
XOAI21X1_141 INVX2_34/Y AND2X2_48/B OR2X2_62/Y gnd OAI21X1_141/Y vdd OAI21X1
XNAND2X1_255 AND2X2_77/A AND2X2_77/B gnd NAND3X1_228/B vdd NAND2X1
XNOR2X1_174 OR2X2_125/A OR2X2_125/B gnd NOR2X1_174/Y vdd NOR2X1
XNOR3X1_54 INVX1_166/Y NOR3X1_54/B AND2X2_87/Y gnd NOR3X1_54/Y vdd NOR3X1
XDFFPOSX1_321 XNOR2X1_182/B CLKBUF1_34/Y INVX1_567/Y gnd vdd DFFPOSX1
XXOR2X1_318 vdd XOR2X1_318/B gnd XOR2X1_318/Y vdd XOR2X1
XINVX1_503 INVX1_503/A gnd INVX1_503/Y vdd INVX1
XXNOR2X1_126 XNOR2X1_126/A INVX2_52/Y gnd XOR2X1_147/A vdd XNOR2X1
XXNOR2X1_48 XNOR2X1_47/Y OR2X2_39/Y gnd INVX1_65/A vdd XNOR2X1
XOAI21X1_105 AND2X2_37/Y NOR2X1_74/Y INVX1_70/Y gnd OAI21X1_105/Y vdd OAI21X1
XNOR2X1_138 gnd OR2X2_97/B gnd NOR3X1_49/B vdd NOR2X1
XFILL_21_6_0 gnd vdd FILL
XNAND2X1_219 AND2X2_66/B AND2X2_66/A gnd AOI21X1_137/C vdd NAND2X1
XFILL_1_7_0 gnd vdd FILL
XFILL_19_8_1 gnd vdd FILL
XDFFPOSX1_285 INVX1_267/A CLKBUF1_23/Y OR2X2_137/A gnd vdd DFFPOSX1
XNOR3X1_18 NOR3X1_9/A MUX2X1_18/Y NOR3X1_9/C gnd NOR3X1_18/Y vdd NOR3X1
XINVX1_467 INVX1_467/A gnd INVX1_467/Y vdd INVX1
XOAI21X1_646 AND2X2_198/Y NOR2X1_451/Y INVX1_594/A gnd NAND3X1_544/B vdd OAI21X1
XXOR2X1_282 BUFX2_238/A gnd gnd XOR2X1_282/Y vdd XOR2X1
XXNOR2X1_12 XNOR2X1_12/A OR2X2_7/Y gnd INVX1_21/A vdd XNOR2X1
XNOR2X1_102 OR2X2_68/A OR2X2_68/B gnd NOR2X1_102/Y vdd NOR2X1
XFILL_31_1_0 gnd vdd FILL
XNAND2X1_183 NAND3X1_161/Y NAND3X1_163/Y gnd INVX2_37/A vdd NAND2X1
XFILL_29_3_1 gnd vdd FILL
XOR2X2_70 OR2X2_70/A OR2X2_70/B gnd OR2X2_70/Y vdd OR2X2
XFILL_9_4_1 gnd vdd FILL
XAOI21X1_81 INVX2_26/Y AOI21X1_81/B AOI21X1_81/C gnd AOI21X1_81/Y vdd AOI21X1
XDFFPOSX1_249 XOR2X1_161/B CLKBUF1_21/Y OR2X2_141/A gnd vdd DFFPOSX1
XOAI21X1_610 INVX1_532/Y bloque_bytes[37] INVX1_533/Y gnd AOI21X1_375/C vdd OAI21X1
XINVX1_431 INVX1_431/A gnd INVX1_431/Y vdd INVX1
XBUFX2_84 gnd gnd BUFX2_84/Y vdd BUFX2
XXOR2X1_246 BUFX2_222/A gnd gnd XOR2X1_246/Y vdd XOR2X1
XNAND2X1_147 OR2X2_55/B OR2X2_55/A gnd NAND2X1_147/Y vdd NAND2X1
XAOI21X1_383 AOI21X1_383/A AOI21X1_383/B XNOR2X1_242/A gnd INVX1_565/A vdd AOI21X1
XAOI21X1_45 INVX2_17/Y NAND2X1_58/B NAND2X1_60/Y gnd NAND3X1_57/A vdd AOI21X1
XDFFPOSX1_213 INVX1_134/A CLKBUF1_50/Y INVX1_571/A gnd vdd DFFPOSX1
XOR2X2_34 gnd OR2X2_34/B gnd OR2X2_34/Y vdd OR2X2
XOAI21X1_574 INVX2_82/A NOR2X1_398/A BUFX4_31/Y gnd OAI21X1_574/Y vdd OAI21X1
XINVX1_395 INVX1_395/A gnd INVX1_395/Y vdd INVX1
XXOR2X1_210 BUFX2_206/A gnd gnd XOR2X1_210/Y vdd XOR2X1
XBUFX2_48 gnd gnd BUFX2_48/Y vdd BUFX2
XNAND2X1_688 NAND2X1_688/A NAND2X1_688/B gnd NAND3X1_526/B vdd NAND2X1
XNAND2X1_111 OR2X2_40/B OR2X2_40/A gnd NAND2X1_112/A vdd NAND2X1
XOAI21X1_93 NOR3X1_35/C NOR3X1_35/B INVX1_66/Y gnd OAI21X1_93/Y vdd OAI21X1
XAOI21X1_347 INVX2_80/Y NAND3X1_501/Y AOI21X1_347/C gnd DFFPOSX1_87/D vdd AOI21X1
XNAND3X1_520 INVX1_558/A XNOR2X1_235/Y XNOR2X1_239/Y gnd NAND3X1_520/Y vdd NAND3X1
XDFFPOSX1_177 XOR2X1_71/B CLKBUF1_29/Y bloque_bytes[39] gnd vdd DFFPOSX1
XINVX1_359 INVX1_359/A gnd INVX1_359/Y vdd INVX1
XOAI21X1_538 NOR2X1_341/Y NOR2X1_340/B AOI22X1_21/C gnd XOR2X1_287/A vdd OAI21X1
XXOR2X1_174 BUFX2_186/A gnd gnd NOR2X1_207/B vdd XOR2X1
XNAND2X1_652 XNOR2X1_210/Y NAND2X1_652/B gnd NAND2X1_652/Y vdd NAND2X1
XFILL_26_8_1 gnd vdd FILL
XBUFX2_12 BUFX2_12/A gnd hash[11] vdd BUFX2
XFILL_28_6_0 gnd vdd FILL
XFILL_6_9_1 gnd vdd FILL
XFILL_8_7_0 gnd vdd FILL
XAOI21X1_311 NAND3X1_464/Y AOI21X1_311/B INVX1_446/Y gnd AOI21X1_312/A vdd AOI21X1
XOAI21X1_57 AOI21X1_46/Y OAI21X1_56/Y INVX1_40/Y gnd OAI21X1_57/Y vdd OAI21X1
XNAND2X1_72 NAND2X1_72/A OR2X2_23/Y gnd OR2X2_24/A vdd NAND2X1
XDFFPOSX1_141 INVX1_35/A CLKBUF1_7/Y bloque_bytes[67] gnd vdd DFFPOSX1
XDFFPOSX1_75 AND2X2_165/B CLKBUF1_3/Y NOR2X1_401/Y gnd vdd DFFPOSX1
XNAND3X1_484 INVX1_456/Y NAND3X1_477/Y NOR3X1_86/Y gnd AOI21X1_320/B vdd NAND3X1
XINVX1_323 NOR3X1_71/B gnd INVX1_323/Y vdd INVX1
XOAI21X1_502 BUFX2_224/A XOR2X1_257/Y INVX1_406/A gnd AOI22X1_19/B vdd OAI21X1
XXOR2X1_138 XOR2X1_138/A BUFX2_165/A gnd XOR2X1_138/Y vdd XOR2X1
XNAND2X1_616 AND2X2_161/B INVX2_82/Y gnd NAND2X1_616/Y vdd NAND2X1
XFILL_36_3_1 gnd vdd FILL
XNAND2X1_36 NAND2X1_36/A OR2X2_8/Y gnd INVX1_18/A vdd NAND2X1
XAOI21X1_275 INVX1_369/A AOI21X1_275/B INVX1_364/Y gnd NOR2X1_292/B vdd AOI21X1
XNAND3X1_448 INVX1_411/Y INVX1_414/Y AND2X2_145/A gnd NAND2X1_551/B vdd NAND3X1
XOAI21X1_21 XNOR2X1_8/A OAI21X1_21/B NOR2X1_25/Y gnd NOR2X1_26/B vdd OAI21X1
XDFFPOSX1_39 INVX1_574/A CLKBUF1_9/Y AND2X2_164/Y gnd vdd DFFPOSX1
XDFFPOSX1_105 NOR2X1_1/B CLKBUF1_28/Y XOR2X1_307/Y gnd vdd DFFPOSX1
XXOR2X1_102 OR2X2_92/A gnd gnd XOR2X1_102/Y vdd XOR2X1
XINVX1_287 INVX1_287/A gnd INVX1_287/Y vdd INVX1
XXOR2X1_82 OR2X2_76/A gnd gnd XOR2X1_82/Y vdd XOR2X1
XOAI21X1_466 BUFX2_217/A XOR2X1_240/Y INVX1_372/A gnd OAI21X1_466/Y vdd OAI21X1
XAOI22X1_14 INVX1_314/A AOI22X1_14/B AOI22X1_14/C INVX1_312/A gnd INVX1_318/A vdd
+ AOI22X1
XNAND2X1_580 INVX1_444/Y NOR2X1_342/Y gnd INVX1_447/A vdd NAND2X1
XAOI21X1_239 NAND3X1_347/Y AOI21X1_239/B INVX1_275/Y gnd AOI21X1_240/A vdd AOI21X1
XNAND3X1_412 INVX1_363/A OAI21X1_457/Y NAND3X1_412/C gnd NAND3X1_419/B vdd NAND3X1
XAND2X2_8 gnd OR2X2_9/B gnd AND2X2_8/Y vdd AND2X2
XFILL_2_3 gnd vdd FILL
XFILL_10_1_1 gnd vdd FILL
XAND2X2_182 INVX1_529/A AND2X2_182/B gnd INVX1_545/A vdd AND2X2
XINVX1_251 INVX1_251/A gnd INVX1_251/Y vdd INVX1
XOAI21X1_430 NOR2X1_269/A NOR3X1_71/Y AOI21X1_265/Y gnd AOI21X1_266/B vdd OAI21X1
XXOR2X1_46 XOR2X1_46/A OR2X2_36/A gnd OR2X2_44/B vdd XOR2X1
XNAND3X1_77 INVX1_55/A NAND2X1_97/Y OR2X2_33/Y gnd NAND3X1_77/Y vdd NAND3X1
XOR2X2_129 OR2X2_129/A OR2X2_129/B gnd OR2X2_129/Y vdd OR2X2
XNAND2X1_544 INVX1_398/A NOR2X1_312/Y gnd AOI21X1_294/B vdd NAND2X1
XAOI21X1_203 AOI22X1_8/D AOI21X1_203/B INVX1_193/Y gnd NOR2X1_184/B vdd AOI21X1
XFILL_35_6_0 gnd vdd FILL
XINVX1_97 OR2X2_64/Y gnd INVX1_97/Y vdd INVX1
XFILL_33_8_1 gnd vdd FILL
XNAND3X1_376 INVX1_310/A INVX1_308/Y INVX1_309/Y gnd AOI21X1_252/B vdd NAND3X1
XXOR2X1_10 XOR2X1_10/A XOR2X1_10/B gnd XOR2X1_15/A vdd XOR2X1
XINVX1_215 INVX1_215/A gnd INVX1_215/Y vdd INVX1
XNOR2X1_427 bloque_bytes[10] NOR2X1_427/B gnd INVX1_554/A vdd NOR2X1
XAND2X2_146 AND2X2_146/A INVX1_415/Y gnd NOR3X1_82/A vdd AND2X2
XOAI21X1_394 gnd XOR2X1_207/Y INVX1_301/A gnd OAI21X1_394/Y vdd OAI21X1
XNAND3X1_41 INVX1_33/A NAND3X1_41/B OR2X2_17/Y gnd NAND3X1_42/A vdd NAND3X1
XNAND2X1_508 INVX1_372/Y NOR2X1_295/Y gnd NAND2X1_508/Y vdd NAND2X1
XNAND3X1_340 AOI22X1_11/B INVX1_257/A INVX1_255/Y gnd AOI21X1_233/B vdd NAND3X1
XAOI21X1_167 AOI21X1_167/A OR2X2_106/Y INVX1_155/A gnd NOR2X1_153/A vdd AOI21X1
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XINVX1_179 INVX1_179/A gnd INVX1_179/Y vdd INVX1
XNOR2X1_391 AND2X2_163/B NOR2X1_390/Y gnd NOR2X1_391/Y vdd NOR2X1
XAND2X2_110 AND2X2_110/A INVX1_244/Y gnd NOR3X1_64/A vdd AND2X2
XOAI21X1_358 NOR3X1_66/C INVX2_63/Y NOR3X1_66/A gnd AND2X2_116/A vdd OAI21X1
XNAND2X1_472 INVX1_333/Y NOR2X1_272/B gnd NAND2X1_473/A vdd NAND2X1
XAOI21X1_131 NAND3X1_187/B OR2X2_82/Y INVX1_122/A gnd NOR2X1_123/A vdd AOI21X1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XNAND3X1_304 INVX1_204/Y INVX1_203/A OAI21X1_297/Y gnd AND2X2_101/B vdd NAND3X1
XAND2X2_83 OR2X2_108/A OR2X2_108/B gnd AND2X2_83/Y vdd AND2X2
XOAI21X1_322 NOR3X1_61/A NOR3X1_61/B OAI21X1_328/B gnd NOR2X1_206/A vdd OAI21X1
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XFILL_17_1_1 gnd vdd FILL
XNAND2X1_436 NAND2X1_436/A AOI22X1_13/C gnd NAND2X1_436/Y vdd NAND2X1
XNOR2X1_355 BUFX2_237/A NOR2X1_355/B gnd NOR2X1_355/Y vdd NOR2X1
XNAND3X1_268 INVX1_169/Y NAND3X1_270/B OR2X2_117/Y gnd NAND3X1_269/C vdd NAND3X1
XAND2X2_47 OR2X2_60/A OR2X2_60/B gnd AND2X2_47/Y vdd AND2X2
XNOR3X1_9 NOR3X1_9/A MUX2X1_9/Y NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XBUFX2_269 XOR2X1_98/B gnd BUFX2_269/Y vdd BUFX2
XINVX1_107 INVX1_107/A gnd INVX1_107/Y vdd INVX1
XOAI21X1_286 gnd NOR2X1_183/B INVX1_191/Y gnd NAND3X1_295/B vdd OAI21X1
XBUFX4_32 reset gnd BUFX4_32/Y vdd BUFX4
XNOR2X1_319 BUFX2_225/A NOR2X1_319/B gnd NOR2X1_319/Y vdd NOR2X1
XNAND2X1_400 INVX1_263/Y AND2X2_114/A gnd NAND3X1_345/B vdd NAND2X1
XAOI22X1_5 INVX2_10/Y target[3] INVX1_9/Y target[2] gnd AOI22X1_5/Y vdd AOI22X1
XAND2X2_11 XOR2X1_2/A OR2X2_12/B gnd AND2X2_11/Y vdd AND2X2
XNAND3X1_232 INVX1_147/Y NAND3X1_234/B OR2X2_101/Y gnd NAND3X1_233/C vdd NAND3X1
XBUFX2_233 BUFX2_233/A gnd BUFX2_233/Y vdd BUFX2
XNOR2X1_86 INVX1_84/Y NOR2X1_86/B gnd NOR2X1_87/B vdd NOR2X1
XOAI21X1_250 OAI21X1_250/A NAND3X1_258/Y INVX1_173/A gnd XOR2X1_150/A vdd OAI21X1
XNAND2X1_364 INVX1_226/Y AND2X2_107/A gnd NAND3X1_319/C vdd NAND2X1
XINVX2_71 INVX2_71/A gnd INVX2_71/Y vdd INVX2
XNOR2X1_283 BUFX2_213/A XOR2X1_231/Y gnd NOR2X1_283/Y vdd NOR2X1
XFILL_28_1 gnd vdd FILL
XBUFX2_197 XOR2X1_28/B gnd BUFX2_197/Y vdd BUFX2
XNOR2X1_50 gnd OR2X2_27/B gnd NOR2X1_50/Y vdd NOR2X1
XNAND3X1_196 INVX1_125/Y NAND2X1_220/Y OR2X2_85/Y gnd NAND3X1_196/Y vdd NAND3X1
XFILL_14_6_1 gnd vdd FILL
XFILL_16_4_0 gnd vdd FILL
XXNOR2X1_235 XNOR2X1_235/A NOR2X1_410/A gnd XNOR2X1_235/Y vdd XNOR2X1
XOAI21X1_214 NOR3X1_50/C NOR3X1_50/B INVX1_144/Y gnd NAND3X1_224/A vdd OAI21X1
XNOR2X1_247 BUFX2_201/A XOR2X1_204/Y gnd NOR2X1_247/Y vdd NOR2X1
XNAND2X1_328 INVX1_192/A NAND2X1_328/B gnd NOR3X1_57/B vdd NAND2X1
XINVX2_35 INVX2_35/A gnd INVX2_35/Y vdd INVX2
XCLKBUF1_38 BUFX4_6/Y gnd CLKBUF1_38/Y vdd CLKBUF1
XNAND3X1_160 INVX1_103/Y NAND3X1_162/B OR2X2_69/Y gnd NAND3X1_160/Y vdd NAND3X1
XBUFX2_161 BUFX2_161/A gnd BUFX2_161/Y vdd BUFX2
XINVX1_576 INVX1_576/A gnd INVX1_576/Y vdd INVX1
XXNOR2X1_5 XNOR2X1_5/A INVX2_11/Y gnd OR2X2_20/A vdd XNOR2X1
XFILL_6_0_0 gnd vdd FILL
XFILL_24_1_1 gnd vdd FILL
XNOR2X1_14 OAI22X1_8/Y NOR2X1_14/B gnd NOR2X1_14/Y vdd NOR2X1
XXNOR2X1_199 XNOR2X1_199/A XNOR2X1_199/B gnd INVX1_433/A vdd XNOR2X1
XFILL_4_2_1 gnd vdd FILL
XNAND2X1_292 gnd OR2X2_115/B gnd NAND3X1_262/B vdd NAND2X1
XNOR2X1_211 BUFX2_185/A NOR2X1_211/B gnd NOR2X1_211/Y vdd NOR2X1
XOAI21X1_178 AND2X2_62/Y NOR3X1_45/B INVX1_121/Y gnd OAI21X1_178/Y vdd OAI21X1
XINVX4_2 INVX4_2/A gnd INVX4_2/Y vdd INVX4
XNOR3X1_91 OR2X2_129/Y NOR3X1_91/B NOR3X1_91/C gnd NOR3X1_91/Y vdd NOR3X1
XBUFX2_125 gnd gnd BUFX2_125/Y vdd BUFX2
XNAND3X1_124 INVX1_81/Y NAND3X1_126/B OR2X2_53/Y gnd NAND3X1_124/Y vdd NAND3X1
XINVX1_540 INVX1_540/A gnd INVX1_540/Y vdd INVX1
XDFFPOSX1_358 INVX1_443/A CLKBUF1_13/Y OR2X2_153/Y gnd vdd DFFPOSX1
XBUFX4_7 clk gnd BUFX4_7/Y vdd BUFX4
XXNOR2X1_163 XNOR2X1_163/A XNOR2X1_163/B gnd INVX1_262/A vdd XNOR2X1
XOAI21X1_142 OAI21X1_142/A OAI21X1_141/Y INVX1_95/Y gnd NAND3X1_148/C vdd OAI21X1
XXNOR2X1_85 gnd XOR2X1_82/Y gnd XNOR2X1_85/Y vdd XNOR2X1
XFILL_13_9_0 gnd vdd FILL
XNAND2X1_256 INVX2_48/Y OAI21X1_221/Y gnd XNOR2X1_116/A vdd NAND2X1
XNOR2X1_175 NOR2X1_175/A INVX1_181/Y gnd NOR2X1_175/Y vdd NOR2X1
XNOR3X1_55 NOR3X1_55/A NOR3X1_55/B NOR3X1_55/C gnd NOR3X1_55/Y vdd NOR3X1
XDFFPOSX1_322 INVX1_358/A CLKBUF1_45/Y INVX1_568/Y gnd vdd DFFPOSX1
XXNOR2X1_127 BUFX2_165/A XOR2X1_128/Y gnd OR2X2_111/A vdd XNOR2X1
XINVX1_504 INVX1_504/A gnd INVX1_504/Y vdd INVX1
XXNOR2X1_49 gnd XOR2X1_42/Y gnd AOI21X1_81/B vdd XNOR2X1
XOAI21X1_106 XNOR2X1_53/A AOI21X1_82/C NOR2X1_75/Y gnd NOR2X1_76/B vdd OAI21X1
XNOR2X1_139 gnd OR2X2_98/B gnd NOR3X1_50/B vdd NOR2X1
XFILL_23_4_0 gnd vdd FILL
XFILL_3_5_0 gnd vdd FILL
XNAND2X1_220 OR2X2_85/A OR2X2_85/B gnd NAND2X1_220/Y vdd NAND2X1
XFILL_21_6_1 gnd vdd FILL
XNOR3X1_19 BUFX4_25/Y MUX2X1_19/Y BUFX4_21/Y gnd NOR3X1_19/Y vdd NOR3X1
XFILL_1_7_1 gnd vdd FILL
XOAI21X1_647 AND2X2_198/Y NOR2X1_451/Y INVX1_594/Y gnd NAND3X1_546/A vdd OAI21X1
XDFFPOSX1_286 INVX1_272/A CLKBUF1_23/Y OR2X2_138/A gnd vdd DFFPOSX1
XINVX1_468 INVX1_468/A gnd INVX1_468/Y vdd INVX1
XXNOR2X1_13 gnd XOR2X1_2/Y gnd XNOR2X1_14/A vdd XNOR2X1
XXOR2X1_283 XOR2X1_283/A BUFX2_231/A gnd INVX1_461/A vdd XOR2X1
XNOR2X1_103 NOR2X1_103/A NOR3X1_42/Y gnd NOR2X1_103/Y vdd NOR2X1
XNAND2X1_184 OAI21X1_156/Y OR2X2_72/B gnd OR2X2_70/A vdd NAND2X1
XFILL_31_1_1 gnd vdd FILL
XDFFPOSX1_250 INVX1_187/A CLKBUF1_11/Y OR2X2_142/A gnd vdd DFFPOSX1
XOR2X2_71 OR2X2_71/A OR2X2_71/B gnd OR2X2_71/Y vdd OR2X2
XAOI21X1_82 AOI21X1_82/A AOI21X1_82/B AOI21X1_82/C gnd AOI21X1_82/Y vdd AOI21X1
XOAI21X1_611 AND2X2_176/Y NOR2X1_408/Y OAI21X1_611/C gnd NOR2X1_426/B vdd OAI21X1
XXOR2X1_247 XOR2X1_247/A BUFX2_215/A gnd INVX1_385/A vdd XOR2X1
XINVX1_432 INVX1_432/A gnd INVX1_432/Y vdd INVX1
XBUFX2_85 gnd gnd BUFX2_85/Y vdd BUFX2
XNAND2X1_148 NAND2X1_147/Y OR2X2_55/Y gnd OR2X2_56/A vdd NAND2X1
XAOI21X1_384 AOI21X1_384/A OR2X2_140/Y NAND3X1_508/Y gnd INVX1_566/A vdd AOI21X1
XAOI21X1_46 AOI21X1_44/Y AOI21X1_46/B AOI21X1_46/C gnd AOI21X1_46/Y vdd AOI21X1
XOR2X2_35 gnd OR2X2_35/B gnd OR2X2_35/Y vdd OR2X2
XDFFPOSX1_214 INVX1_135/A CLKBUF1_10/Y INVX1_572/A gnd vdd DFFPOSX1
XINVX1_396 INVX1_396/A gnd INVX1_396/Y vdd INVX1
XOAI21X1_575 NOR2X1_389/Y AND2X2_162/B BUFX4_31/Y gnd AOI21X1_330/C vdd OAI21X1
XNAND2X1_689 NAND3X1_526/B INVX1_566/A gnd NAND2X1_689/Y vdd NAND2X1
XFILL_20_9_0 gnd vdd FILL
XXOR2X1_211 XOR2X1_211/A INVX1_289/A gnd INVX1_309/A vdd XOR2X1
XBUFX2_49 gnd gnd BUFX2_49/Y vdd BUFX2
XNAND2X1_112 NAND2X1_112/A OR2X2_40/Y gnd INVX1_62/A vdd NAND2X1
XAOI21X1_348 INVX2_81/Y AOI21X1_348/B OAI21X1_588/Y gnd AOI21X1_348/Y vdd AOI21X1
XOAI21X1_94 NOR2X1_73/B NOR2X1_73/A NOR3X1_35/Y gnd OAI21X1_94/Y vdd OAI21X1
XNAND3X1_521 INVX1_560/A XNOR2X1_236/Y NAND3X1_521/C gnd NAND3X1_521/Y vdd NAND3X1
XDFFPOSX1_178 INVX2_32/A CLKBUF1_40/Y bloque_bytes[24] gnd vdd DFFPOSX1
XINVX1_360 INVX1_360/A gnd INVX1_360/Y vdd INVX1
XAOI21X1_10 AOI21X1_9/Y AOI21X1_5/Y MUX2X1_9/S gnd BUFX4_18/A vdd AOI21X1
XFILL_30_4_0 gnd vdd FILL
XOAI21X1_539 BUFX2_232/A NOR2X1_342/B INVX1_444/Y gnd OAI21X1_539/Y vdd OAI21X1
XXOR2X1_175 XOR2X1_175/A BUFX2_179/A gnd INVX1_233/A vdd XOR2X1
XNAND2X1_653 XNOR2X1_211/Y NAND2X1_653/B gnd NAND2X1_653/Y vdd NAND2X1
XBUFX2_13 BUFX2_13/A gnd hash[12] vdd BUFX2
XFILL_28_6_1 gnd vdd FILL
XNAND2X1_73 OR2X2_24/B OR2X2_24/A gnd NAND2X1_74/A vdd NAND2X1
XFILL_8_7_1 gnd vdd FILL
XNAND3X1_485 INVX1_459/A OAI21X1_555/Y NAND3X1_480/Y gnd NAND2X1_607/A vdd NAND3X1
XAOI21X1_312 AOI21X1_312/A AOI21X1_312/B AOI21X1_312/C gnd OAI21X1_543/A vdd AOI21X1
XOAI21X1_58 NOR2X1_47/A INVX1_42/Y INVX1_43/Y gnd OAI21X1_58/Y vdd OAI21X1
XDFFPOSX1_142 INVX1_36/A CLKBUF1_7/Y bloque_bytes[68] gnd vdd DFFPOSX1
XDFFPOSX1_76 AND2X2_166/B CLKBUF1_30/Y DFFPOSX1_76/D gnd vdd DFFPOSX1
XXOR2X1_139 XOR2X1_139/A BUFX2_166/A gnd XOR2X1_139/Y vdd XOR2X1
XINVX1_324 INVX1_324/A gnd INVX1_324/Y vdd INVX1
XOAI21X1_503 gnd XOR2X1_254/Y INVX1_398/Y gnd OAI21X1_503/Y vdd OAI21X1
XNAND2X1_617 AND2X2_161/B INVX1_476/A gnd NOR2X1_398/A vdd NAND2X1
XOAI21X1_22 INVX2_13/Y AND2X2_6/B OR2X2_6/Y gnd OAI21X1_23/B vdd OAI21X1
XNAND2X1_37 INVX2_13/A AND2X2_6/Y gnd OAI21X1_21/B vdd NAND2X1
XNAND3X1_449 INVX2_71/A NAND3X1_449/B NAND2X1_554/Y gnd NOR3X1_81/A vdd NAND3X1
XAOI21X1_276 NAND3X1_420/B NAND3X1_420/C INVX1_364/A gnd NOR2X1_292/A vdd AOI21X1
XDFFPOSX1_40 INVX1_575/A CLKBUF1_15/Y NOR2X1_365/Y gnd vdd DFFPOSX1
XINVX1_288 INVX1_288/A gnd INVX1_288/Y vdd INVX1
XOAI21X1_467 OAI21X1_467/A INVX1_375/A INVX1_374/Y gnd AND2X2_137/A vdd OAI21X1
XDFFPOSX1_106 INVX1_10/A CLKBUF1_42/Y INVX1_584/Y gnd vdd DFFPOSX1
XXOR2X1_103 OR2X2_93/A gnd gnd OR2X2_89/B vdd XOR2X1
XXOR2X1_83 OR2X2_77/A gnd gnd OR2X2_73/B vdd XOR2X1
XNAND2X1_581 NAND3X1_469/Y NAND3X1_470/Y gnd XOR2X1_287/B vdd NAND2X1
XAOI21X1_240 AOI21X1_240/A AOI21X1_240/B NAND2X1_412/Y gnd OAI21X1_372/A vdd AOI21X1
XFILL_27_9_0 gnd vdd FILL
XAOI22X1_15 INVX1_333/A AOI22X1_15/B AOI22X1_15/C INVX1_331/A gnd INVX1_337/A vdd
+ AOI22X1
XNAND3X1_413 INVX1_364/A NAND2X1_501/Y INVX1_363/Y gnd INVX1_370/A vdd NAND3X1
XAND2X2_9 gnd AND2X2_9/B gnd AND2X2_9/Y vdd AND2X2
XINVX1_252 INVX1_252/A gnd INVX1_252/Y vdd INVX1
XAND2X2_183 INVX1_538/A AND2X2_183/B gnd INVX1_550/A vdd AND2X2
XOAI21X1_431 OAI21X1_431/A INVX1_335/A INVX1_338/A gnd OAI21X1_431/Y vdd OAI21X1
XXOR2X1_47 XOR2X1_47/A OR2X2_37/A gnd OR2X2_45/B vdd XOR2X1
XNAND3X1_78 NAND3X1_77/Y OAI21X1_76/Y NAND3X1_78/C gnd OAI21X1_85/B vdd NAND3X1
XOR2X2_130 OR2X2_130/A INVX2_81/Y gnd OR2X2_130/Y vdd OR2X2
XNAND2X1_545 XOR2X1_269/B NOR2X1_316/Y gnd AOI21X1_296/C vdd NAND2X1
XAOI21X1_204 AOI21X1_204/A AOI21X1_204/B INVX1_193/A gnd NOR2X1_184/A vdd AOI21X1
XFILL_35_6_1 gnd vdd FILL
XNAND3X1_377 INVX1_312/A NAND3X1_375/Y INVX1_307/Y gnd AOI22X1_14/C vdd NAND3X1
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XXOR2X1_11 vdd XOR2X1_11/B gnd XOR2X1_11/Y vdd XOR2X1
XNAND3X1_42 NAND3X1_42/A NAND3X1_42/B NAND3X1_42/C gnd OAI21X1_46/B vdd NAND3X1
XINVX1_216 INVX1_216/A gnd INVX1_216/Y vdd INVX1
XNOR2X1_428 bloque_bytes[13] NOR2X1_428/B gnd INVX1_555/A vdd NOR2X1
XAND2X2_147 NOR2X1_323/Y INVX1_416/Y gnd NOR3X1_82/C vdd AND2X2
XOAI21X1_395 gnd XOR2X1_208/Y INVX1_302/A gnd INVX2_65/A vdd OAI21X1
XNAND2X1_509 OAI21X1_466/Y NAND2X1_508/Y gnd NOR2X1_296/B vdd NAND2X1
XNAND3X1_341 INVX1_247/Y NAND3X1_334/Y NOR3X1_64/Y gnd AOI21X1_232/B vdd NAND3X1
XAOI21X1_168 AOI21X1_168/A AOI21X1_168/B NAND3X1_242/C gnd NOR2X1_151/A vdd AOI21X1
XCLKBUF1_1 BUFX4_6/Y gnd CLKBUF1_1/Y vdd CLKBUF1
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XINVX1_180 INVX1_180/A gnd INVX1_180/Y vdd INVX1
XAND2X2_111 AND2X2_111/A INVX1_245/Y gnd NOR3X1_64/C vdd AND2X2
XOAI21X1_359 gnd NOR2X1_228/B INVX1_265/A gnd INVX1_268/A vdd OAI21X1
XFILL_11_2_0 gnd vdd FILL
XNOR2X1_392 NOR2X1_391/Y NOR2X1_392/B gnd NOR2X1_392/Y vdd NOR2X1
XNAND2X1_473 NAND2X1_473/A INVX1_335/Y gnd INVX1_336/A vdd NAND2X1
XAND2X2_84 AND2X2_84/A AND2X2_84/B gnd AND2X2_84/Y vdd AND2X2
XAOI21X1_132 OAI21X1_183/Y NAND3X1_190/Y NAND3X1_187/Y gnd NOR2X1_121/A vdd AOI21X1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XNAND3X1_305 INVX1_202/Y INVX1_205/Y AND2X2_101/A gnd NAND2X1_342/B vdd NAND3X1
XOAI21X1_323 NOR3X1_62/A NOR3X1_62/C INVX2_61/A gnd NOR2X1_205/A vdd OAI21X1
XINVX1_144 INVX1_144/A gnd INVX1_144/Y vdd INVX1
XFILL_34_9_0 gnd vdd FILL
XNOR2X1_356 INVX1_466/Y NOR2X1_356/B gnd INVX1_468/A vdd NOR2X1
XNAND2X1_437 NAND2X1_437/A NAND3X1_370/Y gnd XOR2X1_223/A vdd NAND2X1
XBUFX2_270 XOR2X1_99/B gnd BUFX2_270/Y vdd BUFX2
XNAND3X1_269 NAND3X1_267/A NAND3X1_269/B NAND3X1_269/C gnd AOI21X1_185/A vdd NAND3X1
XAND2X2_48 AND2X2_48/A AND2X2_48/B gnd AND2X2_48/Y vdd AND2X2
XINVX1_108 OR2X2_72/Y gnd INVX1_108/Y vdd INVX1
XBUFX4_33 reset gnd BUFX4_33/Y vdd BUFX4
XOAI21X1_287 gnd NOR2X1_183/B INVX1_191/A gnd INVX1_193/A vdd OAI21X1
XNAND2X1_401 OAI21X1_356/Y NAND3X1_345/B gnd BUFX2_203/A vdd NAND2X1
XAOI22X1_6 INVX2_6/Y INVX2_10/A INVX1_9/A INVX2_7/Y gnd AOI22X1_6/Y vdd AOI22X1
XNOR2X1_320 INVX1_409/Y NOR2X1_320/B gnd INVX1_411/A vdd NOR2X1
XAND2X2_12 AND2X2_12/A AND2X2_12/B gnd AND2X2_12/Y vdd AND2X2
XFILL_6_1 gnd vdd FILL
XNAND3X1_233 NAND3X1_233/A NAND3X1_233/B NAND3X1_233/C gnd AOI21X1_161/A vdd NAND3X1
XBUFX2_234 BUFX2_234/A gnd BUFX2_234/Y vdd BUFX2
XNOR2X1_87 NOR2X1_87/A NOR2X1_87/B gnd NOR2X1_87/Y vdd NOR2X1
XOAI21X1_251 AND2X2_88/Y NOR2X1_160/Y INVX1_167/Y gnd AOI21X1_180/A vdd OAI21X1
XNAND2X1_365 INVX1_227/Y NOR2X1_204/Y gnd NAND2X1_365/Y vdd NAND2X1
XNOR2X1_284 INVX1_352/Y NOR2X1_284/B gnd INVX1_354/A vdd NOR2X1
XINVX2_72 INVX2_72/A gnd INVX2_72/Y vdd INVX2
XFILL_18_2_0 gnd vdd FILL
XNAND3X1_197 NAND3X1_197/A OAI21X1_189/Y NAND3X1_196/Y gnd AOI21X1_137/A vdd NAND3X1
XNOR2X1_51 NOR2X1_51/A INVX2_21/A gnd XOR2X1_40/B vdd NOR2X1
XBUFX2_198 XOR2X1_15/A gnd BUFX2_198/Y vdd BUFX2
XFILL_16_4_1 gnd vdd FILL
XXNOR2X1_236 XNOR2X1_236/A NOR2X1_411/A gnd XNOR2X1_236/Y vdd XNOR2X1
XINVX2_36 INVX2_36/A gnd INVX2_36/Y vdd INVX2
XOAI21X1_215 NOR3X1_50/Y NOR2X1_143/A NAND2X1_250/B gnd NAND2X1_253/B vdd OAI21X1
XNOR2X1_248 INVX1_295/Y NOR2X1_248/B gnd INVX1_297/A vdd NOR2X1
XNAND2X1_329 INVX1_191/A NOR2X1_183/Y gnd NAND2X1_329/Y vdd NAND2X1
XNAND3X1_161 NAND3X1_161/A OAI21X1_155/Y NAND3X1_160/Y gnd NAND3X1_161/Y vdd NAND3X1
XBUFX2_162 BUFX2_162/A gnd BUFX2_162/Y vdd BUFX2
XINVX1_577 INVX1_577/A gnd INVX1_577/Y vdd INVX1
XCLKBUF1_39 BUFX4_5/Y gnd CLKBUF1_39/Y vdd CLKBUF1
XXNOR2X1_6 XNOR2X1_6/A XNOR2X1_6/B gnd OR2X2_21/A vdd XNOR2X1
XFILL_6_0_1 gnd vdd FILL
XOAI21X1_179 NOR3X1_46/Y NOR2X1_123/A NOR3X1_45/Y gnd OAI21X1_179/Y vdd OAI21X1
XNOR2X1_15 NOR2X1_15/A NOR2X1_15/B gnd NAND3X1_4/C vdd NOR2X1
XXNOR2X1_200 NOR2X1_338/A NAND2X1_578/Y gnd BUFX2_246/A vdd XNOR2X1
XNOR2X1_212 INVX1_238/Y NOR2X1_212/B gnd INVX1_240/A vdd NOR2X1
XNAND2X1_293 AND2X2_89/A AND2X2_89/B gnd NAND3X1_264/B vdd NAND2X1
XNOR3X1_92 NOR3X1_92/A INVX1_492/A NOR3X1_95/C gnd NOR3X1_93/C vdd NOR3X1
XDFFPOSX1_359 INVX1_444/A CLKBUF1_13/Y NAND2X1_692/Y gnd vdd DFFPOSX1
XNAND3X1_125 NAND3X1_123/A OAI21X1_121/Y NAND3X1_124/Y gnd AOI21X1_89/A vdd NAND3X1
XBUFX2_126 gnd gnd BUFX2_126/Y vdd BUFX2
XINVX1_541 INVX1_541/A gnd INVX1_541/Y vdd INVX1
XBUFX4_8 BUFX4_8/A gnd BUFX4_8/Y vdd BUFX4
XXNOR2X1_164 NOR2X1_230/A NAND2X1_407/Y gnd BUFX2_206/A vdd XNOR2X1
XFILL_15_7_0 gnd vdd FILL
XOAI21X1_143 NOR2X1_97/A INVX1_97/Y INVX1_98/Y gnd OAI21X1_143/Y vdd OAI21X1
XXNOR2X1_86 XNOR2X1_85/Y INVX2_38/Y gnd OR2X2_92/A vdd XNOR2X1
XFILL_13_9_1 gnd vdd FILL
XNOR2X1_176 INVX1_183/Y NOR2X1_176/B gnd NOR2X1_177/B vdd NOR2X1
XNAND2X1_257 AND2X2_78/B AND2X2_78/A gnd OAI21X1_222/B vdd NAND2X1
XINVX1_505 bloque_bytes[39] gnd INVX1_505/Y vdd INVX1
XNOR3X1_56 NOR3X1_56/A NOR3X1_56/B AND2X2_93/Y gnd NOR3X1_56/Y vdd NOR3X1
XDFFPOSX1_323 INVX1_359/A CLKBUF1_8/Y INVX1_569/Y gnd vdd DFFPOSX1
XXNOR2X1_128 XOR2X1_141/Y XOR2X1_129/Y gnd XNOR2X1_129/A vdd XNOR2X1
XOAI21X1_107 INVX2_28/Y AND2X2_36/B OR2X2_46/Y gnd OAI21X1_107/Y vdd OAI21X1
XXNOR2X1_50 AOI21X1_81/B INVX2_26/Y gnd OR2X2_60/A vdd XNOR2X1
XNOR2X1_140 gnd OR2X2_99/B gnd NOR2X1_140/Y vdd NOR2X1
XFILL_23_4_1 gnd vdd FILL
XFILL_25_2_0 gnd vdd FILL
XFILL_3_5_1 gnd vdd FILL
XFILL_5_3_0 gnd vdd FILL
XNAND2X1_221 AOI21X1_137/A AOI21X1_137/B gnd INVX2_43/A vdd NAND2X1
XNOR3X1_20 NOR3X1_9/A MUX2X1_20/Y NOR3X1_9/C gnd NOR3X1_20/Y vdd NOR3X1
XOAI21X1_648 XNOR2X1_255/A OAI21X1_648/B NOR2X1_452/Y gnd NOR2X1_453/B vdd OAI21X1
XDFFPOSX1_287 INVX1_273/A CLKBUF1_2/Y NOR2X1_428/B gnd vdd DFFPOSX1
XINVX1_469 INVX1_469/A gnd INVX1_469/Y vdd INVX1
XXNOR2X1_14 XNOR2X1_14/A INVX2_14/Y gnd OR2X2_28/A vdd XNOR2X1
XXOR2X1_284 XOR2X1_278/Y BUFX2_232/A gnd XOR2X1_284/Y vdd XOR2X1
XNOR2X1_104 OR2X2_69/A OR2X2_69/B gnd NOR2X1_104/Y vdd NOR2X1
XNAND2X1_185 OR2X2_71/B OR2X2_71/A gnd NAND2X1_185/Y vdd NAND2X1
XAOI21X1_83 AOI21X1_83/A OR2X2_50/Y INVX1_78/A gnd NOR2X1_83/A vdd AOI21X1
XDFFPOSX1_251 INVX1_188/A CLKBUF1_31/Y OR2X2_143/A gnd vdd DFFPOSX1
XOR2X2_72 OR2X2_72/A OR2X2_72/B gnd OR2X2_72/Y vdd OR2X2
XOAI21X1_612 INVX1_536/Y bloque_bytes[26] INVX1_537/Y gnd AOI21X1_376/C vdd OAI21X1
XXOR2X1_248 XOR2X1_242/Y BUFX2_216/A gnd NOR2X1_306/B vdd XOR2X1
XINVX1_433 INVX1_433/A gnd INVX1_433/Y vdd INVX1
XBUFX2_86 gnd gnd BUFX2_86/Y vdd BUFX2
XNAND2X1_149 OR2X2_56/B OR2X2_56/A gnd NAND2X1_149/Y vdd NAND2X1
XAOI21X1_385 AOI21X1_385/A OR2X2_141/Y AOI21X1_385/C gnd INVX1_567/A vdd AOI21X1
XAOI21X1_47 NAND2X1_80/Y OR2X2_26/Y INVX1_45/A gnd NOR2X1_53/A vdd AOI21X1
XOR2X2_36 OR2X2_36/A OR2X2_36/B gnd OR2X2_36/Y vdd OR2X2
XOAI21X1_576 INVX2_83/A INVX2_75/A BUFX4_32/Y gnd OAI21X1_576/Y vdd OAI21X1
XDFFPOSX1_215 INVX1_136/A CLKBUF1_50/Y INVX2_88/A gnd vdd DFFPOSX1
XFILL_22_7_0 gnd vdd FILL
XINVX1_397 INVX1_397/A gnd INVX1_397/Y vdd INVX1
XFILL_2_8_0 gnd vdd FILL
XFILL_20_9_1 gnd vdd FILL
XNAND2X1_690 INVX1_543/Y INVX1_567/A gnd NAND2X1_690/Y vdd NAND2X1
XXOR2X1_212 XOR2X1_206/Y BUFX2_200/A gnd XOR2X1_212/Y vdd XOR2X1
XBUFX2_50 gnd gnd BUFX2_50/Y vdd BUFX2
XNAND2X1_113 INVX2_25/A AND2X2_30/Y gnd OAI21X1_89/B vdd NAND2X1
XAOI21X1_349 NOR2X1_407/Y NOR3X1_90/Y INVX1_485/A gnd NOR3X1_96/B vdd AOI21X1
XOAI21X1_95 NOR3X1_36/C NOR3X1_36/B INVX1_67/Y gnd NAND3X1_99/B vdd OAI21X1
XNAND3X1_522 INVX1_537/Y NAND2X1_659/B INVX1_561/A gnd NAND3X1_522/Y vdd NAND3X1
XDFFPOSX1_179 INVX1_88/A CLKBUF1_13/Y bloque_bytes[25] gnd vdd DFFPOSX1
XFILL_32_2_0 gnd vdd FILL
XAOI21X1_11 NAND3X1_7/B OR2X2_2/Y INVX1_12/A gnd OAI21X1_9/B vdd AOI21X1
XINVX1_361 INVX1_361/A gnd INVX1_361/Y vdd INVX1
XFILL_30_4_1 gnd vdd FILL
XOAI21X1_540 BUFX2_232/A NOR2X1_342/B INVX1_444/A gnd AOI22X1_21/B vdd OAI21X1
XXOR2X1_176 XOR2X1_176/A BUFX2_180/A gnd NOR2X1_210/B vdd XOR2X1
XNAND2X1_654 NAND2X1_654/A AOI21X1_374/Y gnd XNOR2X1_238/A vdd NAND2X1
XBUFX2_14 BUFX2_14/A gnd hash[13] vdd BUFX2
XNAND2X1_74 NAND2X1_74/A OR2X2_24/Y gnd INVX1_40/A vdd NAND2X1
XNAND3X1_486 INVX1_470/Y INVX1_469/A AOI21X1_322/B gnd AND2X2_157/B vdd NAND3X1
XAOI21X1_313 NAND3X1_469/Y NAND3X1_470/Y NAND2X1_588/Y gnd AOI21X1_313/Y vdd AOI21X1
XDFFPOSX1_143 INVX1_37/A CLKBUF1_7/Y bloque_bytes[69] gnd vdd DFFPOSX1
XOAI21X1_59 NOR3X1_31/C NOR3X1_31/B INVX1_44/Y gnd NAND3X1_60/B vdd OAI21X1
XDFFPOSX1_77 INVX1_479/A CLKBUF1_30/Y DFFPOSX1_77/D gnd vdd DFFPOSX1
XINVX1_325 INVX1_325/A gnd INVX1_325/Y vdd INVX1
XNAND2X1_618 AND2X2_163/B NOR2X1_390/Y gnd NOR2X1_393/B vdd NAND2X1
XXOR2X1_140 XOR2X1_140/A XOR2X1_140/B gnd BUFX2_174/A vdd XOR2X1
XOAI21X1_504 BUFX2_225/A NOR2X1_319/B INVX1_410/A gnd OAI21X1_504/Y vdd OAI21X1
XNAND2X1_38 NAND2X1_38/A OAI21X1_24/Y gnd XOR2X1_19/A vdd NAND2X1
XOAI21X1_23 OAI21X1_23/A OAI21X1_23/B INVX1_18/Y gnd NAND3X1_22/C vdd OAI21X1
XDFFPOSX1_41 INVX1_543/A CLKBUF1_3/Y NOR2X1_366/Y gnd vdd DFFPOSX1
XNAND3X1_450 INVX1_420/A NAND2X1_555/Y INVX2_71/Y gnd OAI21X1_512/C vdd NAND3X1
XAOI21X1_277 INVX1_364/A NAND2X1_501/Y INVX1_363/Y gnd NOR3X1_75/C vdd AOI21X1
XFILL_19_1 gnd vdd FILL
XINVX1_289 INVX1_289/A gnd INVX1_289/Y vdd INVX1
XOAI21X1_468 NOR2X1_293/A NOR3X1_75/Y AOI21X1_281/Y gnd AOI21X1_282/B vdd OAI21X1
XDFFPOSX1_107 MUX2X1_18/B CLKBUF1_42/Y NOR2X1_440/Y gnd vdd DFFPOSX1
XXOR2X1_104 BUFX2_157/A gnd gnd OR2X2_90/B vdd XOR2X1
XNAND2X1_582 INVX1_436/A NOR2X1_336/Y gnd AOI21X1_310/B vdd NAND2X1
XXOR2X1_84 XOR2X1_98/B gnd gnd OR2X2_74/B vdd XOR2X1
XFILL_9_8_0 gnd vdd FILL
XAOI21X1_241 AOI21X1_241/A NAND2X1_410/B NAND2X1_417/Y gnd OAI21X1_373/C vdd AOI21X1
XFILL_27_9_1 gnd vdd FILL
XAOI22X1_16 INVX1_352/A AOI22X1_16/B AOI22X1_16/C INVX1_350/A gnd INVX1_356/A vdd
+ AOI22X1
XFILL_29_7_0 gnd vdd FILL
XNAND3X1_414 INVX1_365/Y INVX1_366/Y INVX1_367/Y gnd AOI21X1_275/B vdd NAND3X1
XXOR2X1_48 XOR2X1_48/A BUFX2_249/A gnd XOR2X1_48/Y vdd XOR2X1
XINVX1_253 INVX1_253/A gnd INVX1_253/Y vdd INVX1
XAND2X2_184 INVX1_539/A AND2X2_184/B gnd INVX1_551/A vdd AND2X2
XOAI21X1_432 gnd XOR2X1_225/Y INVX1_339/A gnd OAI21X1_432/Y vdd OAI21X1
XNAND3X1_79 INVX1_56/A NAND2X1_99/Y OR2X2_34/Y gnd NAND3X1_79/Y vdd NAND3X1
XOR2X2_131 bloque_bytes[72] bloque_bytes[32] gnd OR2X2_131/Y vdd OR2X2
XNAND2X1_546 INVX1_410/Y NOR2X1_319/Y gnd NAND2X1_546/Y vdd NAND2X1
XAOI21X1_205 INVX1_193/A NAND3X1_296/B INVX1_192/Y gnd NOR3X1_57/C vdd AOI21X1
XNAND3X1_378 INVX1_312/A NAND3X1_378/B NAND3X1_378/C gnd AOI21X1_257/A vdd NAND3X1
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XOAI21X1_396 NOR3X1_70/C INVX2_65/Y NOR3X1_70/A gnd AND2X2_124/A vdd OAI21X1
XMUX2X1_1 BUFX2_1/A MUX2X1_1/B MUX2X1_8/S gnd MUX2X1_1/Y vdd MUX2X1
XXOR2X1_12 OR2X2_20/A gnd gnd XOR2X1_12/Y vdd XOR2X1
XNAND3X1_43 INVX1_34/A NAND2X1_61/Y OR2X2_18/Y gnd AOI21X1_36/C vdd NAND3X1
XNOR2X1_429 bloque_bytes[14] NOR2X1_429/B gnd INVX1_556/A vdd NOR2X1
XAND2X2_148 AND2X2_148/A NOR3X1_81/A gnd BUFX2_236/A vdd AND2X2
XNAND2X1_510 INVX1_371/Y NOR2X1_296/B gnd NAND2X1_510/Y vdd NAND2X1
XAOI21X1_169 AOI21X1_169/A AOI21X1_169/B NOR3X1_52/Y gnd INVX2_51/A vdd AOI21X1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XNAND3X1_342 INVX1_250/A AOI21X1_228/A AOI21X1_228/B gnd NAND3X1_342/Y vdd NAND3X1
XFILL_11_2_1 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XINVX1_181 INVX1_181/A gnd INVX1_181/Y vdd INVX1
XAND2X2_112 AND2X2_112/A NOR3X1_63/A gnd BUFX2_200/A vdd AND2X2
XCLKBUF1_2 BUFX4_5/Y gnd CLKBUF1_2/Y vdd CLKBUF1
XOAI21X1_360 NOR3X1_65/A NOR3X1_65/B OAI21X1_366/B gnd NOR2X1_230/A vdd OAI21X1
XNOR2X1_393 INVX1_477/Y NOR2X1_393/B gnd NOR3X1_87/C vdd NOR2X1
XNAND2X1_474 NAND2X1_474/A AOI22X1_15/C gnd NAND2X1_474/Y vdd NAND2X1
XAOI21X1_133 AOI21X1_133/A AOI21X1_133/B NOR3X1_46/Y gnd INVX2_42/A vdd AOI21X1
XNAND3X1_306 INVX2_60/A NAND3X1_306/B NAND3X1_306/C gnd NOR3X1_59/A vdd NAND3X1
XAND2X2_85 BUFX2_164/A OR2X2_109/B gnd AND2X2_85/Y vdd AND2X2
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XFILL_36_7_0 gnd vdd FILL
XOAI21X1_324 gnd NOR2X1_207/B INVX1_229/Y gnd OAI21X1_324/Y vdd OAI21X1
XINVX1_145 INVX1_145/A gnd INVX1_145/Y vdd INVX1
XNOR2X1_357 BUFX2_238/A NOR2X1_357/B gnd NOR2X1_357/Y vdd NOR2X1
XFILL_34_9_1 gnd vdd FILL
XNAND2X1_438 INVX1_301/Y AND2X2_122/A gnd NAND2X1_439/B vdd NAND2X1
XBUFX2_271 OR2X2_84/A gnd BUFX2_271/Y vdd BUFX2
XNAND3X1_270 INVX1_169/A NAND3X1_270/B OR2X2_117/Y gnd OR2X2_120/B vdd NAND3X1
XAND2X2_49 OR2X2_61/A OR2X2_61/B gnd AND2X2_49/Y vdd AND2X2
XINVX1_109 INVX1_109/A gnd INVX1_109/Y vdd INVX1
XOAI21X1_288 INVX1_194/A INVX1_195/A INVX1_196/A gnd AOI22X1_8/D vdd OAI21X1
XNAND2X1_402 INVX1_264/Y AND2X2_115/A gnd NAND3X1_345/C vdd NAND2X1
XAOI22X1_7 OAI22X1_6/Y NAND3X1_2/A NOR2X1_13/Y AOI22X1_7/D gnd AOI22X1_7/Y vdd AOI22X1
XNOR2X1_321 BUFX2_226/A XOR2X1_259/Y gnd NOR2X1_321/Y vdd NOR2X1
XAND2X2_13 XOR2X1_3/A OR2X2_13/B gnd AND2X2_13/Y vdd AND2X2
XFILL_10_5_0 gnd vdd FILL
XFILL_6_2 gnd vdd FILL
XNAND3X1_234 INVX1_147/A NAND3X1_234/B OR2X2_101/Y gnd OR2X2_104/B vdd NAND3X1
XNOR2X1_88 gnd OR2X2_57/B gnd NOR2X1_88/Y vdd NOR2X1
XBUFX2_235 INVX1_460/A gnd BUFX2_235/Y vdd BUFX2
XOAI21X1_252 AND2X2_88/Y NOR2X1_160/Y INVX1_167/A gnd OAI21X1_252/Y vdd OAI21X1
XNOR2X1_285 BUFX2_214/A XOR2X1_232/Y gnd NOR2X1_285/Y vdd NOR2X1
XNAND2X1_366 INVX1_230/A NAND2X1_365/Y gnd NOR3X1_61/B vdd NAND2X1
XFILL_20_0_0 gnd vdd FILL
XINVX2_73 INVX2_73/A gnd INVX2_73/Y vdd INVX2
XFILL_0_1_0 gnd vdd FILL
XNAND3X1_198 INVX1_125/A NAND2X1_220/Y OR2X2_85/Y gnd OR2X2_88/B vdd NAND3X1
XFILL_18_2_1 gnd vdd FILL
XBUFX2_199 INVX1_289/A gnd BUFX2_199/Y vdd BUFX2
XNOR2X1_52 OR2X2_28/A OR2X2_28/B gnd NOR2X1_52/Y vdd NOR2X1
XXNOR2X1_237 NAND2X1_653/Y AOI21X1_353/C gnd NAND3X1_523/B vdd XNOR2X1
XINVX2_37 INVX2_37/A gnd INVX2_37/Y vdd INVX2
XNAND2X1_330 INVX1_191/Y NOR2X1_183/Y gnd NAND3X1_296/B vdd NAND2X1
XOAI21X1_216 OAI21X1_216/A XNOR2X1_115/B INVX1_151/A gnd XOR2X1_130/A vdd OAI21X1
XNOR2X1_249 BUFX2_202/A XOR2X1_205/Y gnd NOR2X1_249/Y vdd NOR2X1
XNAND3X1_162 INVX1_103/A NAND3X1_162/B OR2X2_69/Y gnd OR2X2_72/B vdd NAND3X1
XBUFX2_163 OR2X2_108/A gnd BUFX2_163/Y vdd BUFX2
XCLKBUF1_40 BUFX4_4/Y gnd CLKBUF1_40/Y vdd CLKBUF1
XINVX1_578 gnd gnd INVX1_578/Y vdd INVX1
XXNOR2X1_7 XNOR2X1_7/A XNOR2X1_7/B gnd XOR2X1_28/B vdd XNOR2X1
XOAI21X1_180 NOR3X1_46/C NOR3X1_46/B NOR3X1_46/A gnd NAND3X1_189/B vdd OAI21X1
XNOR2X1_16 NOR2X1_16/A NOR2X1_16/B gnd NOR2X1_16/Y vdd NOR2X1
XXNOR2X1_201 NOR2X1_341/Y NOR2X1_340/Y gnd XOR2X1_292/A vdd XNOR2X1
XNAND2X1_294 INVX2_54/Y OAI21X1_255/Y gnd NAND2X1_294/Y vdd NAND2X1
XNOR2X1_213 BUFX2_186/A NOR2X1_213/B gnd NOR2X1_213/Y vdd NOR2X1
XNAND3X1_126 INVX1_81/A NAND3X1_126/B OR2X2_53/Y gnd OR2X2_56/B vdd NAND3X1
XNOR3X1_93 BUFX4_17/Y NOR3X1_93/B NOR3X1_93/C gnd NOR3X1_93/Y vdd NOR3X1
XDFFPOSX1_360 INVX1_448/A CLKBUF1_51/Y NAND2X1_693/Y gnd vdd DFFPOSX1
XBUFX2_127 gnd gnd BUFX2_127/Y vdd BUFX2
XINVX1_542 bloque_bytes[71] gnd INVX1_542/Y vdd INVX1
XXNOR2X1_165 NOR2X1_233/Y NOR2X1_232/Y gnd XOR2X1_211/A vdd XNOR2X1
XBUFX4_9 BUFX4_8/A gnd BUFX4_9/Y vdd BUFX4
XOAI21X1_144 NOR3X1_41/C NOR3X1_41/B INVX1_99/Y gnd OAI21X1_144/Y vdd OAI21X1
XFILL_15_7_1 gnd vdd FILL
XNOR2X1_177 NOR2X1_177/A NOR2X1_177/B gnd XOR2X1_168/A vdd NOR2X1
XFILL_17_5_0 gnd vdd FILL
XXNOR2X1_87 XNOR2X1_87/A XNOR2X1_87/B gnd OR2X2_93/A vdd XNOR2X1
XNOR3X1_57 NOR3X1_57/A NOR3X1_57/B NOR3X1_57/C gnd NOR3X1_57/Y vdd NOR3X1
XNAND2X1_258 OR2X2_101/A OR2X2_101/B gnd NAND3X1_234/B vdd NAND2X1
XINVX1_506 bloque_bytes[56] gnd INVX1_506/Y vdd INVX1
XDFFPOSX1_324 INVX1_360/A CLKBUF1_46/Y INVX1_570/Y gnd vdd DFFPOSX1
XOAI21X1_108 AOI21X1_82/Y OAI21X1_107/Y INVX1_73/Y gnd NAND3X1_112/C vdd OAI21X1
XXNOR2X1_51 AOI21X1_81/C NAND3X1_96/C gnd OR2X2_61/A vdd XNOR2X1
XXNOR2X1_129 XNOR2X1_129/A OR2X2_111/Y gnd INVX1_164/A vdd XNOR2X1
XFILL_25_2_1 gnd vdd FILL
XFILL_27_0_0 gnd vdd FILL
XFILL_5_3_1 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XNAND2X1_222 NAND2X1_222/A OR2X2_88/B gnd OR2X2_86/A vdd NAND2X1
XNOR2X1_141 NOR2X1_141/A INVX2_48/A gnd XOR2X1_130/B vdd NOR2X1
XDFFPOSX1_288 INVX1_277/A CLKBUF1_17/Y NOR2X1_429/B gnd vdd DFFPOSX1
XNOR3X1_21 BUFX4_27/Y MUX2X1_21/Y BUFX4_20/Y gnd NOR3X1_21/Y vdd NOR3X1
XOAI21X1_649 INVX2_94/Y AND2X2_197/B INVX1_595/A gnd OAI21X1_650/B vdd OAI21X1
XXOR2X1_285 AND2X2_149/Y BUFX2_233/A gnd NOR2X1_355/B vdd XOR2X1
XINVX1_470 INVX1_470/A gnd INVX1_470/Y vdd INVX1
XXNOR2X1_15 XNOR2X1_15/A NAND3X1_24/C gnd OR2X2_29/A vdd XNOR2X1
XNAND2X1_186 NAND2X1_185/Y OR2X2_71/Y gnd OR2X2_72/A vdd NAND2X1
XNOR2X1_105 NOR2X1_105/A INVX1_104/Y gnd NOR2X1_105/Y vdd NOR2X1
XAOI21X1_84 AOI21X1_84/A AOI21X1_84/B AOI21X1_84/C gnd NOR2X1_81/A vdd AOI21X1
XDFFPOSX1_252 INVX1_189/A CLKBUF1_44/Y OAI21X1_591/Y gnd vdd DFFPOSX1
XOR2X2_73 gnd OR2X2_73/B gnd OR2X2_73/Y vdd OR2X2
XINVX1_434 INVX1_434/A gnd INVX1_434/Y vdd INVX1
XOAI21X1_613 INVX1_542/Y bloque_bytes[31] INVX1_543/Y gnd AOI21X1_377/C vdd OAI21X1
XXOR2X1_249 AND2X2_133/Y BUFX2_217/A gnd XOR2X1_249/Y vdd XOR2X1
XBUFX2_87 gnd gnd BUFX2_87/Y vdd BUFX2
XAOI21X1_386 AOI21X1_386/A OR2X2_142/Y AOI21X1_386/C gnd INVX1_568/A vdd AOI21X1
XNAND2X1_150 NAND2X1_149/Y OR2X2_56/Y gnd INVX1_84/A vdd NAND2X1
XFILL_24_5_0 gnd vdd FILL
XAOI21X1_48 NAND3X1_67/A NAND3X1_64/Y AOI21X1_48/C gnd NOR2X1_51/A vdd AOI21X1
XFILL_4_6_0 gnd vdd FILL
XOR2X2_37 OR2X2_37/A OR2X2_37/B gnd OR2X2_37/Y vdd OR2X2
XDFFPOSX1_216 INVX1_138/A CLKBUF1_24/Y INVX2_89/A gnd vdd DFFPOSX1
XOAI21X1_577 INVX2_83/Y INVX2_75/Y INVX2_76/Y gnd AND2X2_170/A vdd OAI21X1
XFILL_22_7_1 gnd vdd FILL
XINVX1_398 INVX1_398/A gnd INVX1_398/Y vdd INVX1
XFILL_2_8_1 gnd vdd FILL
XBUFX2_51 gnd gnd BUFX2_51/Y vdd BUFX2
XXOR2X1_213 AND2X2_117/Y BUFX2_201/A gnd XOR2X1_213/Y vdd XOR2X1
XINVX8_1 INVX8_1/A gnd INVX8_1/Y vdd INVX8
XNAND2X1_691 NAND2X1_652/B INVX1_554/A gnd NAND2X1_691/Y vdd NAND2X1
XNAND2X1_114 NAND3X1_94/Y OAI21X1_92/Y gnd XOR2X1_59/A vdd NAND2X1
XAOI21X1_350 bloque_bytes[64] INVX1_493/Y NOR2X1_410/A gnd OAI21X1_589/C vdd AOI21X1
XNAND3X1_523 INVX1_563/A NAND3X1_523/B XNOR2X1_241/Y gnd NAND3X1_523/Y vdd NAND3X1
XFILL_34_0_0 gnd vdd FILL
XOAI21X1_1 INVX1_2/A INVX1_1/Y XNOR2X1_1/Y gnd NOR2X1_2/B vdd OAI21X1
XAOI21X1_12 AOI21X1_12/A AOI21X1_12/B NAND3X1_8/C gnd NOR2X1_21/A vdd AOI21X1
XOAI21X1_96 NOR2X1_73/B NOR2X1_73/A NAND3X1_96/A gnd OAI21X1_96/Y vdd OAI21X1
XDFFPOSX1_180 INVX1_89/A CLKBUF1_51/Y bloque_bytes[26] gnd vdd DFFPOSX1
XFILL_32_2_1 gnd vdd FILL
XXOR2X1_177 AND2X2_101/Y BUFX2_181/A gnd NOR2X1_211/B vdd XOR2X1
XOAI21X1_541 gnd NOR2X1_336/B INVX1_436/Y gnd AOI21X1_310/A vdd OAI21X1
XINVX1_362 INVX1_362/A gnd INVX1_362/Y vdd INVX1
XNAND2X1_655 bloque_bytes[39] INVX1_535/Y gnd AND2X2_177/B vdd NAND2X1
XBUFX2_15 BUFX2_15/A gnd hash[14] vdd BUFX2
XNAND2X1_75 INVX2_19/A AND2X2_18/Y gnd AOI21X1_46/C vdd NAND2X1
XOAI21X1_60 NOR2X1_53/B NOR2X1_53/A NOR3X1_31/Y gnd NAND2X1_81/B vdd OAI21X1
XDFFPOSX1_78 INVX1_480/A CLKBUF1_9/Y AOI21X1_338/Y gnd vdd DFFPOSX1
XNAND3X1_487 INVX1_468/Y INVX1_471/Y AND2X2_157/A gnd NAND2X1_608/B vdd NAND3X1
XAOI21X1_314 INVX1_451/Y AOI21X1_314/B INVX1_450/A gnd OAI21X1_545/A vdd AOI21X1
XDFFPOSX1_144 INVX1_39/A CLKBUF1_1/Y bloque_bytes[70] gnd vdd DFFPOSX1
XINVX1_326 INVX1_326/A gnd INVX1_326/Y vdd INVX1
XOAI21X1_505 OAI21X1_505/A INVX1_413/A INVX1_412/Y gnd AND2X2_145/A vdd OAI21X1
XNAND2X1_619 INVX8_1/A NOR2X1_393/B gnd NOR2X1_392/B vdd NAND2X1
XXOR2X1_141 BUFX2_166/A XOR2X1_141/B gnd XOR2X1_141/Y vdd XOR2X1
XAOI21X1_278 OAI21X1_465/Y NAND2X1_506/Y INVX2_68/A gnd AOI21X1_279/B vdd AOI21X1
XNAND2X1_39 INVX2_14/Y XNOR2X1_14/A gnd NAND3X1_24/C vdd NAND2X1
XOAI21X1_24 NOR2X1_27/A INVX1_20/Y INVX1_21/Y gnd OAI21X1_24/Y vdd OAI21X1
XDFFPOSX1_42 INVX1_501/A CLKBUF1_3/Y NOR2X1_367/Y gnd vdd DFFPOSX1
XDFFPOSX1_108 INVX1_9/A CLKBUF1_48/Y XNOR2X1_245/Y gnd vdd DFFPOSX1
XNAND3X1_451 INVX1_420/A NAND3X1_451/B NAND3X1_451/C gnd AOI21X1_303/A vdd NAND3X1
XFILL_19_2 gnd vdd FILL
XINVX1_290 INVX1_290/A gnd INVX1_290/Y vdd INVX1
XOAI21X1_469 OAI21X1_469/A INVX1_373/A INVX1_376/A gnd NAND2X1_513/A vdd OAI21X1
XXOR2X1_105 BUFX2_158/A gnd gnd OR2X2_91/B vdd XOR2X1
XXOR2X1_85 XOR2X1_99/B gnd gnd OR2X2_75/B vdd XOR2X1
XFILL_31_5_0 gnd vdd FILL
XNAND2X1_583 XOR2X1_287/B NOR2X1_340/Y gnd AOI21X1_312/C vdd NAND2X1
XFILL_29_7_1 gnd vdd FILL
XFILL_9_8_1 gnd vdd FILL
XAOI21X1_242 INVX1_280/Y NAND3X1_356/C INVX1_279/A gnd AOI21X1_242/Y vdd AOI21X1
XNAND3X1_415 INVX1_367/A INVX1_365/Y INVX1_366/Y gnd NAND3X1_420/C vdd NAND3X1
XAOI22X1_17 INVX1_371/A AOI22X1_17/B AOI22X1_17/C INVX1_369/A gnd INVX1_375/A vdd
+ AOI22X1
XXOR2X1_49 XOR2X1_49/A XOR2X1_30/Y gnd XOR2X1_49/Y vdd XOR2X1
XNAND3X1_80 OAI21X1_78/Y NAND3X1_77/Y NAND3X1_79/Y gnd NAND3X1_80/Y vdd NAND3X1
XAND2X2_185 INVX1_540/A AND2X2_185/B gnd INVX1_552/A vdd AND2X2
XINVX1_254 INVX1_254/A gnd INVX1_254/Y vdd INVX1
XOAI21X1_433 gnd NOR2X1_275/B INVX1_340/A gnd INVX2_67/A vdd OAI21X1
XOR2X2_132 bloque_bytes[73] bloque_bytes[33] gnd OR2X2_132/Y vdd OR2X2
XNAND2X1_547 OAI21X1_504/Y NAND2X1_546/Y gnd NOR2X1_320/B vdd NAND2X1
XAOI21X1_206 AOI21X1_206/A AOI21X1_206/B INVX2_59/A gnd AOI21X1_207/B vdd AOI21X1
XNAND3X1_379 AOI22X1_14/B INVX1_314/A INVX1_312/Y gnd AOI21X1_257/B vdd NAND3X1
XINVX1_218 INVX1_218/A gnd INVX1_218/Y vdd INVX1
XOAI21X1_397 gnd NOR2X1_252/B INVX1_303/A gnd INVX1_306/A vdd OAI21X1
XMUX2X1_2 BUFX2_2/A MUX2X1_2/B MUX2X1_3/S gnd NOR3X1_2/B vdd MUX2X1
XAND2X2_149 AND2X2_149/A AND2X2_149/B gnd AND2X2_149/Y vdd AND2X2
XXOR2X1_13 OR2X2_21/A gnd gnd OR2X2_17/B vdd XOR2X1
XNAND3X1_44 NAND3X1_44/A NAND3X1_42/A AOI21X1_36/C gnd NAND2X1_62/A vdd NAND3X1
XNOR2X1_430 INVX1_528/A bloque_bytes[15] gnd NOR2X1_430/Y vdd NOR2X1
XNAND2X1_511 NAND2X1_510/Y INVX1_373/Y gnd INVX1_374/A vdd NAND2X1
XAOI21X1_170 NAND3X1_245/B OR2X2_107/Y INVX1_156/A gnd NAND3X1_249/C vdd AOI21X1
XINVX1_64 OR2X2_40/Y gnd INVX1_64/Y vdd INVX1
XNAND3X1_343 INVX1_261/Y INVX1_260/A NAND3X1_343/C gnd AND2X2_113/B vdd NAND3X1
XNOR2X1_394 NOR2X1_394/A INVX2_82/A gnd NOR2X1_395/B vdd NOR2X1
XFILL_13_0_1 gnd vdd FILL
XINVX1_182 INVX1_182/A gnd OR2X2_127/B vdd INVX1
XCLKBUF1_3 BUFX4_3/Y gnd CLKBUF1_3/Y vdd CLKBUF1
XAND2X2_113 AND2X2_113/A AND2X2_113/B gnd AND2X2_113/Y vdd AND2X2
XOAI21X1_361 NOR3X1_66/A NOR3X1_66/C INVX2_63/A gnd NOR2X1_229/A vdd OAI21X1
XNAND2X1_475 OAI21X1_431/Y NAND3X1_396/Y gnd XOR2X1_241/A vdd NAND2X1
XAOI21X1_134 NAND2X1_216/Y OR2X2_83/Y INVX1_123/A gnd AOI21X1_134/Y vdd AOI21X1
XAND2X2_86 gnd OR2X2_113/B gnd NOR3X1_53/C vdd AND2X2
XNAND3X1_307 INVX1_211/A NAND2X1_347/B INVX2_60/Y gnd OAI21X1_309/B vdd NAND3X1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XINVX1_146 INVX1_146/A gnd INVX1_146/Y vdd INVX1
XFILL_36_7_1 gnd vdd FILL
XNOR2X1_358 BUFX4_13/Y INVX1_472/Y gnd NOR2X1_358/Y vdd NOR2X1
XOAI21X1_325 gnd NOR2X1_207/B INVX1_229/A gnd INVX1_231/A vdd OAI21X1
XNAND2X1_439 OAI21X1_394/Y NAND2X1_439/B gnd INVX1_346/A vdd NAND2X1
XAND2X2_50 gnd OR2X2_65/B gnd NOR3X1_41/C vdd AND2X2
XNAND3X1_271 NAND3X1_271/A OR2X2_120/B OR2X2_118/B gnd AOI21X1_185/B vdd NAND3X1
XBUFX2_272 OR2X2_85/A gnd BUFX2_272/Y vdd BUFX2
XOAI21X1_289 INVX1_194/A INVX1_195/A INVX1_196/Y gnd AOI21X1_204/A vdd OAI21X1
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XFILL_12_3_0 gnd vdd FILL
XAOI22X1_8 INVX1_200/A AOI22X1_8/B AOI22X1_8/C AOI22X1_8/D gnd INVX1_204/A vdd AOI22X1
XNOR2X1_322 gnd NOR2X1_322/B gnd AND2X2_146/A vdd NOR2X1
XNAND2X1_403 INVX1_265/Y NOR2X1_228/Y gnd NAND2X1_404/B vdd NAND2X1
XAND2X2_14 gnd OR2X2_17/B gnd AND2X2_14/Y vdd AND2X2
XFILL_10_5_1 gnd vdd FILL
XNAND3X1_235 NAND3X1_235/A OR2X2_104/B OR2X2_102/B gnd AOI21X1_161/B vdd NAND3X1
XNOR2X1_89 gnd OR2X2_58/B gnd NOR2X1_89/Y vdd NOR2X1
XBUFX2_236 BUFX2_236/A gnd BUFX2_236/Y vdd BUFX2
XINVX2_74 INVX2_74/A gnd INVX2_74/Y vdd INVX2
XOAI21X1_253 AND2X2_89/Y NOR2X1_162/Y INVX1_168/A gnd NAND3X1_265/C vdd OAI21X1
XNOR2X1_286 gnd XOR2X1_234/Y gnd NOR2X1_286/Y vdd NOR2X1
XNAND2X1_367 INVX1_229/A NOR2X1_207/Y gnd NAND3X1_321/C vdd NAND2X1
XFILL_20_0_1 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XNAND3X1_199 NAND2X1_222/A OR2X2_88/B OR2X2_86/B gnd AOI21X1_137/B vdd NAND3X1
XBUFX2_200 BUFX2_200/A gnd BUFX2_200/Y vdd BUFX2
XNOR2X1_53 NOR2X1_53/A NOR2X1_53/B gnd NOR2X1_53/Y vdd NOR2X1
XOAI21X1_217 AND2X2_76/Y NOR2X1_140/Y INVX1_145/Y gnd AOI21X1_156/A vdd OAI21X1
XXNOR2X1_238 XNOR2X1_238/A AOI21X1_354/C gnd XNOR2X1_238/Y vdd XNOR2X1
XNAND2X1_331 NAND2X1_331/A INVX1_199/A gnd XNOR2X1_148/B vdd NAND2X1
XINVX2_38 INVX2_38/A gnd INVX2_38/Y vdd INVX2
XNOR2X1_250 gnd XOR2X1_207/Y gnd AND2X2_122/A vdd NOR2X1
XXNOR2X1_8 XNOR2X1_8/A AND2X2_6/Y gnd XOR2X1_16/A vdd XNOR2X1
XNAND3X1_163 OAI21X1_156/Y OR2X2_72/B OR2X2_70/B gnd NAND3X1_163/Y vdd NAND3X1
XBUFX2_164 BUFX2_164/A gnd BUFX2_164/Y vdd BUFX2
XNOR2X1_17 NOR3X1_3/A NOR3X1_3/C gnd NOR2X1_17/Y vdd NOR2X1
XXNOR2X1_202 NOR2X1_345/Y XNOR2X1_202/B gnd XNOR2X1_202/Y vdd XNOR2X1
XINVX1_579 INVX1_579/A gnd INVX1_579/Y vdd INVX1
XCLKBUF1_41 BUFX4_2/Y gnd CLKBUF1_41/Y vdd CLKBUF1
XOAI21X1_181 NOR3X1_46/Y NOR2X1_123/A NAND3X1_185/Y gnd NAND2X1_215/B vdd OAI21X1
XNOR2X1_214 gnd NOR2X1_214/B gnd AND2X2_110/A vdd NOR2X1
XNAND2X1_295 AND2X2_90/B AND2X2_90/A gnd OAI21X1_256/B vdd NAND2X1
XBUFX2_128 gnd gnd BUFX2_128/Y vdd BUFX2
XNAND3X1_127 OAI21X1_122/Y OR2X2_56/B OR2X2_54/B gnd AOI21X1_89/B vdd NAND3X1
XNOR3X1_94 INVX1_491/A NOR3X1_91/C NOR3X1_94/C gnd NOR3X1_94/Y vdd NOR3X1
XINVX1_543 INVX1_543/A gnd INVX1_543/Y vdd INVX1
XDFFPOSX1_361 XNOR2X1_202/B CLKBUF1_22/Y OR2X2_154/Y gnd vdd DFFPOSX1
XFILL_17_5_1 gnd vdd FILL
XXNOR2X1_166 NOR2X1_237/Y XNOR2X1_166/B gnd XNOR2X1_167/A vdd XNOR2X1
XFILL_19_3_0 gnd vdd FILL
XXNOR2X1_88 XNOR2X1_88/A XNOR2X1_88/B gnd BUFX2_157/A vdd XNOR2X1
XOAI21X1_145 NOR3X1_42/Y NOR2X1_103/A NOR3X1_41/Y gnd OAI21X1_145/Y vdd OAI21X1
XNOR2X1_178 gnd NOR2X1_178/B gnd AND2X2_98/A vdd NOR2X1
XNAND2X1_259 AOI21X1_161/A AOI21X1_161/B gnd INVX2_49/A vdd NAND2X1
XFILL_10_1 gnd vdd FILL
XNOR3X1_58 NOR3X1_58/A INVX2_59/Y NOR3X1_58/C gnd NOR3X1_58/Y vdd NOR3X1
XDFFPOSX1_325 INVX1_362/A CLKBUF1_46/Y NAND2X1_675/Y gnd vdd DFFPOSX1
XINVX1_507 INVX1_507/A gnd INVX1_507/Y vdd INVX1
XOAI21X1_109 NOR2X1_77/A INVX1_75/Y INVX1_76/Y gnd OAI21X1_109/Y vdd OAI21X1
XXNOR2X1_52 XNOR2X1_52/A XNOR2X1_52/B gnd XOR2X1_78/B vdd XNOR2X1
XXNOR2X1_130 gnd XOR2X1_132/Y gnd XNOR2X1_131/A vdd XNOR2X1
XFILL_27_0_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XNAND2X1_223 OR2X2_87/B OR2X2_87/A gnd NAND2X1_223/Y vdd NAND2X1
XNOR2X1_142 AND2X2_77/A AND2X2_77/B gnd NOR2X1_142/Y vdd NOR2X1
XDFFPOSX1_289 XNOR2X1_166/B CLKBUF1_27/Y INVX1_545/Y gnd vdd DFFPOSX1
XNOR3X1_22 NOR3X1_3/A NOR3X1_22/B NOR3X1_3/C gnd NOR3X1_22/Y vdd NOR3X1
XOAI21X1_650 OAI21X1_650/A OAI21X1_650/B INVX1_597/Y gnd NAND3X1_549/C vdd OAI21X1
XXOR2X1_286 XOR2X1_286/A BUFX2_234/A gnd NOR2X1_357/B vdd XOR2X1
XINVX1_471 INVX1_471/A gnd INVX1_471/Y vdd INVX1
XXNOR2X1_16 XNOR2X1_16/A XNOR2X1_16/B gnd BUFX2_241/A vdd XNOR2X1
XNOR2X1_106 INVX1_106/Y NOR2X1_106/B gnd NOR2X1_107/B vdd NOR2X1
XFILL_32_1 gnd vdd FILL
XNAND2X1_187 OR2X2_72/B OR2X2_72/A gnd NAND2X1_187/Y vdd NAND2X1
XFILL_16_8_0 gnd vdd FILL
XAOI21X1_85 AOI21X1_85/A AOI21X1_85/B NOR3X1_38/Y gnd INVX2_30/A vdd AOI21X1
XDFFPOSX1_253 INVX1_191/A CLKBUF1_44/Y NOR2X1_412/B gnd vdd DFFPOSX1
XOAI21X1_614 AND2X2_178/Y NOR2X1_416/Y INVX1_508/A gnd OR2X2_135/A vdd OAI21X1
XINVX1_435 INVX1_435/A gnd INVX1_435/Y vdd INVX1
XOR2X2_74 gnd OR2X2_74/B gnd OR2X2_74/Y vdd OR2X2
XBUFX2_88 gnd gnd BUFX2_88/Y vdd BUFX2
XXOR2X1_250 XOR2X1_250/A BUFX2_218/A gnd NOR2X1_309/B vdd XOR2X1
XNAND2X1_151 INVX2_31/A AND2X2_42/Y gnd AOI21X1_94/C vdd NAND2X1
XAOI21X1_387 OAI21X1_624/Y OR2X2_143/Y AOI21X1_387/C gnd INVX1_569/A vdd AOI21X1
XFILL_26_3_0 gnd vdd FILL
XFILL_6_4_0 gnd vdd FILL
XDFFPOSX1_217 XOR2X1_121/B CLKBUF1_14/Y OR2X2_144/B gnd vdd DFFPOSX1
XFILL_24_5_1 gnd vdd FILL
XAOI21X1_49 AOI21X1_49/A NAND3X1_65/Y NOR2X1_53/B gnd INVX2_21/A vdd AOI21X1
XFILL_4_6_1 gnd vdd FILL
XOR2X2_38 OR2X2_38/A OR2X2_38/B gnd OR2X2_38/Y vdd OR2X2
XOAI21X1_578 INVX2_83/Y INVX1_490/A INVX8_1/A gnd NOR2X1_401/B vdd OAI21X1
XXOR2X1_214 XOR2X1_214/A BUFX2_202/A gnd XOR2X1_214/Y vdd XOR2X1
XINVX1_399 INVX1_399/A gnd INVX1_399/Y vdd INVX1
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XBUFX2_52 gnd gnd BUFX2_52/Y vdd BUFX2
XNAND2X1_692 OAI21X1_611/C INVX1_555/A gnd NAND2X1_692/Y vdd NAND2X1
XNAND2X1_115 INVX2_26/Y AOI21X1_81/B gnd NAND3X1_96/C vdd NAND2X1
XOAI21X1_97 OAI21X1_97/A XNOR2X1_52/B INVX1_74/A gnd XOR2X1_60/A vdd OAI21X1
XAOI21X1_351 bloque_bytes[65] INVX1_494/Y NOR2X1_411/A gnd OAI21X1_590/C vdd AOI21X1
XNAND3X1_524 INVX1_565/A XNOR2X1_238/Y XNOR2X1_242/Y gnd NAND3X1_524/Y vdd NAND3X1
XFILL_34_0_1 gnd vdd FILL
XOAI21X1_2 OAI21X1_2/A OAI21X1_2/B AOI21X1_2/Y gnd NAND2X1_7/B vdd OAI21X1
XAOI21X1_13 AOI21X1_13/A AOI21X1_13/B OAI21X1_9/A gnd INVX2_12/A vdd AOI21X1
XDFFPOSX1_181 INVX1_90/A CLKBUF1_18/Y bloque_bytes[27] gnd vdd DFFPOSX1
XINVX1_363 INVX1_363/A gnd INVX1_363/Y vdd INVX1
XNAND2X1_656 XNOR2X1_213/Y AND2X2_177/Y gnd NAND2X1_656/Y vdd NAND2X1
XXOR2X1_178 XOR2X1_178/A BUFX2_182/A gnd NOR2X1_213/B vdd XOR2X1
XOAI21X1_542 BUFX2_233/A NOR2X1_343/B INVX1_448/A gnd XNOR2X1_203/B vdd OAI21X1
XAOI21X1_315 INVX1_464/A AOI21X1_315/B INVX1_459/Y gnd NOR2X1_352/B vdd AOI21X1
XBUFX2_16 BUFX2_16/A gnd hash[15] vdd BUFX2
XNAND2X1_76 NAND3X1_58/Y OAI21X1_58/Y gnd XOR2X1_39/A vdd NAND2X1
XOAI21X1_61 AND2X2_21/Y NOR2X1_49/Y INVX1_45/Y gnd NAND3X1_63/B vdd OAI21X1
XNAND3X1_488 INVX1_473/A AND2X2_168/Y NOR2X1_384/A gnd INVX4_2/A vdd NAND3X1
XDFFPOSX1_79 INVX2_77/A CLKBUF1_24/Y AOI21X1_339/Y gnd vdd DFFPOSX1
XDFFPOSX1_145 XOR2X1_31/B CLKBUF1_1/Y bloque_bytes[71] gnd vdd DFFPOSX1
XINVX1_327 BUFX2_207/A gnd INVX1_327/Y vdd INVX1
XOAI21X1_506 NOR2X1_317/A NOR3X1_79/Y OAI21X1_506/C gnd NAND3X1_447/C vdd OAI21X1
XNAND2X1_620 AND2X2_164/B NOR2X1_395/B gnd NOR2X1_397/B vdd NAND2X1
XXOR2X1_142 BUFX2_171/A gnd gnd XOR2X1_142/Y vdd XOR2X1
XFILL_23_8_0 gnd vdd FILL
XNAND2X1_40 gnd OR2X2_9/B gnd NAND2X1_40/Y vdd NAND2X1
XFILL_3_9_0 gnd vdd FILL
XAOI21X1_279 NAND3X1_419/B AOI21X1_279/B INVX1_370/Y gnd AOI21X1_280/A vdd AOI21X1
XNAND3X1_452 INVX1_421/A NAND3X1_452/B INVX1_420/Y gnd INVX1_427/A vdd NAND3X1
XOAI21X1_25 AND2X2_8/Y NOR2X1_28/Y INVX1_22/Y gnd NAND2X1_41/A vdd OAI21X1
XDFFPOSX1_43 INVX1_502/A CLKBUF1_3/Y AND2X2_165/Y gnd vdd DFFPOSX1
XDFFPOSX1_109 INVX2_10/A CLKBUF1_28/Y XNOR2X1_246/Y gnd vdd DFFPOSX1
XXOR2X1_86 XOR2X1_86/A OR2X2_68/A gnd OR2X2_76/B vdd XOR2X1
XXOR2X1_106 XOR2X1_106/A OR2X2_84/A gnd OR2X2_92/B vdd XOR2X1
XINVX1_291 INVX1_291/A gnd INVX1_291/Y vdd INVX1
XFILL_33_3_0 gnd vdd FILL
XOAI21X1_470 gnd XOR2X1_243/Y INVX1_377/A gnd OAI21X1_470/Y vdd OAI21X1
XAOI22X1_18 INVX1_390/A AOI22X1_18/B AOI22X1_18/C INVX1_388/A gnd INVX1_394/A vdd
+ AOI22X1
XFILL_31_5_1 gnd vdd FILL
XNAND2X1_584 INVX1_448/Y NOR2X1_343/Y gnd NAND2X1_585/B vdd NAND2X1
XAOI21X1_243 INVX1_293/A NAND3X1_362/Y INVX1_288/Y gnd NOR2X1_244/B vdd AOI21X1
XNAND3X1_416 INVX1_369/A AOI21X1_275/B INVX1_364/Y gnd AOI22X1_17/C vdd NAND3X1
XINVX1_255 INVX1_255/A gnd INVX1_255/Y vdd INVX1
XOAI21X1_434 NOR3X1_74/C INVX2_67/Y NOR3X1_74/A gnd AND2X2_132/A vdd OAI21X1
XXOR2X1_50 XOR2X1_50/A XOR2X1_50/B gnd XOR2X1_71/A vdd XOR2X1
XNAND3X1_81 NAND3X1_79/Y OAI21X1_78/Y NOR3X1_33/Y gnd INVX1_63/A vdd NAND3X1
XAND2X2_186 INVX1_541/A AND2X2_186/B gnd INVX1_553/A vdd AND2X2
XNAND2X1_548 INVX1_409/Y NOR2X1_320/B gnd NAND2X1_548/Y vdd NAND2X1
XAOI21X1_207 NAND2X1_331/A AOI21X1_207/B INVX1_199/Y gnd AOI21X1_207/Y vdd AOI21X1
XOR2X2_133 bloque_bytes[75] bloque_bytes[35] gnd OR2X2_133/Y vdd OR2X2
XNAND3X1_380 INVX1_304/Y AOI21X1_255/A NOR3X1_70/Y gnd AOI21X1_256/B vdd NAND3X1
XMUX2X1_3 BUFX2_3/A MUX2X1_3/B MUX2X1_3/S gnd MUX2X1_3/Y vdd MUX2X1
XINVX1_219 INVX1_219/A gnd INVX1_219/Y vdd INVX1
XAND2X2_150 NOR2X1_334/Y INVX1_434/Y gnd NOR3X1_84/A vdd AND2X2
XOAI21X1_398 NOR3X1_69/A NOR3X1_69/B OAI21X1_404/B gnd NOR2X1_254/A vdd OAI21X1
XXOR2X1_14 XOR2X1_28/B gnd gnd OR2X2_18/B vdd XOR2X1
XNAND3X1_45 AOI21X1_36/C NAND3X1_44/A NOR3X1_29/Y gnd INVX1_41/A vdd NAND3X1
XNOR2X1_431 INVX1_507/A NOR2X1_431/B gnd NOR2X1_431/Y vdd NOR2X1
XNAND2X1_512 NAND2X1_512/A AOI22X1_17/C gnd NAND2X1_512/Y vdd NAND2X1
XNAND3X1_344 INVX1_259/Y INVX1_262/Y AND2X2_113/A gnd NAND3X1_344/Y vdd NAND3X1
XAOI21X1_171 NOR3X1_51/Y NOR2X1_153/Y NOR2X1_151/A gnd OAI21X1_238/C vdd AOI21X1
XFILL_30_8_0 gnd vdd FILL
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XNOR2X1_395 AND2X2_164/B NOR2X1_395/B gnd NOR2X1_395/Y vdd NOR2X1
XINVX1_183 INVX1_183/A gnd INVX1_183/Y vdd INVX1
XAND2X2_114 AND2X2_114/A INVX1_263/Y gnd NOR3X1_66/A vdd AND2X2
XOAI21X1_362 gnd XOR2X1_192/Y INVX1_267/Y gnd OAI21X1_362/Y vdd OAI21X1
XCLKBUF1_4 BUFX4_2/Y gnd CLKBUF1_4/Y vdd CLKBUF1
XNAND2X1_476 INVX1_339/Y NOR2X1_274/Y gnd NAND3X1_397/B vdd NAND2X1
XAND2X2_87 gnd OR2X2_114/B gnd AND2X2_87/Y vdd AND2X2
XAOI21X1_135 NOR3X1_45/Y NOR2X1_123/Y NOR2X1_121/A gnd OAI21X1_187/C vdd AOI21X1
XNAND3X1_308 INVX1_211/A NAND3X1_308/B NAND3X1_308/C gnd NAND2X1_350/A vdd NAND3X1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XOAI21X1_326 BUFX2_183/A INVX1_233/A INVX1_234/A gnd INVX1_236/A vdd OAI21X1
XINVX1_147 INVX1_147/A gnd INVX1_147/Y vdd INVX1
XNOR2X1_359 BUFX4_13/Y INVX2_74/Y gnd NOR2X1_359/Y vdd NOR2X1
XNAND2X1_440 INVX1_302/Y AND2X2_123/A gnd NAND3X1_371/C vdd NAND2X1
XAND2X2_51 gnd OR2X2_66/B gnd NOR3X1_42/C vdd AND2X2
XNAND3X1_272 INVX2_54/Y NAND3X1_272/B OAI21X1_255/Y gnd NAND3X1_272/Y vdd NAND3X1
XBUFX2_273 XOR2X1_94/A gnd BUFX2_273/Y vdd BUFX2
XOAI21X1_290 NOR3X1_57/C OAI21X1_284/C INVX1_199/A gnd NOR2X1_185/A vdd OAI21X1
XNOR2X1_323 gnd NOR2X1_323/B gnd NOR2X1_323/Y vdd NOR2X1
XINVX1_111 INVX1_111/A gnd INVX1_111/Y vdd INVX1
XFILL_12_3_1 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XAOI22X1_9 INVX1_219/A AOI22X1_9/B AOI22X1_9/C INVX1_217/A gnd INVX1_223/A vdd AOI22X1
XNAND2X1_404 INVX1_268/A NAND2X1_404/B gnd NOR3X1_65/B vdd NAND2X1
XAND2X2_15 gnd OR2X2_18/B gnd NOR3X1_30/C vdd AND2X2
XNAND3X1_236 INVX2_48/Y NAND3X1_236/B OAI21X1_221/Y gnd AOI21X1_163/B vdd NAND3X1
XBUFX2_237 BUFX2_237/A gnd BUFX2_237/Y vdd BUFX2
XNOR2X1_90 gnd OR2X2_59/B gnd NOR2X1_90/Y vdd NOR2X1
XOAI21X1_254 AND2X2_89/Y NOR2X1_162/Y INVX1_168/Y gnd NAND3X1_267/A vdd OAI21X1
XNAND2X1_368 INVX1_229/Y NOR2X1_207/Y gnd NAND3X1_322/B vdd NAND2X1
XINVX2_75 INVX2_75/A gnd INVX2_75/Y vdd INVX2
XNOR2X1_287 gnd NOR2X1_287/B gnd NOR2X1_287/Y vdd NOR2X1
XNAND3X1_200 INVX2_42/Y NAND3X1_200/B NAND3X1_200/C gnd AOI21X1_139/B vdd NAND3X1
XBUFX2_201 BUFX2_201/A gnd BUFX2_201/Y vdd BUFX2
XNOR2X1_54 OR2X2_29/A OR2X2_29/B gnd NOR2X1_54/Y vdd NOR2X1
XOAI21X1_218 AND2X2_76/Y NOR2X1_140/Y INVX1_145/A gnd AOI21X1_157/A vdd OAI21X1
XXNOR2X1_239 AOI21X1_379/C OR2X2_142/A gnd XNOR2X1_239/Y vdd XNOR2X1
XNAND2X1_332 INVX1_197/A NOR2X1_186/Y gnd NAND3X1_300/C vdd NAND2X1
XINVX2_39 INVX2_39/A gnd INVX2_39/Y vdd INVX2
XNOR2X1_251 gnd XOR2X1_208/Y gnd AND2X2_123/A vdd NOR2X1
XNAND3X1_164 INVX2_36/Y NAND3X1_164/B NAND3X1_164/C gnd AOI21X1_115/B vdd NAND3X1
XNOR2X1_18 gnd OR2X2_1/B gnd NOR3X1_25/B vdd NOR2X1
XXNOR2X1_9 XNOR2X1_9/A INVX2_13/Y gnd XOR2X1_17/A vdd XNOR2X1
XFILL_11_6_0 gnd vdd FILL
XBUFX2_165 BUFX2_165/A gnd BUFX2_165/Y vdd BUFX2
XCLKBUF1_42 BUFX4_2/Y gnd CLKBUF1_42/Y vdd CLKBUF1
XXNOR2X1_203 XNOR2X1_202/Y XNOR2X1_203/B gnd INVX1_452/A vdd XNOR2X1
XINVX1_580 gnd gnd INVX1_580/Y vdd INVX1
XOAI21X1_182 OAI21X1_182/A XNOR2X1_97/B INVX1_129/A gnd XOR2X1_110/A vdd OAI21X1
XNOR2X1_215 gnd NOR2X1_215/B gnd AND2X2_111/A vdd NOR2X1
XNOR3X1_95 NOR3X1_95/A OR2X2_130/Y NOR3X1_95/C gnd NOR3X1_95/Y vdd NOR3X1
XNAND2X1_296 OR2X2_117/A OR2X2_117/B gnd NAND3X1_270/B vdd NAND2X1
XBUFX2_129 gnd gnd BUFX2_129/Y vdd BUFX2
XNAND3X1_128 INVX2_30/Y AOI21X1_89/Y NAND3X1_128/C gnd AOI21X1_91/B vdd NAND3X1
XINVX1_544 INVX1_544/A gnd INVX1_544/Y vdd INVX1
XFILL_21_1_0 gnd vdd FILL
XDFFPOSX1_362 INVX1_453/A CLKBUF1_40/Y NAND3X1_520/Y gnd vdd DFFPOSX1
XFILL_1_2_0 gnd vdd FILL
XOAI21X1_146 NOR3X1_42/C NOR3X1_42/B NOR3X1_42/A gnd OAI21X1_146/Y vdd OAI21X1
XXNOR2X1_167 XNOR2X1_167/A OAI21X1_371/Y gnd INVX1_281/A vdd XNOR2X1
XFILL_19_3_1 gnd vdd FILL
XXNOR2X1_89 XNOR2X1_89/A AND2X2_60/Y gnd XOR2X1_106/A vdd XNOR2X1
XNOR2X1_179 gnd NOR2X1_179/B gnd AND2X2_99/A vdd NOR2X1
XNAND2X1_260 NAND3X1_235/A OR2X2_104/B gnd OR2X2_102/A vdd NAND2X1
XNOR3X1_59 NOR3X1_59/A NOR3X1_59/B NOR3X1_59/C gnd NOR3X1_59/Y vdd NOR3X1
XDFFPOSX1_326 INVX1_367/A CLKBUF1_8/Y NAND2X1_676/Y gnd vdd DFFPOSX1
XXNOR2X1_131 XNOR2X1_131/A INVX2_53/Y gnd INVX1_194/A vdd XNOR2X1
XINVX1_508 INVX1_508/A gnd INVX1_508/Y vdd INVX1
XOAI21X1_110 NOR3X1_37/C NOR3X1_37/B INVX1_77/Y gnd OAI21X1_110/Y vdd OAI21X1
XXNOR2X1_53 XNOR2X1_53/A AND2X2_36/Y gnd XOR2X1_66/A vdd XNOR2X1
XNAND2X1_224 NAND2X1_223/Y OR2X2_87/Y gnd OR2X2_88/A vdd NAND2X1
XNOR2X1_143 NOR2X1_143/A NOR3X1_50/Y gnd NOR2X1_143/Y vdd NOR2X1
XOAI21X1_651 NOR2X1_454/A INVX1_599/Y INVX1_600/Y gnd NAND2X1_722/B vdd OAI21X1
XINVX1_472 INVX1_472/A gnd INVX1_472/Y vdd INVX1
XDFFPOSX1_290 INVX1_282/A CLKBUF1_8/Y AOI21X1_379/C gnd vdd DFFPOSX1
XNOR3X1_23 BUFX4_27/Y NOR3X1_23/B BUFX4_20/Y gnd NOR3X1_23/Y vdd NOR3X1
XXNOR2X1_17 OAI21X1_35/A AND2X2_12/Y gnd XOR2X1_26/A vdd XNOR2X1
XXOR2X1_287 XOR2X1_287/A XOR2X1_287/B gnd XOR2X1_287/Y vdd XOR2X1
XNOR2X1_107 NOR2X1_107/A NOR2X1_107/B gnd XOR2X1_98/A vdd NOR2X1
XFILL_18_6_0 gnd vdd FILL
XFILL_32_2 gnd vdd FILL
XNAND2X1_188 NAND2X1_187/Y OR2X2_72/Y gnd INVX1_106/A vdd NAND2X1
XFILL_16_8_1 gnd vdd FILL
XAOI21X1_86 AOI21X1_86/A OR2X2_51/Y INVX1_79/A gnd AOI21X1_86/Y vdd AOI21X1
XDFFPOSX1_254 INVX1_196/A CLKBUF1_31/Y NOR2X1_413/B gnd vdd DFFPOSX1
XOAI21X1_615 AND2X2_179/Y NOR2X1_417/Y INVX1_511/A gnd OR2X2_136/A vdd OAI21X1
XINVX1_436 INVX1_436/A gnd INVX1_436/Y vdd INVX1
XOR2X2_75 gnd OR2X2_75/B gnd OR2X2_75/Y vdd OR2X2
XBUFX2_89 gnd gnd BUFX2_89/Y vdd BUFX2
XXOR2X1_251 XOR2X1_251/A XOR2X1_251/B gnd XOR2X1_251/Y vdd XOR2X1
XNAND2X1_152 NAND2X1_152/A NAND2X1_152/B gnd XOR2X1_79/A vdd NAND2X1
XAOI21X1_388 NAND2X1_673/Y AOI21X1_388/B AOI21X1_388/C gnd INVX1_570/A vdd AOI21X1
XFILL_26_3_1 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XAOI21X1_50 NAND3X1_64/B OR2X2_27/Y INVX1_46/A gnd NAND3X1_69/C vdd AOI21X1
XFILL_6_4_1 gnd vdd FILL
XFILL_8_2_0 gnd vdd FILL
XDFFPOSX1_218 INVX2_47/A CLKBUF1_3/Y INVX1_501/A gnd vdd DFFPOSX1
XOR2X2_39 OR2X2_39/A INVX1_61/Y gnd OR2X2_39/Y vdd OR2X2
XOAI21X1_579 AND2X2_171/Y AND2X2_166/B INVX8_1/A gnd AOI21X1_336/C vdd OAI21X1
XXOR2X1_215 XOR2X1_215/A XOR2X1_215/B gnd XOR2X1_215/Y vdd XOR2X1
XINVX1_400 INVX1_400/A gnd INVX1_400/Y vdd INVX1
XNAND2X1_693 AOI21X1_378/Y INVX1_556/A gnd NAND2X1_693/Y vdd NAND2X1
XBUFX2_53 gnd gnd BUFX2_53/Y vdd BUFX2
XNAND2X1_116 gnd OR2X2_41/B gnd NAND3X1_95/B vdd NAND2X1
XOAI21X1_98 AND2X2_34/Y NOR2X1_70/Y INVX1_68/Y gnd OAI21X1_98/Y vdd OAI21X1
XNAND3X1_525 INVX1_576/Y XNOR2X1_234/Y INVX1_546/A gnd NAND3X1_525/Y vdd NAND3X1
XAOI21X1_352 bloque_bytes[66] INVX1_495/Y INVX1_537/A gnd OAI21X1_591/C vdd AOI21X1
XOAI21X1_3 NOR2X1_6/Y NAND2X1_9/Y OAI21X1_3/C gnd AOI21X1_4/A vdd OAI21X1
XAOI21X1_14 AOI21X1_14/A OR2X2_3/Y INVX1_13/A gnd NAND3X1_15/C vdd AOI21X1
XDFFPOSX1_182 INVX1_91/A CLKBUF1_40/Y bloque_bytes[28] gnd vdd DFFPOSX1
XINVX1_364 INVX1_364/A gnd INVX1_364/Y vdd INVX1
XOAI21X1_543 OAI21X1_543/A INVX1_451/A INVX1_450/Y gnd AND2X2_153/A vdd OAI21X1
XNAND2X1_657 NAND2X1_657/A NOR2X1_410/Y gnd NOR2X1_431/B vdd NAND2X1
XXOR2X1_179 XOR2X1_179/A XOR2X1_179/B gnd XOR2X1_185/A vdd XOR2X1
XBUFX2_17 BUFX2_17/A gnd hash[16] vdd BUFX2
XAOI21X1_316 OAI21X1_555/Y NAND3X1_480/Y INVX1_459/A gnd NOR2X1_352/A vdd AOI21X1
XOAI21X1_62 NOR2X1_53/B NOR2X1_53/A OAI21X1_62/C gnd NAND2X1_82/B vdd OAI21X1
XDFFPOSX1_146 INVX2_20/A CLKBUF1_12/Y bloque_bytes[56] gnd vdd DFFPOSX1
XNAND2X1_77 INVX2_20/Y AOI21X1_57/B gnd NAND3X1_60/C vdd NAND2X1
XDFFPOSX1_80 INVX1_481/A CLKBUF1_16/Y DFFPOSX1_80/D gnd vdd DFFPOSX1
XNAND3X1_489 INVX1_475/Y AND2X2_169/Y INVX4_2/Y gnd AOI21X1_327/B vdd NAND3X1
XFILL_25_6_0 gnd vdd FILL
XINVX1_328 INVX1_328/A gnd INVX1_328/Y vdd INVX1
XOAI21X1_507 OAI21X1_507/A INVX1_411/A INVX1_414/A gnd NAND2X1_551/A vdd OAI21X1
XFILL_3_9_1 gnd vdd FILL
XFILL_5_7_0 gnd vdd FILL
XNAND2X1_621 BUFX4_30/Y NOR2X1_397/B gnd NOR2X1_396/B vdd NAND2X1
XXOR2X1_143 OR2X2_125/A gnd gnd AND2X2_92/B vdd XOR2X1
XFILL_23_8_1 gnd vdd FILL
XNAND2X1_41 NAND2X1_41/A NAND2X1_41/B gnd XNOR2X1_15/A vdd NAND2X1
XOAI21X1_26 NOR2X1_33/B NOR2X1_33/A NOR3X1_27/Y gnd NAND2X1_43/B vdd OAI21X1
XNAND3X1_453 INVX1_422/Y INVX1_423/Y INVX1_424/Y gnd NAND3X1_455/B vdd NAND3X1
XAOI21X1_280 AOI21X1_280/A AOI21X1_280/B NAND2X1_507/Y gnd OAI21X1_467/A vdd AOI21X1
XDFFPOSX1_44 INVX1_531/A CLKBUF1_36/Y AND2X2_166/Y gnd vdd DFFPOSX1
XINVX1_292 INVX1_292/A gnd INVX1_292/Y vdd INVX1
XFILL_35_1_0 gnd vdd FILL
XDFFPOSX1_110 INVX1_8/A CLKBUF1_28/Y AND2X2_191/Y gnd vdd DFFPOSX1
XXOR2X1_87 XOR2X1_87/A OR2X2_69/A gnd OR2X2_77/B vdd XOR2X1
XXOR2X1_107 XNOR2X1_90/Y OR2X2_85/A gnd OR2X2_93/B vdd XOR2X1
XFILL_33_3_1 gnd vdd FILL
XOAI21X1_471 gnd XOR2X1_244/Y INVX1_378/A gnd INVX2_69/A vdd OAI21X1
XNAND2X1_585 XNOR2X1_203/B NAND2X1_585/B gnd NOR2X1_344/B vdd NAND2X1
XAOI22X1_19 INVX1_409/A AOI22X1_19/B AOI22X1_19/C INVX1_407/A gnd INVX1_413/A vdd
+ AOI22X1
XAOI21X1_244 OAI21X1_384/Y NAND3X1_363/Y INVX1_288/A gnd NOR2X1_244/A vdd AOI21X1
XNAND3X1_417 INVX1_369/A OAI21X1_463/Y NAND3X1_417/C gnd NAND3X1_417/Y vdd NAND3X1
XAND2X2_187 INVX1_528/A bloque_bytes[15] gnd AND2X2_187/Y vdd AND2X2
XINVX1_256 INVX1_256/A gnd INVX1_256/Y vdd INVX1
XOAI21X1_435 gnd NOR2X1_276/B INVX1_341/A gnd INVX1_344/A vdd OAI21X1
XXOR2X1_51 XOR2X1_30/Y XOR2X1_51/B gnd XOR2X1_51/Y vdd XOR2X1
XNAND3X1_82 INVX1_57/A NAND3X1_83/B OR2X2_35/Y gnd AOI21X1_60/B vdd NAND3X1
XOR2X2_134 bloque_bytes[76] bloque_bytes[36] gnd OR2X2_134/Y vdd OR2X2
XNAND2X1_549 NAND2X1_548/Y INVX1_411/Y gnd INVX1_412/A vdd NAND2X1
XAOI21X1_208 AOI21X1_207/Y NAND3X1_302/Y AOI21X1_208/C gnd AOI21X1_208/Y vdd AOI21X1
XNAND3X1_381 INVX1_307/A OAI21X1_403/Y AOI21X1_252/B gnd NAND3X1_381/Y vdd NAND3X1
XMUX2X1_4 BUFX2_4/A MUX2X1_4/B MUX2X1_8/S gnd MUX2X1_4/Y vdd MUX2X1
XXOR2X1_15 XOR2X1_15/A gnd gnd OR2X2_19/B vdd XOR2X1
XINVX1_220 INVX1_220/A gnd INVX1_220/Y vdd INVX1
XNOR2X1_432 INVX1_510/A NOR2X1_432/B gnd NOR2X1_432/Y vdd NOR2X1
XAND2X2_151 NOR2X1_335/Y INVX1_435/Y gnd NOR3X1_84/C vdd AND2X2
XOAI21X1_399 NOR3X1_70/A NOR3X1_70/C INVX2_65/A gnd NOR2X1_253/A vdd OAI21X1
XNAND3X1_46 INVX1_35/A NAND3X1_46/B OR2X2_19/Y gnd AOI21X1_36/B vdd NAND3X1
XNAND2X1_513 NAND2X1_513/A NAND2X1_513/B gnd XOR2X1_259/A vdd NAND2X1
XAOI21X1_172 NAND3X1_248/B OR2X2_108/Y INVX1_157/A gnd OR2X2_110/B vdd AOI21X1
XNAND3X1_345 INVX2_63/A NAND3X1_345/B NAND3X1_345/C gnd NOR3X1_65/A vdd NAND3X1
XFILL_32_6_0 gnd vdd FILL
XFILL_30_8_1 gnd vdd FILL
XCLKBUF1_5 BUFX4_7/Y gnd CLKBUF1_5/Y vdd CLKBUF1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XINVX1_184 INVX1_184/A gnd INVX1_184/Y vdd INVX1
XOAI21X1_363 gnd XOR2X1_192/Y INVX1_267/A gnd INVX1_269/A vdd OAI21X1
XNAND3X1_10 INVX1_13/A AOI21X1_14/A OR2X2_3/Y gnd AOI21X1_12/B vdd NAND3X1
XNOR2X1_396 NOR2X1_395/Y NOR2X1_396/B gnd NOR2X1_396/Y vdd NOR2X1
XAND2X2_115 AND2X2_115/A INVX1_264/Y gnd NOR3X1_66/C vdd AND2X2
XNAND2X1_477 OAI21X1_432/Y NAND3X1_397/B gnd BUFX2_219/A vdd NAND2X1
XAOI21X1_136 AOI21X1_136/A OR2X2_84/Y INVX1_124/A gnd OR2X2_86/B vdd AOI21X1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XAND2X2_88 gnd OR2X2_115/B gnd AND2X2_88/Y vdd AND2X2
XNAND3X1_309 INVX1_212/A NAND3X1_309/B INVX1_211/Y gnd INVX1_218/A vdd NAND3X1
XOAI21X1_327 BUFX2_183/A INVX1_233/A INVX1_234/Y gnd OAI21X1_327/Y vdd OAI21X1
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XNOR2X1_360 BUFX4_13/Y INVX1_473/Y gnd NOR2X1_360/Y vdd NOR2X1
XNAND2X1_441 INVX1_303/Y NOR2X1_252/Y gnd NAND2X1_442/B vdd NAND2X1
XAND2X2_52 gnd OR2X2_67/B gnd AND2X2_52/Y vdd AND2X2
XNAND3X1_273 AOI21X1_189/Y NAND3X1_273/B XOR2X1_150/B gnd NAND3X1_273/Y vdd NAND3X1
XAOI21X1_100 AOI21X1_100/A OR2X2_60/Y INVX1_91/A gnd OR2X2_62/B vdd AOI21X1
XBUFX2_274 XOR2X1_90/Y gnd BUFX2_274/Y vdd BUFX2
XFILL_23_1 gnd vdd FILL
XOAI21X1_291 NOR2X1_185/Y NOR2X1_184/B AOI22X1_8/C gnd XOR2X1_170/A vdd OAI21X1
XFILL_14_1_1 gnd vdd FILL
XNOR2X1_324 gnd NOR2X1_324/B gnd NOR2X1_324/Y vdd NOR2X1
XINVX1_112 INVX1_112/A gnd INVX1_112/Y vdd INVX1
XNAND2X1_405 INVX1_267/A NOR2X1_231/Y gnd NAND2X1_405/Y vdd NAND2X1
XAND2X2_16 gnd OR2X2_19/B gnd AND2X2_16/Y vdd AND2X2
XNAND3X1_237 NAND3X1_237/A XNOR2X1_115/A XOR2X1_130/B gnd AOI21X1_166/B vdd NAND3X1
XBUFX2_238 BUFX2_238/A gnd BUFX2_238/Y vdd BUFX2
XOAI21X1_255 OAI21X1_250/A NAND3X1_258/Y AOI21X1_183/Y gnd OAI21X1_255/Y vdd OAI21X1
XNOR2X1_91 NOR2X1_91/A INVX2_33/A gnd NOR2X1_91/Y vdd NOR2X1
XNAND2X1_369 AOI21X1_223/A INVX1_237/A gnd NAND2X1_369/Y vdd NAND2X1
XINVX2_76 INVX2_76/A gnd INVX2_76/Y vdd INVX2
XNOR2X1_288 gnd XOR2X1_236/Y gnd NOR2X1_288/Y vdd NOR2X1
XNOR2X1_55 NOR2X1_55/A INVX1_49/Y gnd NOR2X1_55/Y vdd NOR2X1
XNAND3X1_201 NAND3X1_201/A XNOR2X1_97/A XOR2X1_110/B gnd AOI21X1_142/B vdd NAND3X1
XBUFX2_202 BUFX2_202/A gnd BUFX2_202/Y vdd BUFX2
XXNOR2X1_240 NAND3X1_504/Y OR2X2_143/A gnd NAND3X1_521/C vdd XNOR2X1
XOAI21X1_219 AND2X2_77/Y NOR2X1_142/Y INVX1_146/A gnd NAND3X1_229/C vdd OAI21X1
XNOR2X1_252 gnd NOR2X1_252/B gnd NOR2X1_252/Y vdd NOR2X1
XNAND2X1_333 INVX1_197/Y NOR2X1_186/Y gnd INVX1_200/A vdd NAND2X1
XINVX2_40 INVX2_40/A gnd INVX2_40/Y vdd INVX2
XNAND3X1_165 NAND3X1_165/A XNOR2X1_79/A XOR2X1_90/B gnd AOI21X1_118/B vdd NAND3X1
XFILL_13_4_0 gnd vdd FILL
XBUFX2_166 BUFX2_166/A gnd BUFX2_166/Y vdd BUFX2
XCLKBUF1_43 BUFX4_2/Y gnd CLKBUF1_43/Y vdd CLKBUF1
XINVX1_581 INVX1_581/A gnd INVX1_581/Y vdd INVX1
XNOR2X1_19 gnd OR2X2_2/B gnd NOR3X1_26/B vdd NOR2X1
XFILL_11_6_1 gnd vdd FILL
XXNOR2X1_204 NOR2X1_350/A NAND2X1_597/Y gnd INVX1_587/A vdd XNOR2X1
XOAI21X1_183 AND2X2_64/Y NOR2X1_120/Y INVX1_123/Y gnd OAI21X1_183/Y vdd OAI21X1
XNAND2X1_297 AOI21X1_185/A AOI21X1_185/B gnd INVX2_55/A vdd NAND2X1
XNOR2X1_216 gnd XOR2X1_182/Y gnd NOR2X1_216/Y vdd NOR2X1
XNOR3X1_96 BUFX4_17/Y NOR3X1_96/B NOR3X1_95/Y gnd NOR3X1_96/Y vdd NOR3X1
XDFFPOSX1_363 INVX1_454/A CLKBUF1_8/Y NAND3X1_521/Y gnd vdd DFFPOSX1
XFILL_3_0_0 gnd vdd FILL
XNAND3X1_129 AOI21X1_93/Y XNOR2X1_61/A NOR2X1_81/Y gnd AOI21X1_94/B vdd NAND3X1
XINVX1_545 INVX1_545/A gnd INVX1_545/Y vdd INVX1
XFILL_21_1_1 gnd vdd FILL
XBUFX2_130 gnd gnd BUFX2_130/Y vdd BUFX2
XFILL_1_2_1 gnd vdd FILL
XOAI21X1_147 NOR3X1_42/Y NOR2X1_103/A NAND3X1_152/B gnd NAND2X1_177/B vdd OAI21X1
XXNOR2X1_90 XNOR2X1_90/A INVX2_40/Y gnd XNOR2X1_90/Y vdd XNOR2X1
XXNOR2X1_168 NOR2X1_242/A XNOR2X1_168/B gnd BUFX2_210/A vdd XNOR2X1
XNOR2X1_180 gnd NOR2X1_180/B gnd NOR2X1_180/Y vdd NOR2X1
XNAND2X1_261 INVX1_149/Y OR2X2_103/A gnd NAND2X1_262/A vdd NAND2X1
XNOR3X1_60 NOR3X1_60/A INVX2_60/Y NOR3X1_60/C gnd NOR3X1_60/Y vdd NOR3X1
XDFFPOSX1_327 INVX1_368/A CLKBUF1_46/Y NAND2X1_677/Y gnd vdd DFFPOSX1
XINVX1_509 bloque_bytes[57] gnd INVX1_509/Y vdd INVX1
XXNOR2X1_132 NAND2X1_288/Y NAND3X1_258/C gnd BUFX2_176/A vdd XNOR2X1
XOAI21X1_111 NOR3X1_38/Y NOR2X1_83/A NOR3X1_37/Y gnd OAI21X1_111/Y vdd OAI21X1
XXNOR2X1_54 XNOR2X1_54/A INVX2_28/Y gnd XOR2X1_67/A vdd XNOR2X1
XFILL_10_9_0 gnd vdd FILL
XNOR2X1_144 OR2X2_101/A OR2X2_101/B gnd NOR2X1_144/Y vdd NOR2X1
XNAND2X1_225 OR2X2_88/B OR2X2_88/A gnd NAND2X1_226/A vdd NAND2X1
XNOR3X1_24 NOR3X1_3/A MUX2X1_24/Y NOR3X1_3/C gnd NOR3X1_24/Y vdd NOR3X1
XINVX1_473 INVX1_473/A gnd INVX1_473/Y vdd INVX1
XDFFPOSX1_291 INVX1_283/A CLKBUF1_23/Y NAND3X1_504/Y gnd vdd DFFPOSX1
XXNOR2X1_18 OAI21X1_35/Y INVX2_16/Y gnd XOR2X1_27/A vdd XNOR2X1
XXOR2X1_288 BUFX2_243/A gnd gnd INVX1_584/A vdd XOR2X1
XNAND2X1_189 INVX2_37/A AND2X2_54/Y gnd NAND2X1_189/Y vdd NAND2X1
XFILL_18_6_1 gnd vdd FILL
XFILL_20_4_0 gnd vdd FILL
XNOR2X1_108 gnd OR2X2_73/B gnd NOR3X1_43/B vdd NOR2X1
XFILL_0_5_0 gnd vdd FILL
XAOI21X1_87 NOR3X1_37/Y NOR2X1_83/Y NOR2X1_81/A gnd AOI21X1_87/Y vdd AOI21X1
XDFFPOSX1_255 INVX1_197/A CLKBUF1_11/Y INVX1_576/A gnd vdd DFFPOSX1
XOAI21X1_616 NOR2X1_418/Y NOR2X1_419/Y INVX1_514/A gnd NOR2X1_427/B vdd OAI21X1
XOR2X2_76 OR2X2_76/A OR2X2_76/B gnd OR2X2_76/Y vdd OR2X2
XXOR2X1_252 BUFX2_223/A gnd gnd NOR2X1_310/B vdd XOR2X1
XINVX1_437 INVX1_437/A gnd INVX1_437/Y vdd INVX1
XBUFX2_90 gnd gnd BUFX2_90/Y vdd BUFX2
XFILL_28_1_1 gnd vdd FILL
XFILL_8_2_1 gnd vdd FILL
XAOI21X1_389 AOI21X1_389/A OR2X2_144/Y NAND3X1_513/Y gnd INVX1_573/A vdd AOI21X1
XNAND2X1_153 INVX2_32/Y XNOR2X1_67/Y gnd XNOR2X1_69/B vdd NAND2X1
XAOI21X1_51 NOR3X1_31/Y NOR2X1_53/Y NOR2X1_51/A gnd OAI21X1_68/C vdd AOI21X1
XOR2X2_40 OR2X2_40/A OR2X2_40/B gnd OR2X2_40/Y vdd OR2X2
XDFFPOSX1_219 INVX1_143/A CLKBUF1_30/Y INVX1_502/A gnd vdd DFFPOSX1
XINVX1_401 INVX1_401/A gnd INVX1_401/Y vdd INVX1
XOAI21X1_580 AND2X2_172/Y INVX1_480/A INVX8_2/A gnd OAI21X1_580/Y vdd OAI21X1
XXOR2X1_216 BUFX2_207/A gnd gnd NOR2X1_262/B vdd XOR2X1
XNAND2X1_694 gnd gnd gnd INVX1_579/A vdd NAND2X1
XAOI21X1_353 bloque_bytes[67] INVX1_496/Y AOI21X1_353/C gnd OAI21X1_592/C vdd AOI21X1
XBUFX2_54 gnd gnd BUFX2_54/Y vdd BUFX2
XOAI21X1_4 INVX1_1/Y INVX1_2/A NOR2X1_7/Y gnd OAI21X1_5/C vdd OAI21X1
XNAND2X1_117 OAI21X1_93/Y NAND3X1_96/A gnd AOI21X1_81/C vdd NAND2X1
XOAI21X1_99 AND2X2_34/Y NOR2X1_70/Y INVX1_68/A gnd OAI21X1_99/Y vdd OAI21X1
XNAND3X1_526 INVX1_577/Y NAND3X1_526/B INVX1_566/A gnd NAND3X1_526/Y vdd NAND3X1
XAOI21X1_15 NOR3X1_25/Y NOR2X1_23/Y NOR2X1_21/A gnd OAI21X1_17/C vdd AOI21X1
XDFFPOSX1_183 INVX1_92/A CLKBUF1_18/Y bloque_bytes[29] gnd vdd DFFPOSX1
XFILL_17_9_0 gnd vdd FILL
XINVX1_365 BUFX2_215/A gnd INVX1_365/Y vdd INVX1
XOAI21X1_544 NOR2X1_341/A NOR3X1_83/Y AOI21X1_313/Y gnd AOI21X1_314/B vdd OAI21X1
XXOR2X1_180 INVX1_251/A gnd gnd NOR2X1_214/B vdd XOR2X1
XNAND2X1_658 XNOR2X1_215/Y NOR2X1_411/Y gnd NOR2X1_432/B vdd NAND2X1
XBUFX2_18 BUFX2_18/A gnd hash[17] vdd BUFX2
XNAND2X1_78 gnd OR2X2_25/B gnd NAND3X1_59/B vdd NAND2X1
XNAND3X1_490 NOR2X1_381/Y NOR2X1_387/Y NOR2X1_388/Y gnd INVX2_82/A vdd NAND3X1
XAOI21X1_317 INVX1_459/A AOI21X1_317/B INVX1_458/Y gnd NOR3X1_85/C vdd AOI21X1
XOAI21X1_63 OAI21X1_63/A OAI21X1_68/B INVX1_52/A gnd XOR2X1_40/A vdd OAI21X1
XDFFPOSX1_147 INVX1_44/A CLKBUF1_12/Y bloque_bytes[57] gnd vdd DFFPOSX1
XDFFPOSX1_81 INVX1_482/A CLKBUF1_15/Y DFFPOSX1_81/D gnd vdd DFFPOSX1
XFILL_27_4_0 gnd vdd FILL
XFILL_7_5_0 gnd vdd FILL
XXOR2X1_144 BUFX2_173/A gnd gnd OR2X2_122/B vdd XOR2X1
XFILL_25_6_1 gnd vdd FILL
XOAI21X1_508 gnd NOR2X1_322/B INVX1_415/A gnd NAND2X1_553/A vdd OAI21X1
XINVX1_329 INVX1_329/A gnd INVX1_329/Y vdd INVX1
XFILL_5_7_1 gnd vdd FILL
XNAND2X1_622 AND2X2_164/B INVX1_478/A gnd NOR2X1_398/B vdd NAND2X1
XOAI21X1_27 AND2X2_9/Y NOR3X1_28/B INVX1_23/Y gnd NAND3X1_26/A vdd OAI21X1
XNAND2X1_42 gnd AND2X2_9/B gnd NAND3X1_25/B vdd NAND2X1
XDFFPOSX1_45 INVX1_503/A CLKBUF1_30/Y NOR2X1_368/Y gnd vdd DFFPOSX1
XNAND3X1_454 INVX1_424/A INVX1_422/Y INVX1_423/Y gnd AOI21X1_300/B vdd NAND3X1
XAOI21X1_281 NAND3X1_417/Y AOI21X1_281/B NAND2X1_512/Y gnd AOI21X1_281/Y vdd AOI21X1
XINVX1_293 INVX1_293/A gnd INVX1_293/Y vdd INVX1
XFILL_35_1_1 gnd vdd FILL
XDFFPOSX1_111 INVX1_7/A CLKBUF1_43/Y XNOR2X1_247/Y gnd vdd DFFPOSX1
XOAI21X1_472 NOR3X1_78/C INVX2_69/Y NOR3X1_78/A gnd AND2X2_140/A vdd OAI21X1
XXOR2X1_108 XOR2X1_108/A XOR2X1_94/A gnd XOR2X1_108/Y vdd XOR2X1
XXOR2X1_88 NOR2X1_97/Y XOR2X1_74/A gnd XOR2X1_88/Y vdd XOR2X1
XNAND2X1_586 INVX1_447/Y NOR2X1_344/B gnd NAND2X1_587/A vdd NAND2X1
XAOI21X1_245 INVX1_288/A AOI21X1_245/B INVX1_287/Y gnd NOR3X1_67/C vdd AOI21X1
XAOI22X1_20 INVX1_428/A AOI22X1_20/B AOI22X1_20/C INVX1_426/A gnd INVX1_432/A vdd
+ AOI22X1
XNAND3X1_418 AOI22X1_17/B INVX1_371/A INVX1_369/Y gnd AOI21X1_281/B vdd NAND3X1
XINVX1_257 INVX1_257/A gnd INVX1_257/Y vdd INVX1
XOAI21X1_436 NOR3X1_73/A INVX1_342/A OAI21X1_442/B gnd NOR2X1_278/A vdd OAI21X1
XAND2X2_188 AND2X2_188/A BUFX2_243/A gnd AND2X2_189/A vdd AND2X2
XXOR2X1_52 OR2X2_52/A gnd gnd XOR2X1_52/Y vdd XOR2X1
XNAND3X1_83 INVX1_57/Y NAND3X1_83/B OR2X2_35/Y gnd AOI21X1_61/B vdd NAND3X1
XOR2X2_135 OR2X2_135/A bloque_bytes[8] gnd OR2X2_145/A vdd OR2X2
XNAND2X1_550 NAND2X1_550/A AOI22X1_19/C gnd NAND2X1_550/Y vdd NAND2X1
XAOI21X1_209 NAND2X1_334/A NAND2X1_334/B AOI21X1_209/C gnd OAI21X1_297/C vdd AOI21X1
XFILL_24_9_0 gnd vdd FILL
XNAND3X1_382 INVX1_318/Y INVX1_317/A NAND3X1_382/C gnd AND2X2_125/B vdd NAND3X1
XMUX2X1_5 BUFX2_5/A MUX2X1_5/B MUX2X1_3/S gnd MUX2X1_5/Y vdd MUX2X1
XNAND3X1_47 INVX1_35/Y NAND3X1_46/B OR2X2_19/Y gnd AOI21X1_37/B vdd NAND3X1
XXOR2X1_16 XOR2X1_16/A XOR2X1_2/A gnd OR2X2_20/B vdd XOR2X1
XINVX1_221 INVX1_221/A gnd INVX1_221/Y vdd INVX1
XNOR2X1_433 INVX1_513/A NOR2X1_433/B gnd NOR2X1_433/Y vdd NOR2X1
XOAI21X1_400 gnd XOR2X1_210/Y INVX1_305/Y gnd OAI21X1_400/Y vdd OAI21X1
XNAND2X1_514 INVX1_377/Y NOR2X1_298/Y gnd NAND3X1_423/B vdd NAND2X1
XAND2X2_152 AND2X2_152/A NOR3X1_83/A gnd BUFX2_244/A vdd AND2X2
XFILL_34_4_0 gnd vdd FILL
XFILL_32_6_1 gnd vdd FILL
XAOI21X1_173 AOI21X1_173/A AOI21X1_173/B OAI21X1_239/B gnd NAND3X1_254/B vdd AOI21X1
XNAND3X1_346 INVX1_268/A NAND2X1_404/B INVX2_63/Y gnd OAI21X1_366/B vdd NAND3X1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XCLKBUF1_6 BUFX4_7/Y gnd CLKBUF1_6/Y vdd CLKBUF1
XINVX1_185 INVX1_185/A gnd INVX1_185/Y vdd INVX1
XOAI21X1_364 BUFX2_191/A INVX1_271/A INVX1_272/A gnd INVX1_274/A vdd OAI21X1
XAND2X2_116 AND2X2_116/A NOR3X1_65/A gnd BUFX2_204/A vdd AND2X2
XNAND3X1_11 INVX1_13/Y AOI21X1_14/A OR2X2_3/Y gnd AOI21X1_13/B vdd NAND3X1
XNOR2X1_397 INVX1_478/Y NOR2X1_397/B gnd NOR3X1_88/C vdd NOR2X1
XNAND2X1_478 INVX1_340/Y NOR2X1_275/Y gnd NAND2X1_478/Y vdd NAND2X1
XAND2X2_89 AND2X2_89/A AND2X2_89/B gnd AND2X2_89/Y vdd AND2X2
XAOI21X1_137 AOI21X1_137/A AOI21X1_137/B AOI21X1_137/C gnd NAND3X1_200/B vdd AOI21X1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XNAND3X1_310 INVX1_213/Y INVX1_214/Y INVX1_215/Y gnd NAND3X1_312/B vdd NAND3X1
XFILL_1_1 gnd vdd FILL
XNOR2X1_361 BUFX4_13/Y INVX1_474/Y gnd NOR2X1_361/Y vdd NOR2X1
XINVX1_149 INVX1_149/A gnd INVX1_149/Y vdd INVX1
XOAI21X1_328 NOR3X1_61/C OAI21X1_328/B INVX1_237/A gnd NOR2X1_209/A vdd OAI21X1
XNAND2X1_442 INVX1_306/A NAND2X1_442/B gnd NOR3X1_69/B vdd NAND2X1
XAND2X2_53 OR2X2_68/A OR2X2_68/B gnd AND2X2_53/Y vdd AND2X2
XNAND3X1_274 INVX1_174/A INVX1_175/A NAND3X1_274/C gnd NAND2X1_304/A vdd NAND3X1
XAOI21X1_101 NAND3X1_143/Y NAND3X1_145/Y AOI21X1_101/C gnd NAND3X1_146/B vdd AOI21X1
XOAI21X1_292 BUFX2_176/A NOR2X1_186/B INVX1_197/Y gnd NAND3X1_300/B vdd OAI21X1
XINVX1_113 INVX1_113/A gnd INVX1_113/Y vdd INVX1
XFILL_31_9_0 gnd vdd FILL
XNAND2X1_406 INVX1_267/Y NOR2X1_231/Y gnd AOI21X1_237/B vdd NAND2X1
XNOR2X1_325 NOR2X1_325/A INVX1_418/Y gnd NOR2X1_325/Y vdd NOR2X1
XBUFX2_239 OR2X2_28/A gnd BUFX2_239/Y vdd BUFX2
XAND2X2_17 OR2X2_20/A OR2X2_20/B gnd AND2X2_17/Y vdd AND2X2
XNAND3X1_238 OR2X2_104/Y INVX1_153/A NAND3X1_238/C gnd NAND2X1_266/A vdd NAND3X1
XOAI21X1_256 NAND2X1_294/Y OAI21X1_256/B AND2X2_90/B gnd OAI21X1_256/Y vdd OAI21X1
XNOR2X1_92 OR2X2_60/A OR2X2_60/B gnd NOR2X1_92/Y vdd NOR2X1
XINVX2_77 INVX2_77/A gnd INVX2_77/Y vdd INVX2
XNAND2X1_370 INVX1_235/A NOR2X1_210/Y gnd NAND3X1_326/C vdd NAND2X1
XNOR2X1_289 NOR2X1_289/A INVX1_361/Y gnd NOR2X1_289/Y vdd NOR2X1
XNAND3X1_202 OR2X2_88/Y INVX1_131/A NAND3X1_202/C gnd NAND2X1_228/A vdd NAND3X1
XNOR2X1_56 INVX1_51/Y NOR2X1_56/B gnd NOR2X1_57/B vdd NOR2X1
XXNOR2X1_241 AOI21X1_382/C NOR2X1_412/B gnd XNOR2X1_241/Y vdd XNOR2X1
XBUFX2_203 BUFX2_203/A gnd BUFX2_203/Y vdd BUFX2
XINVX2_41 INVX2_41/A gnd INVX2_41/Y vdd INVX2
XOAI21X1_220 AND2X2_77/Y NOR2X1_142/Y INVX1_146/Y gnd NAND3X1_233/A vdd OAI21X1
XNOR2X1_253 NOR2X1_253/A INVX1_304/Y gnd NOR2X1_254/B vdd NOR2X1
XNAND2X1_334 NAND2X1_334/A NAND2X1_334/B gnd XOR2X1_170/B vdd NAND2X1
XFILL_15_2_0 gnd vdd FILL
XCLKBUF1_44 BUFX4_1/Y gnd CLKBUF1_44/Y vdd CLKBUF1
XNAND3X1_166 OR2X2_72/Y INVX1_109/A NAND3X1_166/C gnd NAND3X1_166/Y vdd NAND3X1
XBUFX2_167 AND2X2_89/A gnd BUFX2_167/Y vdd BUFX2
XFILL_13_4_1 gnd vdd FILL
XINVX1_582 INVX1_582/A gnd INVX1_582/Y vdd INVX1
XNOR2X1_20 gnd OR2X2_3/B gnd NOR2X1_20/Y vdd NOR2X1
XOAI21X1_184 AND2X2_64/Y NOR2X1_120/Y INVX1_123/A gnd AOI21X1_133/A vdd OAI21X1
XXNOR2X1_205 NOR2X1_353/Y NOR2X1_352/Y gnd INVX1_588/A vdd XNOR2X1
XNAND2X1_298 NAND3X1_271/A OR2X2_120/B gnd OR2X2_118/A vdd NAND2X1
XNOR2X1_217 NOR2X1_217/A INVX1_247/Y gnd NOR2X1_218/B vdd NOR2X1
XNOR3X1_97 INVX1_590/Y NOR3X1_97/B NOR3X1_97/C gnd NOR3X1_97/Y vdd NOR3X1
XDFFPOSX1_364 INVX1_455/A CLKBUF1_22/Y NAND3X1_522/Y gnd vdd DFFPOSX1
XBUFX2_131 gnd gnd BUFX2_131/Y vdd BUFX2
XFILL_3_0_1 gnd vdd FILL
XNAND3X1_130 OR2X2_56/Y INVX1_87/A NAND3X1_130/C gnd NAND2X1_152/A vdd NAND3X1
XINVX1_546 INVX1_546/A gnd INVX1_546/Y vdd INVX1
XXNOR2X1_169 NOR2X1_245/Y NOR2X1_244/Y gnd XOR2X1_220/A vdd XNOR2X1
XOAI21X1_148 OAI21X1_153/A XNOR2X1_79/B INVX1_107/A gnd XOR2X1_90/A vdd OAI21X1
XNOR2X1_181 NOR2X1_181/A INVX1_190/Y gnd NOR2X1_182/B vdd NOR2X1
XXNOR2X1_91 XOR2X1_98/B XOR2X1_88/Y gnd OR2X2_79/A vdd XNOR2X1
XNAND2X1_262 NAND2X1_262/A OR2X2_103/Y gnd OR2X2_104/A vdd NAND2X1
XNOR3X1_61 NOR3X1_61/A NOR3X1_61/B NOR3X1_61/C gnd NOR3X1_61/Y vdd NOR3X1
XINVX1_510 INVX1_510/A gnd INVX1_510/Y vdd INVX1
XDFFPOSX1_328 INVX1_372/A CLKBUF1_2/Y NAND2X1_678/Y gnd vdd DFFPOSX1
XXNOR2X1_55 BUFX2_253/A XOR2X1_48/Y gnd OR2X2_47/A vdd XNOR2X1
XXNOR2X1_133 NAND3X1_273/B NAND3X1_258/Y gnd BUFX2_177/A vdd XNOR2X1
XOAI21X1_112 NOR3X1_38/C NOR2X1_79/Y INVX1_78/Y gnd OAI21X1_112/Y vdd OAI21X1
XFILL_10_9_1 gnd vdd FILL
XFILL_12_7_0 gnd vdd FILL
XNAND2X1_226 NAND2X1_226/A OR2X2_88/Y gnd INVX1_128/A vdd NAND2X1
XNOR2X1_145 NOR2X1_145/A INVX1_148/Y gnd NOR2X1_145/Y vdd NOR2X1
XNOR3X1_25 INVX1_11/Y NOR3X1_25/B AND2X2_2/Y gnd NOR3X1_25/Y vdd NOR3X1
XDFFPOSX1_292 INVX1_284/A CLKBUF1_2/Y AOI21X1_381/C gnd vdd DFFPOSX1
XINVX1_474 INVX1_474/A gnd INVX1_474/Y vdd INVX1
XXNOR2X1_19 XOR2X1_4/A XOR2X1_8/Y gnd OR2X2_15/A vdd XNOR2X1
XFILL_20_4_1 gnd vdd FILL
XFILL_22_2_0 gnd vdd FILL
XXOR2X1_289 BUFX2_244/A gnd gnd XOR2X1_289/Y vdd XOR2X1
XFILL_0_5_1 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XNAND2X1_190 NAND3X1_166/Y OAI21X1_160/Y gnd XOR2X1_99/A vdd NAND2X1
XNOR2X1_109 gnd OR2X2_74/B gnd NOR3X1_44/B vdd NOR2X1
XAOI21X1_88 AOI21X1_88/A OR2X2_52/Y INVX1_80/A gnd OR2X2_54/B vdd AOI21X1
XDFFPOSX1_256 INVX1_201/A CLKBUF1_11/Y INVX1_577/A gnd vdd DFFPOSX1
XOAI21X1_617 AND2X2_180/Y NOR2X1_420/Y INVX1_517/A gnd OR2X2_137/A vdd OAI21X1
XOR2X2_77 OR2X2_77/A OR2X2_77/B gnd OR2X2_77/Y vdd OR2X2
XINVX1_438 INVX1_438/A gnd INVX1_438/Y vdd INVX1
XXOR2X1_253 BUFX2_224/A gnd gnd NOR2X1_311/B vdd XOR2X1
XBUFX2_91 gnd gnd BUFX2_91/Y vdd BUFX2
XAOI21X1_390 NAND2X1_657/A NOR2X1_410/Y INVX1_507/Y gnd OAI21X1_626/B vdd AOI21X1
XNAND2X1_154 gnd OR2X2_57/B gnd NAND2X1_154/Y vdd NAND2X1
XAOI21X1_52 AOI21X1_52/A OR2X2_28/Y INVX1_47/A gnd OR2X2_30/B vdd AOI21X1
XOR2X2_41 gnd OR2X2_41/B gnd OR2X2_41/Y vdd OR2X2
XOAI21X1_581 INVX2_83/Y INVX2_84/A BUFX4_32/Y gnd AOI21X1_339/C vdd OAI21X1
XDFFPOSX1_220 INVX1_144/A CLKBUF1_36/Y INVX1_531/A gnd vdd DFFPOSX1
XINVX1_402 INVX1_402/A gnd INVX1_402/Y vdd INVX1
XBUFX2_55 gnd gnd BUFX2_55/Y vdd BUFX2
XXOR2X1_217 BUFX2_208/A gnd gnd XOR2X1_217/Y vdd XOR2X1
XNAND2X1_695 gnd INVX1_579/Y gnd XNOR2X1_244/A vdd NAND2X1
XNAND2X1_118 gnd OR2X2_42/B gnd NAND3X1_97/B vdd NAND2X1
XAOI21X1_354 bloque_bytes[68] INVX1_497/Y AOI21X1_354/C gnd OAI21X1_593/C vdd AOI21X1
XOAI21X1_5 INVX2_8/Y NOR2X1_1/B OAI21X1_5/C gnd OAI21X1_5/Y vdd OAI21X1
XDFFPOSX1_184 INVX1_94/A CLKBUF1_29/Y bloque_bytes[30] gnd vdd DFFPOSX1
XNAND3X1_527 INVX1_543/Y AOI21X1_393/B INVX1_567/A gnd NAND3X1_527/Y vdd NAND3X1
XFILL_19_7_0 gnd vdd FILL
XAOI21X1_16 NAND3X1_14/B OR2X2_4/Y INVX1_14/A gnd OR2X2_6/B vdd AOI21X1
XFILL_17_9_1 gnd vdd FILL
XXOR2X1_181 BUFX2_188/A gnd gnd NOR2X1_215/B vdd XOR2X1
XINVX1_366 INVX1_366/A gnd INVX1_366/Y vdd INVX1
XOAI21X1_545 OAI21X1_545/A INVX1_449/A INVX1_452/A gnd NAND2X1_589/A vdd OAI21X1
XFILL_14_1 gnd vdd FILL
XNAND2X1_659 XNOR2X1_216/Y NAND2X1_659/B gnd NOR2X1_433/B vdd NAND2X1
XBUFX2_19 BUFX2_19/A gnd hash[18] vdd BUFX2
XOAI21X1_64 AND2X2_22/Y NOR2X1_50/Y INVX1_46/Y gnd NAND3X1_67/A vdd OAI21X1
XNAND2X1_79 NAND3X1_60/B OAI21X1_62/C gnd AOI21X1_57/C vdd NAND2X1
XNAND3X1_491 AND2X2_161/B INVX1_476/A AND2X2_162/B gnd INVX1_488/A vdd NAND3X1
XAOI21X1_318 AOI21X1_318/A NAND2X1_601/Y INVX2_73/A gnd AOI21X1_319/B vdd AOI21X1
XFILL_29_2_0 gnd vdd FILL
XDFFPOSX1_148 INVX1_45/A CLKBUF1_1/Y bloque_bytes[58] gnd vdd DFFPOSX1
XFILL_9_3_0 gnd vdd FILL
XDFFPOSX1_82 INVX2_78/A CLKBUF1_6/Y AOI21X1_342/Y gnd vdd DFFPOSX1
XFILL_27_4_1 gnd vdd FILL
XINVX1_330 INVX1_330/A gnd INVX1_330/Y vdd INVX1
XFILL_7_5_1 gnd vdd FILL
XNAND2X1_623 INVX1_489/Y NOR2X1_398/Y gnd INVX1_491/A vdd NAND2X1
XXOR2X1_145 BUFX2_174/A gnd gnd OR2X2_123/B vdd XOR2X1
XOAI21X1_509 gnd NOR2X1_323/B INVX1_416/A gnd INVX2_71/A vdd OAI21X1
XAOI21X1_282 INVX1_375/Y AOI21X1_282/B INVX1_374/A gnd OAI21X1_469/A vdd AOI21X1
XOAI21X1_28 NOR2X1_33/B NOR2X1_33/A NAND2X1_41/B gnd OAI21X1_28/Y vdd OAI21X1
XNAND2X1_43 NAND3X1_26/Y NAND2X1_43/B gnd XNOR2X1_16/A vdd NAND2X1
XDFFPOSX1_46 INVX1_504/A CLKBUF1_3/Y NOR2X1_369/Y gnd vdd DFFPOSX1
XNAND3X1_455 INVX1_426/A NAND3X1_455/B INVX1_421/Y gnd AOI22X1_20/C vdd NAND3X1
XINVX1_294 INVX1_294/A gnd INVX1_294/Y vdd INVX1
XFILL_36_1 gnd vdd FILL
XOAI21X1_473 gnd NOR2X1_300/B INVX1_379/A gnd INVX1_382/A vdd OAI21X1
XDFFPOSX1_112 INVX1_6/A CLKBUF1_28/Y XNOR2X1_248/Y gnd vdd DFFPOSX1
XXOR2X1_109 XOR2X1_109/A XOR2X1_90/Y gnd XOR2X1_109/Y vdd XOR2X1
XXOR2X1_89 XOR2X1_89/A XOR2X1_75/A gnd XOR2X1_89/Y vdd XOR2X1
XNAND2X1_587 NAND2X1_587/A INVX1_449/Y gnd INVX1_450/A vdd NAND2X1
XAOI21X1_246 OAI21X1_389/Y AOI21X1_246/B INVX2_64/A gnd AOI21X1_247/B vdd AOI21X1
XNAND3X1_419 INVX1_361/Y NAND3X1_419/B NOR3X1_76/Y gnd AOI21X1_280/B vdd NAND3X1
XAOI22X1_21 INVX1_447/A AOI22X1_21/B AOI22X1_21/C INVX1_445/A gnd INVX1_451/A vdd
+ AOI22X1
XDFFPOSX1_10 BUFX2_9/A CLKBUF1_41/Y NOR3X1_9/Y gnd vdd DFFPOSX1
XXOR2X1_53 OR2X2_53/A gnd gnd OR2X2_49/B vdd XOR2X1
XINVX1_258 INVX1_258/A gnd INVX1_258/Y vdd INVX1
XOAI21X1_437 NOR3X1_74/A NOR3X1_74/C INVX2_67/A gnd NOR2X1_277/A vdd OAI21X1
XAND2X2_189 AND2X2_189/A BUFX2_244/A gnd XOR2X1_306/A vdd AND2X2
XNAND3X1_84 INVX1_58/Y NAND3X1_84/B OR2X2_36/Y gnd NAND3X1_84/Y vdd NAND3X1
XFILL_24_9_1 gnd vdd FILL
XOR2X2_136 OR2X2_136/A bloque_bytes[9] gnd OR2X2_151/A vdd OR2X2
XFILL_26_7_0 gnd vdd FILL
XNAND2X1_551 NAND2X1_551/A NAND2X1_551/B gnd XOR2X1_277/A vdd NAND2X1
XFILL_6_8_0 gnd vdd FILL
XAOI21X1_210 INVX1_204/Y OAI21X1_297/Y INVX1_203/A gnd AOI21X1_210/Y vdd AOI21X1
XNAND3X1_383 INVX1_316/Y INVX1_319/Y AND2X2_125/A gnd NAND3X1_383/Y vdd NAND3X1
XINVX1_222 INVX1_222/A gnd INVX1_222/Y vdd INVX1
XMUX2X1_6 BUFX2_6/A MUX2X1_6/B MUX2X1_8/S gnd NOR3X1_6/B vdd MUX2X1
XOAI21X1_401 gnd XOR2X1_210/Y INVX1_305/A gnd INVX1_307/A vdd OAI21X1
XNAND3X1_48 INVX1_36/Y NAND3X1_50/B OR2X2_20/Y gnd NAND3X1_49/B vdd NAND3X1
XXOR2X1_17 XOR2X1_17/A XOR2X1_3/A gnd OR2X2_21/B vdd XOR2X1
XNOR2X1_434 INVX1_528/A NOR2X1_434/B gnd NOR2X1_434/Y vdd NOR2X1
XFILL_36_2_0 gnd vdd FILL
XNAND2X1_515 OAI21X1_470/Y NAND3X1_423/B gnd INVX1_422/A vdd NAND2X1
XAND2X2_153 AND2X2_153/A AND2X2_153/B gnd XOR2X1_294/A vdd AND2X2
XOR2X2_100 AND2X2_77/A AND2X2_77/B gnd OR2X2_100/Y vdd OR2X2
XAOI21X1_174 OR2X2_110/B OR2X2_110/A AND2X2_84/B gnd NOR2X1_155/A vdd AOI21X1
XFILL_34_4_1 gnd vdd FILL
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XNAND3X1_347 INVX1_268/A OAI21X1_362/Y NAND2X1_405/Y gnd NAND3X1_347/Y vdd NAND3X1
XCLKBUF1_7 BUFX4_1/Y gnd CLKBUF1_7/Y vdd CLKBUF1
XINVX1_186 INVX1_186/A gnd INVX1_186/Y vdd INVX1
XOAI21X1_365 BUFX2_191/A INVX1_271/A INVX1_272/Y gnd AOI21X1_236/A vdd OAI21X1
XAND2X2_117 AND2X2_117/A AND2X2_117/B gnd AND2X2_117/Y vdd AND2X2
XNAND3X1_12 INVX1_14/Y NAND3X1_14/B OR2X2_4/Y gnd NAND3X1_12/Y vdd NAND3X1
XNOR2X1_398 NOR2X1_398/A NOR2X1_398/B gnd NOR2X1_398/Y vdd NOR2X1
XNAND2X1_479 INVX1_341/Y NOR2X1_276/Y gnd NAND2X1_480/B vdd NAND2X1
XAND2X2_90 AND2X2_90/A AND2X2_90/B gnd AND2X2_90/Y vdd AND2X2
XAOI21X1_138 OR2X2_86/B OR2X2_86/A AND2X2_66/B gnd NOR2X1_125/A vdd AOI21X1
XNAND3X1_311 INVX1_215/A INVX1_213/Y INVX1_214/Y gnd AOI21X1_212/B vdd NAND3X1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XFILL_10_0_0 gnd vdd FILL
XFILL_1_2 gnd vdd FILL
XNOR2X1_362 BUFX4_13/Y INVX1_475/Y gnd NOR2X1_362/Y vdd NOR2X1
XOAI21X1_329 NOR2X1_209/Y NOR2X1_208/B AOI22X1_10/C gnd XOR2X1_188/A vdd OAI21X1
XINVX1_150 INVX1_150/A gnd INVX1_150/Y vdd INVX1
XNAND2X1_443 INVX1_305/A NOR2X1_255/Y gnd NAND3X1_373/C vdd NAND2X1
XAND2X2_54 AND2X2_54/A AND2X2_54/B gnd AND2X2_54/Y vdd AND2X2
XAOI21X1_102 OR2X2_62/B OR2X2_62/A AND2X2_48/B gnd NOR2X1_95/A vdd AOI21X1
XNAND3X1_275 INVX1_176/A NAND2X1_306/Y OR2X2_121/Y gnd NAND3X1_276/A vdd NAND3X1
XFILL_33_7_0 gnd vdd FILL
XOAI21X1_293 BUFX2_176/A NOR2X1_186/B INVX1_197/A gnd AOI22X1_8/B vdd OAI21X1
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XFILL_31_9_1 gnd vdd FILL
XNAND2X1_407 NAND3X1_347/Y INVX1_275/A gnd NAND2X1_407/Y vdd NAND2X1
XNOR2X1_326 NOR2X1_326/A NOR2X1_325/Y gnd BUFX2_237/A vdd NOR2X1
XAND2X2_18 AND2X2_18/A AND2X2_18/B gnd AND2X2_18/Y vdd AND2X2
XBUFX2_240 OR2X2_29/A gnd BUFX2_240/Y vdd BUFX2
XNOR2X1_93 NOR2X1_93/A NOR3X1_40/Y gnd NOR2X1_93/Y vdd NOR2X1
XNAND3X1_239 INVX1_154/A NAND3X1_239/B OR2X2_105/Y gnd NAND2X1_269/B vdd NAND3X1
XOAI21X1_257 AND2X2_91/Y NOR2X1_164/Y INVX1_169/A gnd NAND3X1_269/B vdd OAI21X1
XINVX2_78 INVX2_78/A gnd INVX2_78/Y vdd INVX2
XNOR2X1_290 NOR2X1_290/A NOR2X1_289/Y gnd BUFX2_225/A vdd NOR2X1
XNAND2X1_371 INVX1_235/Y NOR2X1_210/Y gnd INVX1_238/A vdd NAND2X1
XNAND3X1_203 INVX1_132/A NAND3X1_203/B OR2X2_89/Y gnd NAND2X1_231/B vdd NAND3X1
XBUFX2_204 BUFX2_204/A gnd BUFX2_204/Y vdd BUFX2
XNOR2X1_57 NOR2X1_57/A NOR2X1_57/B gnd XOR2X1_48/A vdd NOR2X1
XXNOR2X1_242 XNOR2X1_242/A NOR2X1_413/B gnd XNOR2X1_242/Y vdd XNOR2X1
XNAND2X1_335 INVX1_189/A NOR2X1_180/Y gnd AOI21X1_206/B vdd NAND2X1
XINVX2_42 INVX2_42/A gnd INVX2_42/Y vdd INVX2
XOAI21X1_221 OAI21X1_216/A XNOR2X1_115/B OAI21X1_221/C gnd OAI21X1_221/Y vdd OAI21X1
XNOR2X1_254 NOR2X1_254/A NOR2X1_254/B gnd BUFX2_213/A vdd NOR2X1
XFILL_15_2_1 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XBUFX2_168 OR2X2_117/A gnd BUFX2_168/Y vdd BUFX2
XCLKBUF1_45 BUFX4_4/Y gnd CLKBUF1_45/Y vdd CLKBUF1
XNAND3X1_167 INVX1_110/A NAND3X1_167/B OR2X2_73/Y gnd NAND3X1_170/B vdd NAND3X1
XINVX1_583 INVX1_583/A gnd INVX1_583/Y vdd INVX1
XNOR2X1_21 NOR2X1_21/A INVX2_12/A gnd XOR2X1_10/B vdd NOR2X1
XXNOR2X1_206 NOR2X1_357/Y XNOR2X1_206/B gnd XNOR2X1_206/Y vdd XNOR2X1
XOAI21X1_185 AND2X2_65/Y NOR2X1_122/Y INVX1_124/A gnd NAND3X1_193/C vdd OAI21X1
XNAND2X1_299 OR2X2_119/B OR2X2_119/A gnd NAND2X1_300/A vdd NAND2X1
XNOR2X1_218 NOR2X1_218/A NOR2X1_218/B gnd BUFX2_201/A vdd NOR2X1
XNOR3X1_98 NOR3X1_98/A NOR3X1_98/B NOR3X1_98/C gnd NOR3X1_98/Y vdd NOR3X1
XINVX1_547 bloque_bytes[78] gnd INVX1_547/Y vdd INVX1
XDFFPOSX1_365 INVX1_457/A CLKBUF1_2/Y NAND3X1_523/Y gnd vdd DFFPOSX1
XNAND3X1_131 INVX1_88/A NAND2X1_154/Y OR2X2_57/Y gnd NAND3X1_134/B vdd NAND3X1
XXNOR2X1_170 NOR2X1_249/Y XNOR2X1_170/B gnd XNOR2X1_170/Y vdd XNOR2X1
XBUFX2_132 gnd gnd BUFX2_132/Y vdd BUFX2
XOAI21X1_149 AND2X2_52/Y NOR2X1_100/Y INVX1_101/Y gnd NAND3X1_157/A vdd OAI21X1
XNOR2X1_182 NOR2X1_182/A NOR2X1_182/B gnd BUFX2_185/A vdd NOR2X1
XXNOR2X1_92 XOR2X1_101/Y XOR2X1_89/Y gnd XNOR2X1_92/Y vdd XNOR2X1
XNAND2X1_263 OR2X2_104/B OR2X2_104/A gnd NAND2X1_264/A vdd NAND2X1
XNOR3X1_62 NOR3X1_62/A INVX2_61/Y NOR3X1_62/C gnd NOR3X1_62/Y vdd NOR3X1
XINVX1_511 INVX1_511/A gnd INVX1_511/Y vdd INVX1
XDFFPOSX1_329 XNOR2X1_186/B CLKBUF1_46/Y INVX1_573/Y gnd vdd DFFPOSX1
XOAI21X1_113 NOR3X1_38/Y NOR2X1_83/A OAI21X1_113/C gnd OAI21X1_113/Y vdd OAI21X1
XXNOR2X1_56 XOR2X1_61/Y XOR2X1_49/Y gnd XNOR2X1_56/Y vdd XNOR2X1
XFILL_12_7_1 gnd vdd FILL
XXNOR2X1_134 NAND2X1_294/Y AND2X2_90/Y gnd XOR2X1_156/A vdd XNOR2X1
XFILL_14_5_0 gnd vdd FILL
XNOR2X1_146 INVX1_150/Y NOR2X1_146/B gnd NOR2X1_147/B vdd NOR2X1
XNAND2X1_227 INVX2_43/A AND2X2_66/Y gnd AOI21X1_142/C vdd NAND2X1
XNOR3X1_26 INVX1_12/Y NOR3X1_26/B AND2X2_3/Y gnd OAI21X1_9/A vdd NOR3X1
XDFFPOSX1_293 INVX1_286/A CLKBUF1_32/Y AOI21X1_382/C gnd vdd DFFPOSX1
XINVX1_475 INVX1_475/A gnd INVX1_475/Y vdd INVX1
XFILL_24_0_0 gnd vdd FILL
XXOR2X1_290 BUFX2_245/A gnd gnd INVX2_91/A vdd XOR2X1
XXNOR2X1_20 XOR2X1_21/Y XOR2X1_9/Y gnd XNOR2X1_21/A vdd XNOR2X1
XFILL_4_1_0 gnd vdd FILL
XFILL_22_2_1 gnd vdd FILL
XNOR2X1_110 gnd OR2X2_75/B gnd NOR2X1_110/Y vdd NOR2X1
XFILL_2_3_1 gnd vdd FILL
XNAND2X1_191 INVX2_38/Y XNOR2X1_85/Y gnd XNOR2X1_87/B vdd NAND2X1
XAOI21X1_89 AOI21X1_89/A AOI21X1_89/B AOI21X1_89/C gnd AOI21X1_89/Y vdd AOI21X1
XDFFPOSX1_257 XNOR2X1_150/B CLKBUF1_47/Y OR2X2_144/A gnd vdd DFFPOSX1
XOAI21X1_618 AND2X2_181/Y NOR2X1_421/Y INVX1_520/A gnd OR2X2_138/A vdd OAI21X1
XOR2X2_78 OR2X2_78/A OR2X2_78/B gnd OR2X2_78/Y vdd OR2X2
XINVX1_439 INVX1_439/A gnd INVX1_439/Y vdd INVX1
XXOR2X1_254 BUFX2_225/A gnd gnd XOR2X1_254/Y vdd XOR2X1
XBUFX2_92 gnd gnd BUFX2_92/Y vdd BUFX2
XAOI21X1_391 XNOR2X1_215/Y NOR2X1_411/Y INVX1_510/Y gnd OAI21X1_627/B vdd AOI21X1
XNAND2X1_155 NAND3X1_132/B NAND3X1_134/B gnd XNOR2X1_69/A vdd NAND2X1
XAOI21X1_53 AOI21X1_53/A AOI21X1_53/B OAI21X1_69/B gnd AOI21X1_53/Y vdd AOI21X1
XOAI21X1_582 AND2X2_173/Y INVX1_481/A BUFX4_30/Y gnd OAI21X1_582/Y vdd OAI21X1
XOR2X2_42 gnd OR2X2_42/B gnd OR2X2_42/Y vdd OR2X2
XDFFPOSX1_221 INVX1_145/A CLKBUF1_36/Y INVX1_503/A gnd vdd DFFPOSX1
XINVX1_403 BUFX2_223/A gnd INVX1_403/Y vdd INVX1
XBUFX2_56 gnd gnd BUFX2_56/Y vdd BUFX2
XXOR2X1_218 BUFX2_209/A gnd gnd NOR2X1_264/B vdd XOR2X1
XNAND2X1_696 INVX2_91/A NOR2X1_440/B gnd OAI21X1_631/A vdd NAND2X1
XNAND2X1_119 NAND3X1_98/Y OAI21X1_94/Y gnd XNOR2X1_52/A vdd NAND2X1
XAOI21X1_355 bloque_bytes[69] INVX1_498/Y INVX1_574/A gnd OAI21X1_594/C vdd AOI21X1
XFILL_21_5_0 gnd vdd FILL
XOAI21X1_6 INVX2_10/Y target[3] NOR2X1_15/A gnd OAI21X1_7/C vdd OAI21X1
XNAND3X1_528 BUFX2_244/A BUFX2_245/A AND2X2_189/A gnd XOR2X1_307/A vdd NAND3X1
XFILL_1_6_0 gnd vdd FILL
XAOI21X1_17 AOI21X1_17/A AOI21X1_17/B OAI21X1_18/B gnd NAND3X1_20/B vdd AOI21X1
XDFFPOSX1_185 XOR2X1_81/B CLKBUF1_12/Y bloque_bytes[31] gnd vdd DFFPOSX1
XFILL_19_7_1 gnd vdd FILL
XXOR2X1_182 BUFX2_189/A gnd gnd XOR2X1_182/Y vdd XOR2X1
XINVX1_367 INVX1_367/A gnd INVX1_367/Y vdd INVX1
XOAI21X1_546 gnd XOR2X1_279/Y INVX1_453/A gnd OAI21X1_546/Y vdd OAI21X1
XFILL_14_2 gnd vdd FILL
XNAND2X1_660 XNOR2X1_217/Y AOI21X1_393/B gnd NOR2X1_434/B vdd NAND2X1
XBUFX2_20 BUFX2_20/A gnd hash[19] vdd BUFX2
XNAND2X1_80 gnd OR2X2_26/B gnd NAND2X1_80/Y vdd NAND2X1
XOAI21X1_65 AND2X2_22/Y NOR2X1_50/Y INVX1_46/A gnd AOI21X1_49/A vdd OAI21X1
XDFFPOSX1_83 INVX2_79/A CLKBUF1_14/Y AND2X2_175/Y gnd vdd DFFPOSX1
XNAND3X1_492 AND2X2_163/B INVX1_477/A INVX1_488/Y gnd NOR2X1_394/A vdd NAND3X1
XAOI21X1_319 NAND3X1_477/Y AOI21X1_319/B INVX1_465/Y gnd AOI21X1_320/A vdd AOI21X1
XFILL_31_0_0 gnd vdd FILL
XFILL_29_2_1 gnd vdd FILL
XDFFPOSX1_149 INVX1_46/A CLKBUF1_29/Y bloque_bytes[59] gnd vdd DFFPOSX1
XFILL_9_3_1 gnd vdd FILL
XOAI21X1_510 NOR3X1_82/C INVX2_71/Y NOR3X1_82/A gnd AND2X2_148/A vdd OAI21X1
XINVX1_331 INVX1_331/A gnd INVX1_331/Y vdd INVX1
XNAND2X1_624 AND2X2_166/B AND2X2_171/Y gnd NAND2X1_624/Y vdd NAND2X1
XXOR2X1_146 XOR2X1_146/A AND2X2_89/A gnd OR2X2_124/B vdd XOR2X1
XAOI21X1_283 INVX1_388/A NAND3X1_429/B INVX1_383/Y gnd NOR2X1_304/B vdd AOI21X1
XOAI21X1_29 OAI21X1_29/A XNOR2X1_16/B INVX1_30/A gnd XOR2X1_20/A vdd OAI21X1
XNAND2X1_44 INVX1_30/A OAI21X1_28/Y gnd OAI21X1_29/A vdd NAND2X1
XDFFPOSX1_47 INVX1_533/A CLKBUF1_26/Y NOR2X1_370/Y gnd vdd DFFPOSX1
XDFFPOSX1_113 INVX1_5/A CLKBUF1_35/Y XOR2X1_308/Y gnd vdd DFFPOSX1
XNAND3X1_456 INVX1_426/A NAND3X1_456/B NAND2X1_560/Y gnd NAND2X1_562/A vdd NAND3X1
XXOR2X1_90 XOR2X1_90/A XOR2X1_90/B gnd XOR2X1_90/Y vdd XOR2X1
XXOR2X1_110 XOR2X1_110/A XOR2X1_110/B gnd BUFX2_162/A vdd XOR2X1
XINVX1_295 INVX1_295/A gnd INVX1_295/Y vdd INVX1
XOAI21X1_474 NOR3X1_77/A INVX1_380/A OAI21X1_474/C gnd NOR2X1_302/A vdd OAI21X1
XNAND2X1_588 NAND2X1_588/A AOI22X1_21/C gnd NAND2X1_588/Y vdd NAND2X1
XAOI21X1_247 NAND3X1_360/Y AOI21X1_247/B INVX1_294/Y gnd AOI21X1_247/Y vdd AOI21X1
XNAND3X1_420 INVX1_364/A NAND3X1_420/B NAND3X1_420/C gnd NAND2X1_512/A vdd NAND3X1
XAOI22X1_22 INVX1_466/A AOI22X1_22/B AOI22X1_22/C INVX1_464/A gnd INVX1_470/A vdd
+ AOI22X1
XINVX1_259 INVX1_259/A gnd INVX1_259/Y vdd INVX1
XDFFPOSX1_11 BUFX2_10/A CLKBUF1_41/Y NOR3X1_10/Y gnd vdd DFFPOSX1
XNAND3X1_85 NAND3X1_85/A NAND3X1_84/Y NAND3X1_85/C gnd AND2X2_30/B vdd NAND3X1
XXOR2X1_54 XOR2X1_54/A gnd gnd OR2X2_50/B vdd XOR2X1
XNAND2X1_552 INVX1_415/Y AND2X2_146/A gnd NAND3X1_449/B vdd NAND2X1
XOAI21X1_438 gnd NOR2X1_279/B INVX1_343/Y gnd OAI21X1_438/Y vdd OAI21X1
XAND2X2_190 INVX1_584/A XOR2X1_289/Y gnd NOR2X1_440/B vdd AND2X2
XFILL_28_5_0 gnd vdd FILL
XFILL_6_8_1 gnd vdd FILL
XFILL_8_6_0 gnd vdd FILL
XOR2X2_137 OR2X2_137/A bloque_bytes[11] gnd OR2X2_137/Y vdd OR2X2
XFILL_26_7_1 gnd vdd FILL
XAOI21X1_211 INVX1_217/A NAND3X1_312/B INVX1_212/Y gnd NOR2X1_196/B vdd AOI21X1
XNAND3X1_384 INVX2_66/A NAND3X1_384/B NAND3X1_384/C gnd NOR3X1_71/A vdd NAND3X1
XINVX1_223 INVX1_223/A gnd INVX1_223/Y vdd INVX1
XMUX2X1_7 BUFX2_7/A MUX2X1_7/B BUFX4_8/Y gnd MUX2X1_7/Y vdd MUX2X1
XAND2X2_154 NOR2X1_346/Y INVX1_453/Y gnd NOR3X1_86/A vdd AND2X2
XOAI21X1_402 BUFX2_203/A INVX1_309/A INVX1_310/A gnd INVX1_312/A vdd OAI21X1
XNAND3X1_49 AOI21X1_36/A NAND3X1_49/B NAND3X1_49/C gnd AND2X2_18/B vdd NAND3X1
XXOR2X1_18 XOR2X1_18/A XOR2X1_4/A gnd XOR2X1_18/Y vdd XOR2X1
XOR2X2_101 OR2X2_101/A OR2X2_101/B gnd OR2X2_101/Y vdd OR2X2
XFILL_36_2_1 gnd vdd FILL
XNAND2X1_516 INVX1_378/Y NOR2X1_299/Y gnd NAND3X1_423/C vdd NAND2X1
XNOR2X1_435 gnd gnd gnd NOR2X1_435/Y vdd NOR2X1
XAOI21X1_175 NOR2X1_155/Y AOI21X1_175/B INVX1_161/A gnd NOR2X1_157/A vdd AOI21X1
XNAND3X1_348 INVX1_269/A AOI21X1_237/B INVX1_268/Y gnd INVX1_275/A vdd NAND3X1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XNOR2X1_399 INVX1_491/A INVX2_82/A gnd INVX2_83/A vdd NOR2X1
XINVX1_187 INVX1_187/A gnd AND2X2_98/B vdd INVX1
XCLKBUF1_8 BUFX4_5/Y gnd CLKBUF1_8/Y vdd CLKBUF1
XAND2X2_118 NOR2X1_238/Y INVX1_282/Y gnd NOR3X1_68/A vdd AND2X2
XOAI21X1_366 NOR3X1_65/C OAI21X1_366/B INVX1_275/A gnd NOR2X1_233/A vdd OAI21X1
XNAND3X1_13 AOI21X1_12/A NAND3X1_12/Y OAI21X1_15/Y gnd AND2X2_6/B vdd NAND3X1
XNAND2X1_480 INVX1_344/A NAND2X1_480/B gnd INVX1_342/A vdd NAND2X1
XAND2X2_91 OR2X2_117/A OR2X2_117/B gnd AND2X2_91/Y vdd AND2X2
XAOI21X1_139 NOR2X1_125/Y AOI21X1_139/B INVX1_128/A gnd NOR2X1_127/A vdd AOI21X1
XNAND3X1_312 INVX1_217/A NAND3X1_312/B INVX1_212/Y gnd AOI22X1_9/C vdd NAND3X1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XFILL_10_0_1 gnd vdd FILL
XOAI21X1_330 BUFX2_184/A NOR2X1_210/B INVX1_235/Y gnd NAND3X1_326/B vdd OAI21X1
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XNOR2X1_363 BUFX4_16/Y INVX1_476/Y gnd NOR2X1_363/Y vdd NOR2X1
XNAND2X1_444 INVX1_305/Y NOR2X1_255/Y gnd AOI21X1_253/B vdd NAND2X1
XAOI21X1_103 NOR2X1_95/Y AOI21X1_103/B INVX1_95/A gnd NOR2X1_97/A vdd AOI21X1
XAND2X2_55 OR2X2_69/A OR2X2_69/B gnd AND2X2_55/Y vdd AND2X2
XNAND3X1_276 NAND3X1_276/A OAI21X1_263/Y NAND3X1_276/C gnd XNOR2X1_142/B vdd NAND3X1
XFILL_35_5_0 gnd vdd FILL
XFILL_33_7_1 gnd vdd FILL
XOAI21X1_294 gnd NOR2X1_180/B INVX1_189/Y gnd AOI21X1_206/A vdd OAI21X1
XINVX1_115 OR2X2_78/Y gnd INVX1_115/Y vdd INVX1
XNAND2X1_408 INVX1_273/A NOR2X1_234/Y gnd NAND3X1_352/C vdd NAND2X1
XNOR2X1_327 gnd NOR2X1_327/B gnd NOR2X1_327/Y vdd NOR2X1
XAND2X2_19 OR2X2_21/A OR2X2_21/B gnd AND2X2_19/Y vdd AND2X2
XNAND3X1_240 NAND2X1_269/B NAND2X1_269/A XNOR2X1_123/B gnd NAND3X1_240/Y vdd NAND3X1
XBUFX2_241 BUFX2_241/A gnd BUFX2_241/Y vdd BUFX2
XNOR2X1_94 OR2X2_61/A OR2X2_61/B gnd NOR2X1_94/Y vdd NOR2X1
XOAI21X1_258 AND2X2_91/Y NOR2X1_164/Y INVX1_169/Y gnd NAND3X1_271/A vdd OAI21X1
XINVX2_79 INVX2_79/A gnd INVX2_79/Y vdd INVX2
XNOR2X1_291 gnd NOR2X1_291/B gnd NOR2X1_291/Y vdd NOR2X1
XNAND2X1_372 NAND2X1_372/A NAND2X1_372/B gnd XOR2X1_188/B vdd NAND2X1
XNAND3X1_204 NAND2X1_231/B NAND2X1_231/A XNOR2X1_105/B gnd XNOR2X1_106/B vdd NAND3X1
XBUFX2_205 BUFX2_205/A gnd BUFX2_205/Y vdd BUFX2
XNOR2X1_58 gnd OR2X2_33/B gnd NOR2X1_58/Y vdd NOR2X1
XOAI21X1_222 XNOR2X1_116/A OAI21X1_222/B AND2X2_78/B gnd XNOR2X1_117/A vdd OAI21X1
XXNOR2X1_243 INVX1_579/A gnd gnd XNOR2X1_243/Y vdd XNOR2X1
XNAND2X1_336 XOR2X1_170/B NOR2X1_184/Y gnd AOI21X1_208/C vdd NAND2X1
XINVX2_43 INVX2_43/A gnd INVX2_43/Y vdd INVX2
XFILL_17_0_1 gnd vdd FILL
XNOR2X1_255 gnd XOR2X1_210/Y gnd NOR2X1_255/Y vdd NOR2X1
XNOR2X1_22 gnd OR2X2_4/B gnd NOR2X1_22/Y vdd NOR2X1
XBUFX2_169 BUFX2_169/A gnd BUFX2_169/Y vdd BUFX2
XNAND3X1_168 NAND3X1_170/B OAI21X1_161/Y XNOR2X1_87/B gnd XNOR2X1_88/B vdd NAND3X1
XINVX1_584 INVX1_584/A gnd INVX1_584/Y vdd INVX1
XXNOR2X1_207 XNOR2X1_206/Y OAI21X1_561/Y gnd INVX1_471/A vdd XNOR2X1
XCLKBUF1_46 BUFX4_5/Y gnd CLKBUF1_46/Y vdd CLKBUF1
XOAI21X1_186 AND2X2_65/Y NOR2X1_122/Y INVX1_124/Y gnd NAND3X1_197/A vdd OAI21X1
XNOR2X1_219 gnd XOR2X1_183/Y gnd NOR2X1_219/Y vdd NOR2X1
XNAND2X1_300 NAND2X1_300/A OR2X2_119/Y gnd OR2X2_120/A vdd NAND2X1
XBUFX2_133 gnd gnd BUFX2_133/Y vdd BUFX2
XINVX1_548 INVX1_548/A gnd INVX1_548/Y vdd INVX1
XCLKBUF1_10 BUFX4_3/Y gnd CLKBUF1_10/Y vdd CLKBUF1
XNAND3X1_132 NAND3X1_134/B NAND3X1_132/B XNOR2X1_69/B gnd XNOR2X1_70/B vdd NAND3X1
XDFFPOSX1_366 INVX1_462/A CLKBUF1_51/Y NAND3X1_524/Y gnd vdd DFFPOSX1
XXNOR2X1_93 XNOR2X1_92/Y OR2X2_79/Y gnd INVX1_120/A vdd XNOR2X1
XXNOR2X1_171 XNOR2X1_170/Y OAI21X1_390/Y gnd INVX1_300/A vdd XNOR2X1
XOAI21X1_150 AND2X2_52/Y NOR2X1_100/Y INVX1_101/A gnd AOI21X1_109/A vdd OAI21X1
XNOR2X1_183 gnd NOR2X1_183/B gnd NOR2X1_183/Y vdd NOR2X1
XNAND2X1_264 NAND2X1_264/A OR2X2_104/Y gnd INVX1_150/A vdd NAND2X1
XNOR3X1_63 NOR3X1_63/A INVX1_247/A NOR3X1_63/C gnd NOR3X1_63/Y vdd NOR3X1
XDFFPOSX1_330 INVX1_377/A CLKBUF1_51/Y OR2X2_145/Y gnd vdd DFFPOSX1
XFILL_27_1 gnd vdd FILL
XINVX1_512 bloque_bytes[58] gnd INVX1_512/Y vdd INVX1
XFILL_16_3_0 gnd vdd FILL
XXNOR2X1_57 XNOR2X1_56/Y OR2X2_47/Y gnd INVX1_76/A vdd XNOR2X1
XOAI21X1_114 OAI21X1_119/A XNOR2X1_61/B INVX1_85/A gnd XOR2X1_70/A vdd OAI21X1
XXNOR2X1_135 OAI21X1_256/Y INVX2_55/Y gnd XOR2X1_157/A vdd XNOR2X1
XFILL_14_5_1 gnd vdd FILL
XNAND2X1_228 NAND2X1_228/A OAI21X1_194/Y gnd XOR2X1_119/A vdd NAND2X1
XNOR2X1_147 NOR2X1_147/A NOR2X1_147/B gnd XOR2X1_138/A vdd NOR2X1
XNOR3X1_27 INVX1_22/Y NOR2X1_28/Y AND2X2_8/Y gnd NOR3X1_27/Y vdd NOR3X1
XDFFPOSX1_294 INVX1_291/A CLKBUF1_23/Y XNOR2X1_242/A gnd vdd DFFPOSX1
XINVX1_476 INVX1_476/A gnd INVX1_476/Y vdd INVX1
XFILL_24_0_1 gnd vdd FILL
XXOR2X1_291 BUFX2_246/A gnd gnd INVX1_581/A vdd XOR2X1
XXNOR2X1_21 XNOR2X1_21/A OR2X2_15/Y gnd INVX1_32/A vdd XNOR2X1
XFILL_4_1_1 gnd vdd FILL
XNOR2X1_111 NOR2X1_111/A INVX2_39/A gnd XOR2X1_100/B vdd NOR2X1
XNAND2X1_192 gnd OR2X2_73/B gnd NAND3X1_167/B vdd NAND2X1
XAOI21X1_90 OR2X2_54/B OR2X2_54/A AND2X2_42/B gnd NOR2X1_85/A vdd AOI21X1
XOAI21X1_619 NOR2X1_422/Y NOR2X1_423/Y INVX1_523/A gnd NOR2X1_428/B vdd OAI21X1
XOR2X2_79 OR2X2_79/A OR2X2_79/B gnd OR2X2_79/Y vdd OR2X2
XDFFPOSX1_258 INVX1_206/A CLKBUF1_32/Y INVX1_508/Y gnd vdd DFFPOSX1
XINVX1_440 INVX1_440/A gnd INVX1_440/Y vdd INVX1
XBUFX2_93 gnd gnd BUFX2_93/Y vdd BUFX2
XXOR2X1_255 BUFX2_226/A gnd gnd XOR2X1_255/Y vdd XOR2X1
XFILL_13_8_0 gnd vdd FILL
XAOI21X1_392 XNOR2X1_216/Y NAND2X1_659/B INVX1_513/Y gnd OAI21X1_628/B vdd AOI21X1
XNAND2X1_156 gnd OR2X2_58/B gnd AOI21X1_95/A vdd NAND2X1
XAOI21X1_54 OR2X2_30/B OR2X2_30/A AND2X2_24/B gnd NOR2X1_55/A vdd AOI21X1
XDFFPOSX1_222 INVX1_146/A CLKBUF1_50/Y INVX1_504/A gnd vdd DFFPOSX1
XOAI21X1_583 OAI21X1_583/A INVX1_481/Y INVX1_482/A gnd OAI21X1_583/Y vdd OAI21X1
XOR2X2_43 gnd OR2X2_43/B gnd OR2X2_43/Y vdd OR2X2
XXOR2X1_219 BUFX2_210/A gnd gnd NOR2X1_267/B vdd XOR2X1
XINVX1_404 INVX1_404/A gnd INVX1_404/Y vdd INVX1
XNAND2X1_697 INVX1_585/A NOR2X1_350/Y gnd NAND2X1_698/A vdd NAND2X1
XBUFX2_57 gnd gnd BUFX2_57/Y vdd BUFX2
XAOI21X1_356 bloque_bytes[70] INVX1_499/Y INVX1_575/A gnd OAI21X1_595/C vdd AOI21X1
XNAND2X1_120 INVX1_74/A OAI21X1_96/Y gnd OAI21X1_97/A vdd NAND2X1
XFILL_21_5_1 gnd vdd FILL
XFILL_23_3_0 gnd vdd FILL
XOAI21X1_7 OAI21X1_7/A AOI21X1_6/Y OAI21X1_7/C gnd OAI21X1_7/Y vdd OAI21X1
XNAND3X1_529 INVX1_582/A NOR2X1_440/B NOR2X1_441/Y gnd AND2X2_191/B vdd NAND3X1
XFILL_1_6_1 gnd vdd FILL
XFILL_3_4_0 gnd vdd FILL
XAOI21X1_18 OR2X2_6/B OR2X2_6/A AND2X2_6/B gnd NOR2X1_25/A vdd AOI21X1
XDFFPOSX1_186 INVX2_35/A CLKBUF1_49/Y bloque_bytes[16] gnd vdd DFFPOSX1
XINVX1_368 INVX1_368/A gnd INVX1_368/Y vdd INVX1
XXOR2X1_183 BUFX2_190/A gnd gnd XOR2X1_183/Y vdd XOR2X1
XNAND2X1_661 bloque_bytes[0] OR2X2_150/B gnd AOI21X1_379/B vdd NAND2X1
XOAI21X1_547 gnd NOR2X1_347/B INVX1_454/A gnd INVX2_73/A vdd OAI21X1
XBUFX2_21 BUFX2_21/A gnd hash[20] vdd BUFX2
XFILL_31_0_1 gnd vdd FILL
XAOI21X1_320 AOI21X1_320/A AOI21X1_320/B NAND2X1_602/Y gnd AOI21X1_320/Y vdd AOI21X1
XOAI21X1_66 AND2X2_23/Y NOR2X1_52/Y INVX1_47/A gnd NAND3X1_67/C vdd OAI21X1
XNAND2X1_81 NAND2X1_81/A NAND2X1_81/B gnd NAND3X1_75/B vdd NAND2X1
XDFFPOSX1_84 AND2X2_167/B CLKBUF1_6/Y NOR2X1_405/Y gnd vdd DFFPOSX1
XNAND3X1_493 AND2X2_162/B AND2X2_163/B INVX1_477/A gnd INVX1_489/A vdd NAND3X1
XDFFPOSX1_150 INVX1_47/A CLKBUF1_29/Y bloque_bytes[60] gnd vdd DFFPOSX1
XINVX1_332 INVX1_332/A gnd INVX1_332/Y vdd INVX1
XOAI21X1_511 gnd NOR2X1_324/B INVX1_417/A gnd INVX1_420/A vdd OAI21X1
XNAND2X1_625 AND2X2_166/B INVX1_479/A gnd NOR2X1_402/A vdd NAND2X1
XXOR2X1_147 XOR2X1_147/A OR2X2_117/A gnd OR2X2_125/B vdd XOR2X1
XNAND2X1_45 gnd OR2X2_11/B gnd NAND3X1_28/B vdd NAND2X1
XAOI21X1_284 OAI21X1_479/Y NAND3X1_433/C INVX1_383/A gnd NOR2X1_304/A vdd AOI21X1
XNAND3X1_457 AOI22X1_20/B INVX1_428/A INVX1_426/Y gnd NAND2X1_562/B vdd NAND3X1
XDFFPOSX1_114 INVX2_92/A CLKBUF1_5/Y bloque_bytes[88] gnd vdd DFFPOSX1
XOAI21X1_30 AND2X2_10/Y NOR2X1_30/Y INVX1_24/Y gnd AOI21X1_24/A vdd OAI21X1
XDFFPOSX1_48 INVX1_548/A CLKBUF1_15/Y NOR2X1_371/Y gnd vdd DFFPOSX1
XXOR2X1_91 XOR2X1_75/A XOR2X1_91/B gnd XOR2X1_91/Y vdd XOR2X1
XXOR2X1_111 XOR2X1_90/Y XOR2X1_111/B gnd XOR2X1_111/Y vdd XOR2X1
XFILL_20_8_0 gnd vdd FILL
XINVX1_296 INVX1_296/A gnd INVX1_296/Y vdd INVX1
XOAI21X1_475 NOR3X1_78/A NOR3X1_78/C INVX2_69/A gnd NOR2X1_301/A vdd OAI21X1
XFILL_0_9_0 gnd vdd FILL
XNAND2X1_589 NAND2X1_589/A NAND2X1_589/B gnd XOR2X1_295/A vdd NAND2X1
XAOI21X1_248 AOI21X1_247/Y AOI21X1_248/B NAND2X1_431/Y gnd OAI21X1_391/A vdd AOI21X1
XDFFPOSX1_12 BUFX2_11/A CLKBUF1_48/Y NOR3X1_11/Y gnd vdd DFFPOSX1
XNAND3X1_421 INVX1_375/Y INVX1_374/A AOI21X1_282/B gnd AND2X2_137/B vdd NAND3X1
XINVX1_260 INVX1_260/A gnd INVX1_260/Y vdd INVX1
XFILL_30_3_0 gnd vdd FILL
XOAI21X1_439 gnd NOR2X1_279/B INVX1_343/A gnd INVX1_345/A vdd OAI21X1
XXOR2X1_55 XOR2X1_71/A gnd gnd OR2X2_51/B vdd XOR2X1
XNAND3X1_86 INVX1_58/A NAND3X1_84/B OR2X2_36/Y gnd NAND3X1_87/B vdd NAND3X1
XOR2X2_138 OR2X2_138/A bloque_bytes[12] gnd OR2X2_138/Y vdd OR2X2
XNAND2X1_553 NAND2X1_553/A NAND3X1_449/B gnd INVX1_460/A vdd NAND2X1
XAND2X2_191 AND2X2_191/A AND2X2_191/B gnd AND2X2_191/Y vdd AND2X2
XFILL_28_5_1 gnd vdd FILL
XFILL_8_6_1 gnd vdd FILL
XAOI21X1_212 AOI21X1_212/A AOI21X1_212/B INVX1_212/A gnd NOR2X1_196/A vdd AOI21X1
XMUX2X1_8 BUFX2_8/A MUX2X1_8/B MUX2X1_8/S gnd NOR3X1_8/B vdd MUX2X1
XNAND3X1_385 INVX1_325/A NAND2X1_460/Y INVX2_66/Y gnd OAI21X1_423/B vdd NAND3X1
XINVX1_224 INVX1_224/A gnd INVX1_224/Y vdd INVX1
XOAI21X1_403 BUFX2_203/A INVX1_309/A INVX1_310/Y gnd OAI21X1_403/Y vdd OAI21X1
XNOR2X1_436 NOR2X1_435/Y INVX1_579/Y gnd NOR2X1_436/Y vdd NOR2X1
XAND2X2_155 NOR2X1_347/Y INVX1_454/Y gnd NOR3X1_86/C vdd AND2X2
XXOR2X1_19 XOR2X1_19/A XOR2X1_5/A gnd XOR2X1_19/Y vdd XOR2X1
XNAND3X1_50 INVX1_36/A NAND3X1_50/B OR2X2_20/Y gnd NAND3X1_51/B vdd NAND3X1
XOR2X2_102 OR2X2_102/A OR2X2_102/B gnd INVX1_148/A vdd OR2X2
XNAND2X1_517 INVX1_379/Y NOR2X1_300/Y gnd NAND2X1_517/Y vdd NAND2X1
XAOI21X1_176 INVX2_51/Y INVX1_162/Y NOR2X1_151/A gnd AOI21X1_178/A vdd AOI21X1
XNAND3X1_349 INVX1_270/Y INVX1_271/Y INVX1_272/Y gnd AOI21X1_235/B vdd NAND3X1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XINVX1_188 INVX1_188/A gnd AND2X2_99/B vdd INVX1
XNAND3X1_14 INVX1_14/A NAND3X1_14/B OR2X2_4/Y gnd NAND3X1_15/B vdd NAND3X1
XCLKBUF1_9 BUFX4_6/Y gnd CLKBUF1_9/Y vdd CLKBUF1
XNOR2X1_400 INVX2_75/Y INVX2_76/Y gnd NOR2X1_400/Y vdd NOR2X1
XOAI21X1_367 NOR2X1_233/Y NOR2X1_232/B AOI22X1_12/C gnd XOR2X1_206/A vdd OAI21X1
XAND2X2_119 NOR2X1_239/Y INVX1_283/Y gnd NOR3X1_68/C vdd AND2X2
XNAND2X1_481 INVX1_343/A NOR2X1_279/Y gnd NAND3X1_399/C vdd NAND2X1
XFILL_7_9_0 gnd vdd FILL
XAOI21X1_140 INVX2_42/Y INVX1_129/Y NOR2X1_121/A gnd AOI21X1_140/Y vdd AOI21X1
XNAND3X1_313 INVX1_217/A NAND3X1_313/B NAND3X1_313/C gnd AOI21X1_217/A vdd NAND3X1
XAND2X2_92 gnd AND2X2_92/B gnd NOR3X1_55/C vdd AND2X2
XFILL_27_8_0 gnd vdd FILL
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XOAI21X1_331 BUFX2_184/A NOR2X1_210/B INVX1_235/A gnd AOI22X1_10/B vdd OAI21X1
XINVX1_152 OR2X2_104/Y gnd INVX1_152/Y vdd INVX1
XNOR2X1_364 BUFX4_14/Y INVX1_477/Y gnd NOR2X1_364/Y vdd NOR2X1
XNAND2X1_445 AOI21X1_255/A INVX1_313/A gnd NAND2X1_445/Y vdd NAND2X1
XAOI21X1_104 INVX2_33/Y INVX1_96/Y NOR2X1_91/A gnd AOI21X1_106/A vdd AOI21X1
XAND2X2_56 gnd OR2X2_73/B gnd AND2X2_56/Y vdd AND2X2
XFILL_35_5_1 gnd vdd FILL
XNAND3X1_277 INVX1_177/A AOI21X1_191/A OR2X2_122/Y gnd NAND3X1_279/A vdd NAND3X1
XOAI21X1_295 BUFX2_177/A NOR2X1_187/B INVX1_201/A gnd XNOR2X1_151/B vdd OAI21X1
XINVX1_116 INVX1_116/A gnd OR2X2_79/B vdd INVX1
XNOR2X1_328 NOR2X1_328/A NOR2X1_328/B gnd NOR2X1_328/Y vdd NOR2X1
XNAND2X1_409 INVX1_273/Y NOR2X1_234/Y gnd INVX1_276/A vdd NAND2X1
XBUFX2_242 XOR2X1_39/B gnd BUFX2_242/Y vdd BUFX2
XAND2X2_20 gnd OR2X2_25/B gnd NOR3X1_31/C vdd AND2X2
XNAND3X1_241 INVX1_155/A AOI21X1_167/A OR2X2_106/Y gnd NAND3X1_242/C vdd NAND3X1
XOAI21X1_259 NAND2X1_294/Y AOI21X1_190/C NOR2X1_165/Y gnd NOR2X1_166/B vdd OAI21X1
XNOR2X1_95 NOR2X1_95/A INVX1_93/Y gnd NOR2X1_95/Y vdd NOR2X1
XINVX2_80 INVX2_80/A gnd INVX2_80/Y vdd INVX2
XFILL_11_1_0 gnd vdd FILL
XNAND2X1_373 INVX1_227/A NOR2X1_204/Y gnd NAND2X1_373/Y vdd NAND2X1
XNOR2X1_292 NOR2X1_292/A NOR2X1_292/B gnd NOR2X1_292/Y vdd NOR2X1
XNAND3X1_205 INVX1_133/A NAND2X1_232/Y OR2X2_90/Y gnd NAND3X1_206/C vdd NAND3X1
XBUFX2_206 BUFX2_206/A gnd BUFX2_206/Y vdd BUFX2
XNOR2X1_59 gnd OR2X2_34/B gnd NOR3X1_34/B vdd NOR2X1
XOAI21X1_223 AND2X2_79/Y NOR2X1_144/Y INVX1_147/A gnd NAND3X1_233/B vdd OAI21X1
XFILL_34_8_0 gnd vdd FILL
XXNOR2X1_244 XNOR2X1_244/A INVX2_90/Y gnd XNOR2X1_244/Y vdd XNOR2X1
XNAND2X1_337 INVX1_201/Y NOR2X1_187/Y gnd NAND2X1_338/B vdd NAND2X1
XINVX2_44 INVX2_44/A gnd INVX2_44/Y vdd INVX2
XNOR2X1_256 NOR2X1_256/A NOR2X1_256/B gnd NOR2X1_256/Y vdd NOR2X1
XINVX1_585 INVX1_585/A gnd INVX1_585/Y vdd INVX1
XNAND3X1_169 INVX1_111/A NAND3X1_169/B OR2X2_74/Y gnd AOI21X1_120/C vdd NAND3X1
XNOR2X1_23 OAI21X1_9/B OAI21X1_9/A gnd NOR2X1_23/Y vdd NOR2X1
XCLKBUF1_47 BUFX4_6/Y gnd CLKBUF1_47/Y vdd CLKBUF1
XBUFX2_170 BUFX2_170/A gnd BUFX2_170/Y vdd BUFX2
XXNOR2X1_208 bloque_bytes[48] bloque_bytes[8] gnd XNOR2X1_208/Y vdd XNOR2X1
XOAI21X1_187 OAI21X1_182/A XNOR2X1_97/B OAI21X1_187/C gnd NAND3X1_200/C vdd OAI21X1
XNOR2X1_220 NOR2X1_220/A NOR2X1_220/B gnd NOR2X1_220/Y vdd NOR2X1
XNAND2X1_301 OR2X2_120/B OR2X2_120/A gnd NAND2X1_302/A vdd NAND2X1
XFILL_5_1 gnd vdd FILL
XBUFX2_134 gnd gnd BUFX2_134/Y vdd BUFX2
XINVX1_549 INVX1_549/A gnd INVX1_549/Y vdd INVX1
XCLKBUF1_11 BUFX4_1/Y gnd CLKBUF1_11/Y vdd CLKBUF1
XNAND3X1_133 INVX1_89/A AOI21X1_95/A OR2X2_58/Y gnd AOI21X1_96/C vdd NAND3X1
XDFFPOSX1_367 INVX1_463/A CLKBUF1_22/Y NAND3X1_525/Y gnd vdd DFFPOSX1
XOAI21X1_151 AND2X2_53/Y NOR2X1_102/Y INVX1_102/A gnd OAI21X1_151/Y vdd OAI21X1
XXNOR2X1_94 gnd XOR2X1_92/Y gnd XNOR2X1_94/Y vdd XNOR2X1
XXNOR2X1_172 NOR2X1_254/A NAND2X1_445/Y gnd BUFX2_214/A vdd XNOR2X1
XNOR2X1_184 NOR2X1_184/A NOR2X1_184/B gnd NOR2X1_184/Y vdd NOR2X1
XNAND2X1_265 INVX2_49/A AND2X2_78/Y gnd AOI21X1_166/C vdd NAND2X1
XFILL_18_1_0 gnd vdd FILL
XNOR3X1_64 NOR3X1_64/A INVX2_62/Y NOR3X1_64/C gnd NOR3X1_64/Y vdd NOR3X1
XFILL_27_2 gnd vdd FILL
XDFFPOSX1_331 INVX1_378/A CLKBUF1_45/Y OR2X2_146/Y gnd vdd DFFPOSX1
XXNOR2X1_136 BUFX2_169/A XOR2X1_138/Y gnd OR2X2_119/A vdd XNOR2X1
XFILL_16_3_1 gnd vdd FILL
XINVX1_513 INVX1_513/A gnd INVX1_513/Y vdd INVX1
XOAI21X1_115 AND2X2_40/Y NOR2X1_80/Y INVX1_79/Y gnd AOI21X1_84/A vdd OAI21X1
XXNOR2X1_58 gnd XOR2X1_52/Y gnd AOI21X1_93/B vdd XNOR2X1
XNOR2X1_148 gnd OR2X2_105/B gnd NOR3X1_51/B vdd NOR2X1
XNAND2X1_229 INVX2_44/Y XNOR2X1_104/A gnd XNOR2X1_105/B vdd NAND2X1
XNOR3X1_28 INVX1_23/Y NOR3X1_28/B AND2X2_9/Y gnd NOR2X1_33/B vdd NOR3X1
XINVX1_477 INVX1_477/A gnd INVX1_477/Y vdd INVX1
XDFFPOSX1_295 INVX1_292/A CLKBUF1_32/Y INVX1_546/Y gnd vdd DFFPOSX1
XXNOR2X1_22 gnd XOR2X1_12/Y gnd NAND2X1_58/B vdd XNOR2X1
XXNOR2X1_100 XOR2X1_94/A XOR2X1_98/Y gnd OR2X2_87/A vdd XNOR2X1
XXOR2X1_292 XOR2X1_292/A INVX1_460/A gnd INVX1_582/A vdd XOR2X1
XNOR2X1_112 OR2X2_76/A OR2X2_76/B gnd NOR2X1_112/Y vdd NOR2X1
XNAND2X1_193 OAI21X1_161/Y NAND3X1_170/B gnd XNOR2X1_87/A vdd NAND2X1
XDFFPOSX1_259 INVX1_207/A CLKBUF1_17/Y INVX1_511/Y gnd vdd DFFPOSX1
XAOI21X1_91 NOR2X1_85/Y AOI21X1_91/B INVX1_84/A gnd NOR2X1_87/A vdd AOI21X1
XOAI21X1_620 NOR2X1_424/Y NOR2X1_425/Y INVX1_526/A gnd NOR2X1_429/B vdd OAI21X1
XOR2X2_80 OR2X2_80/A OR2X2_80/B gnd OR2X2_80/Y vdd OR2X2
XINVX1_441 BUFX2_231/A gnd INVX1_441/Y vdd INVX1
XBUFX2_94 gnd gnd BUFX2_94/Y vdd BUFX2
XXOR2X1_256 XOR2X1_256/A BUFX2_219/A gnd INVX1_404/A vdd XOR2X1
XFILL_13_8_1 gnd vdd FILL
XAOI21X1_393 XNOR2X1_217/Y AOI21X1_393/B INVX1_528/Y gnd AOI21X1_393/Y vdd AOI21X1
XFILL_15_6_0 gnd vdd FILL
XNAND2X1_157 NAND3X1_134/Y NAND2X1_157/B gnd XNOR2X1_70/A vdd NAND2X1
XAOI21X1_55 NOR2X1_55/Y AOI21X1_55/B INVX1_51/A gnd NOR2X1_57/A vdd AOI21X1
XDFFPOSX1_223 INVX1_147/A CLKBUF1_14/Y INVX1_533/A gnd vdd DFFPOSX1
XOR2X2_44 OR2X2_44/A OR2X2_44/B gnd OR2X2_44/Y vdd OR2X2
XOAI21X1_584 NOR3X1_90/Y INVX2_78/A BUFX4_32/Y gnd AOI21X1_342/C vdd OAI21X1
XINVX1_405 INVX1_405/A gnd INVX1_405/Y vdd INVX1
XXOR2X1_220 XOR2X1_220/A BUFX2_203/A gnd INVX1_328/A vdd XOR2X1
XOAI21X1_8 AND2X2_2/Y NOR3X1_25/B INVX1_11/Y gnd NAND3X1_6/B vdd OAI21X1
XFILL_23_3_1 gnd vdd FILL
XFILL_25_1_0 gnd vdd FILL
XBUFX2_58 gnd gnd BUFX2_58/Y vdd BUFX2
XNAND2X1_698 NAND2X1_698/A INVX1_586/Y gnd DFFPOSX1_92/D vdd NAND2X1
XFILL_3_4_1 gnd vdd FILL
XFILL_5_2_0 gnd vdd FILL
XNAND2X1_121 gnd OR2X2_43/B gnd AOI21X1_74/A vdd NAND2X1
XAOI21X1_357 bloque_bytes[71] INVX1_500/Y INVX1_543/A gnd OAI21X1_596/C vdd AOI21X1
XNAND3X1_530 NOR2X1_440/B AND2X2_192/Y NOR2X1_441/Y gnd NOR2X1_442/B vdd NAND3X1
XAOI21X1_19 NOR2X1_25/Y AOI21X1_19/B INVX1_18/A gnd NOR2X1_27/A vdd AOI21X1
XDFFPOSX1_187 INVX1_99/A CLKBUF1_49/Y bloque_bytes[17] gnd vdd DFFPOSX1
XINVX1_369 INVX1_369/A gnd INVX1_369/Y vdd INVX1
XOAI21X1_548 NOR3X1_86/C INVX2_73/Y NOR3X1_86/A gnd AND2X2_156/A vdd OAI21X1
XXOR2X1_184 XOR2X1_184/A BUFX2_183/A gnd INVX1_252/A vdd XOR2X1
XNAND2X1_662 INVX1_557/Y AOI21X1_370/Y gnd AOI21X1_379/A vdd NAND2X1
XBUFX2_22 BUFX2_22/A gnd hash[21] vdd BUFX2
XAOI21X1_321 NAND3X1_482/Y NAND3X1_483/Y AOI21X1_321/C gnd AOI21X1_321/Y vdd AOI21X1
XDFFPOSX1_151 INVX1_48/A CLKBUF1_29/Y bloque_bytes[61] gnd vdd DFFPOSX1
XOAI21X1_67 AND2X2_23/Y NOR2X1_52/Y INVX1_47/Y gnd NAND3X1_69/A vdd OAI21X1
XNAND2X1_82 INVX1_52/A NAND2X1_82/B gnd OAI21X1_63/A vdd NAND2X1
XDFFPOSX1_85 INVX1_483/A CLKBUF1_6/Y NOR3X1_93/Y gnd vdd DFFPOSX1
XNAND3X1_494 INVX2_75/A INVX2_76/A AND2X2_165/B gnd INVX1_490/A vdd NAND3X1
XXOR2X1_148 XOR2X1_148/A BUFX2_169/A gnd XOR2X1_148/Y vdd XOR2X1
XOAI21X1_512 NOR3X1_81/A INVX1_418/A OAI21X1_512/C gnd NOR2X1_326/A vdd OAI21X1
XINVX1_333 INVX1_333/A gnd INVX1_333/Y vdd INVX1
XNAND2X1_626 AND2X2_172/B INVX2_83/A gnd NAND2X1_626/Y vdd NAND2X1
XOAI21X1_31 AND2X2_10/Y NOR2X1_30/Y INVX1_24/A gnd AOI21X1_25/A vdd OAI21X1
XNAND2X1_46 XOR2X1_2/A OR2X2_12/B gnd NAND3X1_30/B vdd NAND2X1
XNAND3X1_458 INVX1_418/Y AOI21X1_303/A NOR3X1_82/Y gnd AOI21X1_304/B vdd NAND3X1
XAOI21X1_285 INVX1_383/A AOI21X1_285/B INVX1_382/Y gnd NOR3X1_77/C vdd AOI21X1
XDFFPOSX1_115 INVX1_590/A CLKBUF1_25/Y bloque_bytes[89] gnd vdd DFFPOSX1
XDFFPOSX1_49 OR2X2_149/B CLKBUF1_6/Y NOR2X1_372/Y gnd vdd DFFPOSX1
XFILL_22_6_0 gnd vdd FILL
XINVX1_297 INVX1_297/A gnd INVX1_297/Y vdd INVX1
XFILL_2_7_0 gnd vdd FILL
XXOR2X1_92 OR2X2_84/A gnd gnd XOR2X1_92/Y vdd XOR2X1
XXOR2X1_112 AND2X2_77/A gnd gnd XOR2X1_112/Y vdd XOR2X1
XFILL_20_8_1 gnd vdd FILL
XOAI21X1_476 gnd XOR2X1_246/Y INVX1_381/Y gnd NAND3X1_425/B vdd OAI21X1
XNAND2X1_590 INVX1_453/Y NOR2X1_346/Y gnd NAND3X1_475/B vdd NAND2X1
XFILL_0_9_1 gnd vdd FILL
XAOI21X1_249 NAND3X1_365/Y AOI21X1_249/B NAND2X1_436/Y gnd AOI21X1_249/Y vdd AOI21X1
XDFFPOSX1_13 BUFX2_12/A CLKBUF1_48/Y NOR3X1_12/Y gnd vdd DFFPOSX1
XNAND2X1_10 NOR2X1_8/Y AOI21X1_3/Y gnd NOR2X1_10/A vdd NAND2X1
XFILL_32_1_0 gnd vdd FILL
XNAND3X1_422 INVX1_373/Y INVX1_376/Y AND2X2_137/A gnd NAND2X1_513/B vdd NAND3X1
XINVX1_261 INVX1_261/A gnd INVX1_261/Y vdd INVX1
XOAI21X1_440 INVX1_346/A INVX1_347/A INVX1_348/A gnd INVX1_350/A vdd OAI21X1
XFILL_30_3_1 gnd vdd FILL
XAND2X2_192 INVX1_582/A AND2X2_192/B gnd AND2X2_192/Y vdd AND2X2
XNAND3X1_87 OAI21X1_84/Y NAND3X1_87/B AOI21X1_62/Y gnd AND2X2_30/A vdd NAND3X1
XXOR2X1_56 XOR2X1_56/A OR2X2_44/A gnd OR2X2_52/B vdd XOR2X1
XOR2X2_139 OR2X2_139/A bloque_bytes[2] gnd OR2X2_139/Y vdd OR2X2
XNAND2X1_554 INVX1_416/Y NOR2X1_323/Y gnd NAND2X1_554/Y vdd NAND2X1
XAOI21X1_213 INVX1_212/A NAND3X1_309/B INVX1_211/Y gnd NOR3X1_59/C vdd AOI21X1
XNAND3X1_386 INVX1_325/A OAI21X1_419/Y NAND2X1_462/Y gnd NAND3X1_386/Y vdd NAND3X1
XMUX2X1_9 BUFX2_9/A INVX1_4/A MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XXOR2X1_20 XOR2X1_20/A XOR2X1_20/B gnd XOR2X1_39/B vdd XOR2X1
XNAND3X1_51 NAND3X1_51/A NAND3X1_51/B NAND3X1_51/C gnd AND2X2_18/A vdd NAND3X1
XINVX1_225 INVX1_225/A gnd INVX1_225/Y vdd INVX1
XOAI21X1_404 NOR3X1_69/C OAI21X1_404/B INVX1_313/A gnd NOR2X1_257/A vdd OAI21X1
XNOR2X1_437 BUFX2_244/A AND2X2_189/A gnd NOR2X1_437/Y vdd NOR2X1
XAND2X2_156 AND2X2_156/A NOR3X1_85/A gnd INVX1_585/A vdd AND2X2
XOR2X2_103 OR2X2_103/A INVX1_149/Y gnd OR2X2_103/Y vdd OR2X2
XNAND2X1_518 INVX1_382/A NAND2X1_517/Y gnd INVX1_380/A vdd NAND2X1
XAOI21X1_177 INVX2_50/Y XNOR2X1_122/A XNOR2X1_123/A gnd AOI21X1_177/Y vdd AOI21X1
XNAND3X1_350 INVX1_272/A INVX1_270/Y INVX1_271/Y gnd AOI21X1_236/B vdd NAND3X1
XINVX1_189 INVX1_189/A gnd INVX1_189/Y vdd INVX1
XINVX1_71 OR2X2_46/Y gnd INVX1_71/Y vdd INVX1
XFILL_18_1 gnd vdd FILL
XOAI21X1_368 BUFX2_192/A XOR2X1_194/Y INVX1_273/Y gnd NAND3X1_352/B vdd OAI21X1
XNAND3X1_15 NAND3X1_17/A NAND3X1_15/B NAND3X1_15/C gnd AND2X2_6/A vdd NAND3X1
XNOR2X1_401 NOR2X1_401/A NOR2X1_401/B gnd NOR2X1_401/Y vdd NOR2X1
XAND2X2_120 AND2X2_120/A NOR3X1_67/A gnd BUFX2_208/A vdd AND2X2
XNAND2X1_482 INVX1_343/Y NOR2X1_279/Y gnd NAND2X1_482/Y vdd NAND2X1
XAOI21X1_141 INVX2_41/Y XNOR2X1_94/Y XNOR2X1_96/A gnd NAND3X1_201/A vdd AOI21X1
XAND2X2_93 gnd OR2X2_122/B gnd AND2X2_93/Y vdd AND2X2
XFILL_27_8_1 gnd vdd FILL
XFILL_29_6_0 gnd vdd FILL
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XFILL_7_9_1 gnd vdd FILL
XFILL_9_7_0 gnd vdd FILL
XNAND3X1_314 AOI22X1_9/B INVX1_219/A INVX1_217/Y gnd AOI21X1_217/B vdd NAND3X1
XINVX1_153 INVX1_153/A gnd INVX1_153/Y vdd INVX1
XOAI21X1_332 gnd NOR2X1_204/B INVX1_227/Y gnd AOI21X1_222/A vdd OAI21X1
XNOR2X1_365 BUFX4_14/Y INVX1_478/Y gnd NOR2X1_365/Y vdd NOR2X1
XNAND2X1_446 INVX1_311/A NOR2X1_258/Y gnd NAND3X1_378/C vdd NAND2X1
XNAND3X1_278 NAND3X1_279/B NAND3X1_276/A NAND3X1_279/A gnd NAND3X1_278/Y vdd NAND3X1
XAOI21X1_105 INVX2_32/Y XNOR2X1_67/Y XNOR2X1_69/A gnd NAND3X1_147/A vdd AOI21X1
XAND2X2_57 gnd OR2X2_74/B gnd AND2X2_57/Y vdd AND2X2
XOAI21X1_296 AOI21X1_208/Y INVX1_204/A INVX1_203/Y gnd AND2X2_101/A vdd OAI21X1
XINVX1_117 INVX1_117/A gnd INVX1_117/Y vdd INVX1
XNOR2X1_329 NOR2X1_329/A NOR3X1_81/Y gnd NOR2X1_329/Y vdd NOR2X1
XNAND2X1_410 AOI21X1_241/A NAND2X1_410/B gnd XOR2X1_206/B vdd NAND2X1
XAND2X2_21 gnd OR2X2_26/B gnd AND2X2_21/Y vdd AND2X2
XNAND3X1_242 NAND3X1_242/A NAND2X1_269/B NAND3X1_242/C gnd NAND2X1_271/A vdd NAND3X1
XBUFX2_243 BUFX2_243/A gnd BUFX2_243/Y vdd BUFX2
XOAI21X1_260 INVX2_55/Y AND2X2_90/B INVX1_170/A gnd OAI21X1_261/B vdd OAI21X1
XNOR2X1_96 INVX1_95/Y NOR2X1_96/B gnd NOR2X1_96/Y vdd NOR2X1
XINVX2_81 INVX2_81/A gnd INVX2_81/Y vdd INVX2
XFILL_11_1_1 gnd vdd FILL
XNAND2X1_374 XOR2X1_188/B NOR2X1_208/Y gnd AOI21X1_224/C vdd NAND2X1
XNOR2X1_293 NOR2X1_293/A NOR3X1_75/Y gnd NOR2X1_293/Y vdd NOR2X1
XNOR2X1_60 gnd OR2X2_35/B gnd NOR2X1_60/Y vdd NOR2X1
XNAND3X1_206 NAND3X1_206/A NAND2X1_231/B NAND3X1_206/C gnd NAND2X1_233/A vdd NAND3X1
XFILL_36_6_0 gnd vdd FILL
XBUFX2_207 BUFX2_207/A gnd BUFX2_207/Y vdd BUFX2
XXNOR2X1_245 NOR2X1_440/B INVX2_91/Y gnd XNOR2X1_245/Y vdd XNOR2X1
XOAI21X1_224 AND2X2_79/Y NOR2X1_144/Y INVX1_147/Y gnd NAND3X1_235/A vdd OAI21X1
XINVX2_45 INVX2_45/A gnd INVX2_45/Y vdd INVX2
XFILL_34_8_1 gnd vdd FILL
XNOR2X1_257 NOR2X1_257/A NOR3X1_69/Y gnd NOR2X1_257/Y vdd NOR2X1
XNAND2X1_338 XNOR2X1_151/B NAND2X1_338/B gnd NOR2X1_188/B vdd NAND2X1
XBUFX2_171 BUFX2_171/A gnd BUFX2_171/Y vdd BUFX2
XCLKBUF1_48 BUFX4_2/Y gnd CLKBUF1_48/Y vdd CLKBUF1
XINVX1_586 INVX1_586/A gnd INVX1_586/Y vdd INVX1
XNAND3X1_170 NAND3X1_170/A NAND3X1_170/B AOI21X1_120/C gnd NAND2X1_195/A vdd NAND3X1
XNOR2X1_24 vdd OR2X2_5/B gnd NOR2X1_24/Y vdd NOR2X1
XXNOR2X1_209 bloque_bytes[49] bloque_bytes[9] gnd XNOR2X1_209/Y vdd XNOR2X1
XNAND2X1_302 NAND2X1_302/A INVX1_174/A gnd INVX1_172/A vdd NAND2X1
XOAI21X1_188 XNOR2X1_98/A AOI21X1_137/C AND2X2_66/B gnd XNOR2X1_99/A vdd OAI21X1
XNOR2X1_221 NOR2X1_221/A NOR3X1_63/Y gnd NOR2X1_221/Y vdd NOR2X1
XFILL_10_4_0 gnd vdd FILL
XDFFPOSX1_368 INVX1_467/A CLKBUF1_19/Y NAND3X1_526/Y gnd vdd DFFPOSX1
XFILL_5_2 gnd vdd FILL
XCLKBUF1_12 BUFX4_1/Y gnd CLKBUF1_12/Y vdd CLKBUF1
XNAND3X1_134 OAI21X1_129/Y NAND3X1_134/B AOI21X1_96/C gnd NAND3X1_134/Y vdd NAND3X1
XBUFX2_135 gnd gnd BUFX2_135/Y vdd BUFX2
XINVX1_550 INVX1_550/A gnd INVX1_550/Y vdd INVX1
XOAI21X1_152 AND2X2_53/Y NOR2X1_102/Y INVX1_102/Y gnd NAND3X1_161/A vdd OAI21X1
XXNOR2X1_95 XNOR2X1_94/Y INVX2_41/Y gnd AND2X2_77/A vdd XNOR2X1
XXNOR2X1_173 NOR2X1_257/Y NOR2X1_256/Y gnd XOR2X1_229/A vdd XNOR2X1
XNOR2X1_185 NOR2X1_185/A NOR3X1_57/Y gnd NOR2X1_185/Y vdd NOR2X1
XNAND2X1_266 NAND2X1_266/A NAND2X1_266/B gnd XOR2X1_139/A vdd NAND2X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_514 INVX1_514/A gnd INVX1_514/Y vdd INVX1
XFILL_18_1_1 gnd vdd FILL
XDFFPOSX1_332 INVX1_379/A CLKBUF1_19/Y NAND2X1_680/Y gnd vdd DFFPOSX1
XNOR3X1_65 NOR3X1_65/A NOR3X1_65/B NOR3X1_65/C gnd NOR3X1_65/Y vdd NOR3X1
XXNOR2X1_137 XOR2X1_151/Y XOR2X1_139/Y gnd XNOR2X1_138/A vdd XNOR2X1
XOAI21X1_116 AND2X2_40/Y NOR2X1_80/Y INVX1_79/A gnd AOI21X1_85/A vdd OAI21X1
XXNOR2X1_59 AOI21X1_93/B INVX2_29/Y gnd OR2X2_68/A vdd XNOR2X1
XNOR2X1_149 gnd AND2X2_81/B gnd NOR3X1_52/B vdd NOR2X1
XNOR3X1_29 INVX1_33/Y NOR3X1_29/B AND2X2_14/Y gnd NOR3X1_29/Y vdd NOR3X1
XNAND2X1_230 gnd OR2X2_89/B gnd NAND3X1_203/B vdd NAND2X1
XINVX1_478 INVX1_478/A gnd INVX1_478/Y vdd INVX1
XDFFPOSX1_296 INVX1_296/A CLKBUF1_21/Y NAND3X1_508/Y gnd vdd DFFPOSX1
XXNOR2X1_23 NAND2X1_58/B INVX2_17/Y gnd OR2X2_36/A vdd XNOR2X1
XXNOR2X1_101 XOR2X1_111/Y XOR2X1_99/Y gnd XNOR2X1_101/Y vdd XNOR2X1
XXOR2X1_293 XOR2X1_287/Y BUFX2_236/A gnd AND2X2_192/B vdd XOR2X1
XNAND2X1_194 gnd OR2X2_74/B gnd NAND3X1_169/B vdd NAND2X1
XNOR2X1_113 NOR2X1_113/A NOR3X1_44/Y gnd NOR2X1_113/Y vdd NOR2X1
XAOI21X1_92 INVX2_30/Y INVX1_85/Y NOR2X1_81/A gnd AOI21X1_92/Y vdd AOI21X1
XDFFPOSX1_260 INVX1_208/A CLKBUF1_17/Y INVX1_514/Y gnd vdd DFFPOSX1
XOR2X2_81 gnd OR2X2_81/B gnd OR2X2_81/Y vdd OR2X2
XOAI21X1_621 INVX1_547/Y bloque_bytes[38] INVX1_548/Y gnd OAI21X1_621/Y vdd OAI21X1
XXOR2X1_257 XOR2X1_251/Y BUFX2_220/A gnd XOR2X1_257/Y vdd XOR2X1
XINVX1_442 INVX1_442/A gnd INVX1_442/Y vdd INVX1
XFILL_15_6_1 gnd vdd FILL
XFILL_17_4_0 gnd vdd FILL
XBUFX2_95 gnd gnd BUFX2_95/Y vdd BUFX2
XAOI21X1_394 AOI21X1_394/A OR2X2_156/Y INVX1_591/A gnd NOR2X1_450/A vdd AOI21X1
XNAND2X1_158 INVX1_96/A NAND2X1_158/B gnd OAI21X1_131/A vdd NAND2X1
XAOI21X1_56 INVX2_21/Y INVX1_52/Y NOR2X1_51/A gnd AOI21X1_58/A vdd AOI21X1
XOR2X2_45 OR2X2_45/A OR2X2_45/B gnd OR2X2_45/Y vdd OR2X2
XOAI21X1_585 NOR3X1_95/C INVX2_78/Y INVX2_79/Y gnd AND2X2_175/A vdd OAI21X1
XDFFPOSX1_224 INVX1_149/A CLKBUF1_9/Y INVX1_548/A gnd vdd DFFPOSX1
XINVX1_406 INVX1_406/A gnd INVX1_406/Y vdd INVX1
XNAND2X1_699 INVX1_587/Y INVX1_586/A gnd NAND2X1_699/Y vdd NAND2X1
XXOR2X1_221 XOR2X1_215/Y BUFX2_204/A gnd XOR2X1_221/Y vdd XOR2X1
XBUFX2_59 gnd gnd BUFX2_59/Y vdd BUFX2
XOAI21X1_9 OAI21X1_9/A OAI21X1_9/B NOR3X1_25/Y gnd OAI21X1_9/Y vdd OAI21X1
XFILL_7_0_0 gnd vdd FILL
XNAND2X1_122 OR2X2_44/A OR2X2_44/B gnd AOI21X1_76/A vdd NAND2X1
XAOI21X1_358 bloque_bytes[74] INVX2_85/Y INVX1_531/A gnd OAI21X1_597/C vdd AOI21X1
XFILL_25_1_1 gnd vdd FILL
XFILL_5_2_1 gnd vdd FILL
XNAND3X1_531 INVX1_587/Y INVX1_588/Y INVX1_586/A gnd NOR2X1_444/B vdd NAND3X1
XAOI21X1_20 INVX2_12/Y INVX1_19/Y NOR2X1_21/A gnd AOI21X1_22/A vdd AOI21X1
XDFFPOSX1_188 INVX1_100/A CLKBUF1_49/Y bloque_bytes[18] gnd vdd DFFPOSX1
XOAI21X1_549 gnd NOR2X1_348/B INVX1_455/A gnd INVX1_458/A vdd OAI21X1
XINVX1_370 INVX1_370/A gnd INVX1_370/Y vdd INVX1
XXOR2X1_185 XOR2X1_185/A BUFX2_184/A gnd NOR2X1_222/B vdd XOR2X1
XNAND2X1_663 bloque_bytes[1] OR2X2_151/B gnd AOI21X1_380/B vdd NAND2X1
XBUFX2_23 BUFX2_23/A gnd hash[22] vdd BUFX2
XNAND2X1_83 gnd OR2X2_27/B gnd NAND3X1_64/B vdd NAND2X1
XNAND3X1_495 INVX1_481/A INVX1_482/Y AND2X2_173/Y gnd AOI21X1_341/B vdd NAND3X1
XAOI21X1_322 INVX1_470/Y AOI21X1_322/B INVX1_469/A gnd OAI21X1_564/A vdd AOI21X1
XDFFPOSX1_152 INVX1_50/A CLKBUF1_29/Y bloque_bytes[62] gnd vdd DFFPOSX1
XOAI21X1_68 OAI21X1_63/A OAI21X1_68/B OAI21X1_68/C gnd NAND3X1_74/C vdd OAI21X1
XDFFPOSX1_86 INVX1_484/A CLKBUF1_6/Y DFFPOSX1_86/D gnd vdd DFFPOSX1
XFILL_14_9_0 gnd vdd FILL
XXOR2X1_149 XOR2X1_149/A BUFX2_170/A gnd XOR2X1_149/Y vdd XOR2X1
XOAI21X1_513 NOR3X1_82/A NOR3X1_82/C INVX2_71/A gnd NOR2X1_325/A vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd hash[0] vdd BUFX2
XINVX1_334 INVX1_334/A gnd INVX1_334/Y vdd INVX1
XNAND2X1_627 INVX8_1/A NAND2X1_626/Y gnd NAND2X1_627/Y vdd NAND2X1
XNAND2X1_47 INVX2_15/Y OAI21X1_34/Y gnd OAI21X1_35/A vdd NAND2X1
XOAI21X1_32 AND2X2_11/Y NOR2X1_32/Y INVX1_25/A gnd OAI21X1_32/Y vdd OAI21X1
XDFFPOSX1_50 OR2X2_142/B CLKBUF1_14/Y NOR2X1_373/Y gnd vdd DFFPOSX1
XFILL_24_4_0 gnd vdd FILL
XAOI21X1_286 OAI21X1_484/Y NAND2X1_525/Y INVX2_69/A gnd AOI21X1_287/B vdd AOI21X1
XNAND3X1_459 INVX1_421/A AOI21X1_300/A AOI21X1_300/B gnd NAND2X1_569/A vdd NAND3X1
XFILL_4_5_0 gnd vdd FILL
XDFFPOSX1_116 INVX1_591/A CLKBUF1_25/Y bloque_bytes[90] gnd vdd DFFPOSX1
XFILL_22_6_1 gnd vdd FILL
XINVX1_298 INVX1_298/A gnd INVX1_298/Y vdd INVX1
XOAI21X1_477 gnd XOR2X1_246/Y INVX1_381/A gnd INVX1_383/A vdd OAI21X1
XFILL_2_7_1 gnd vdd FILL
XXOR2X1_93 OR2X2_85/A gnd gnd OR2X2_81/B vdd XOR2X1
XXOR2X1_113 OR2X2_101/A gnd gnd OR2X2_97/B vdd XOR2X1
XNAND2X1_591 OAI21X1_546/Y NAND3X1_475/B gnd BUFX2_26/A vdd NAND2X1
XAOI21X1_250 INVX1_299/Y AOI21X1_250/B INVX1_298/A gnd OAI21X1_393/A vdd AOI21X1
XDFFPOSX1_14 BUFX2_13/A CLKBUF1_43/Y NOR3X1_13/Y gnd vdd DFFPOSX1
XNAND2X1_11 INVX1_5/A INVX2_8/Y gnd NAND3X1_2/A vdd NAND2X1
XFILL_32_1_1 gnd vdd FILL
XNAND3X1_423 INVX2_69/A NAND3X1_423/B NAND3X1_423/C gnd NOR3X1_77/A vdd NAND3X1
XAND2X2_193 gnd gnd gnd NOR3X1_97/C vdd AND2X2
XXOR2X1_57 XOR2X1_57/A OR2X2_45/A gnd OR2X2_53/B vdd XOR2X1
XINVX1_262 INVX1_262/A gnd INVX1_262/Y vdd INVX1
XOAI21X1_441 INVX1_346/A INVX1_347/A INVX1_348/Y gnd OAI21X1_441/Y vdd OAI21X1
XNAND3X1_88 INVX1_59/Y NAND3X1_88/B OR2X2_37/Y gnd NAND3X1_89/C vdd NAND3X1
XOR2X2_140 OR2X2_140/A bloque_bytes[6] gnd OR2X2_140/Y vdd OR2X2
XNAND2X1_555 INVX1_417/Y NOR2X1_324/Y gnd NAND2X1_555/Y vdd NAND2X1
XAOI21X1_214 AOI21X1_214/A AOI21X1_214/B INVX2_60/A gnd AOI21X1_215/B vdd AOI21X1
XNAND3X1_387 INVX1_326/A AOI21X1_261/B INVX1_325/Y gnd INVX1_332/A vdd NAND3X1
XINVX1_226 INVX1_226/A gnd INVX1_226/Y vdd INVX1
XXOR2X1_21 XOR2X1_5/A XOR2X1_21/B gnd XOR2X1_21/Y vdd XOR2X1
XNAND3X1_52 INVX1_37/Y NAND3X1_52/B OR2X2_21/Y gnd NAND3X1_53/C vdd NAND3X1
XNAND2X1_519 INVX1_381/A NOR2X1_303/Y gnd NAND3X1_425/C vdd NAND2X1
XOAI21X1_405 NOR2X1_257/Y NOR2X1_256/B AOI22X1_14/C gnd XOR2X1_224/A vdd OAI21X1
XAND2X2_157 AND2X2_157/A AND2X2_157/B gnd INVX1_589/A vdd AND2X2
XNOR2X1_438 NOR2X1_437/Y XOR2X1_306/A gnd NOR2X1_438/Y vdd NOR2X1
XOR2X2_104 OR2X2_104/A OR2X2_104/B gnd OR2X2_104/Y vdd OR2X2
XFILL_21_9_0 gnd vdd FILL
XAOI21X1_178 AOI21X1_178/A AOI21X1_178/B NAND2X1_284/Y gnd OAI21X1_244/A vdd AOI21X1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XNAND3X1_351 INVX1_274/A AOI21X1_235/B INVX1_269/Y gnd AOI22X1_12/C vdd NAND3X1
XINVX1_190 NOR3X1_57/B gnd INVX1_190/Y vdd INVX1
XFILL_18_2 gnd vdd FILL
XOAI21X1_369 BUFX2_192/A XOR2X1_194/Y INVX1_273/A gnd AOI22X1_12/B vdd OAI21X1
XAND2X2_121 AND2X2_121/A AND2X2_121/B gnd AND2X2_121/Y vdd AND2X2
XNAND3X1_16 INVX1_15/Y NAND3X1_16/B OR2X2_5/Y gnd NAND3X1_16/Y vdd NAND3X1
XNOR2X1_402 NOR2X1_402/A INVX1_490/A gnd AND2X2_172/B vdd NOR2X1
XNAND2X1_483 NAND3X1_399/Y INVX1_351/A gnd XNOR2X1_180/B vdd NAND2X1
XFILL_31_4_0 gnd vdd FILL
XFILL_9_7_1 gnd vdd FILL
XAOI21X1_142 AOI21X1_140/Y AOI21X1_142/B AOI21X1_142/C gnd AOI21X1_142/Y vdd AOI21X1
XNAND3X1_315 INVX1_209/Y NAND2X1_350/A NOR3X1_60/Y gnd AOI21X1_216/B vdd NAND3X1
XAND2X2_94 gnd OR2X2_123/B gnd AND2X2_94/Y vdd AND2X2
XFILL_29_6_1 gnd vdd FILL
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XOAI21X1_333 BUFX2_185/A NOR2X1_211/B INVX1_239/A gnd NAND2X1_376/A vdd OAI21X1
XNOR2X1_366 BUFX4_16/Y INVX2_75/Y gnd NOR2X1_366/Y vdd NOR2X1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XNAND2X1_447 INVX1_311/Y NOR2X1_258/Y gnd INVX1_314/A vdd NAND2X1
XNAND3X1_279 NAND3X1_279/A NAND3X1_279/B NOR3X1_55/Y gnd INVX1_184/A vdd NAND3X1
XAOI21X1_106 AOI21X1_106/A AOI21X1_106/B OAI21X1_140/B gnd OAI21X1_142/A vdd AOI21X1
XAND2X2_58 gnd OR2X2_75/B gnd AND2X2_58/Y vdd AND2X2
XOAI21X1_297 NOR2X1_185/A NOR3X1_57/Y OAI21X1_297/C gnd OAI21X1_297/Y vdd OAI21X1
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XNAND2X1_411 INVX1_265/A NOR2X1_228/Y gnd AOI21X1_238/B vdd NAND2X1
XNOR2X1_330 BUFX2_228/A NOR2X1_330/B gnd NOR2X1_330/Y vdd NOR2X1
XAND2X2_22 gnd OR2X2_27/B gnd AND2X2_22/Y vdd AND2X2
XNAND3X1_243 NAND3X1_242/C NAND3X1_242/A NOR3X1_51/Y gnd INVX1_162/A vdd NAND3X1
XBUFX2_244 BUFX2_244/A gnd BUFX2_244/Y vdd BUFX2
XFILL_28_9_0 gnd vdd FILL
XOAI21X1_261 OAI21X1_261/A OAI21X1_261/B INVX1_172/Y gnd NAND3X1_274/C vdd OAI21X1
XNOR2X1_97 NOR2X1_97/A NOR2X1_96/Y gnd NOR2X1_97/Y vdd NOR2X1
XNAND2X1_375 INVX1_239/Y NOR2X1_211/Y gnd NAND2X1_375/Y vdd NAND2X1
XINVX2_82 INVX2_82/A gnd INVX2_82/Y vdd INVX2
XNOR2X1_294 BUFX2_216/A NOR2X1_294/B gnd NOR2X1_294/Y vdd NOR2X1
XNAND3X1_207 NAND3X1_206/C NAND3X1_206/A NOR3X1_47/Y gnd INVX1_140/A vdd NAND3X1
XNOR2X1_61 NOR2X1_61/A INVX2_24/A gnd XOR2X1_50/B vdd NOR2X1
XFILL_36_6_1 gnd vdd FILL
XBUFX2_208 BUFX2_208/A gnd BUFX2_208/Y vdd BUFX2
XXNOR2X1_246 OAI21X1_631/A INVX1_581/A gnd XNOR2X1_246/Y vdd XNOR2X1
XOAI21X1_225 XNOR2X1_116/A AOI21X1_166/C NOR2X1_145/Y gnd NOR2X1_146/B vdd OAI21X1
XINVX2_46 INVX2_46/A gnd INVX2_46/Y vdd INVX2
XNOR2X1_258 BUFX2_204/A XOR2X1_212/Y gnd NOR2X1_258/Y vdd NOR2X1
XNAND2X1_339 INVX1_200/Y NOR2X1_188/B gnd NAND2X1_340/A vdd NAND2X1
XCLKBUF1_49 BUFX4_7/Y gnd CLKBUF1_49/Y vdd CLKBUF1
XBUFX2_172 OR2X2_125/A gnd BUFX2_172/Y vdd BUFX2
XINVX1_587 INVX1_587/A gnd INVX1_587/Y vdd INVX1
XNAND3X1_171 AOI21X1_120/C NAND3X1_170/A NOR3X1_43/Y gnd INVX1_118/A vdd NAND3X1
XNOR2X1_25 NOR2X1_25/A INVX1_16/Y gnd NOR2X1_25/Y vdd NOR2X1
XOAI21X1_189 AND2X2_67/Y NOR2X1_124/Y INVX1_125/A gnd OAI21X1_189/Y vdd OAI21X1
XXNOR2X1_210 bloque_bytes[50] bloque_bytes[10] gnd XNOR2X1_210/Y vdd XNOR2X1
XNAND2X1_303 INVX2_55/A AND2X2_90/Y gnd AOI21X1_190/C vdd NAND2X1
XFILL_12_2_0 gnd vdd FILL
XNOR2X1_222 BUFX2_188/A NOR2X1_222/B gnd NOR2X1_222/Y vdd NOR2X1
XINVX2_10 INVX2_10/A gnd INVX2_10/Y vdd INVX2
XFILL_10_4_1 gnd vdd FILL
XDFFPOSX1_369 XNOR2X1_206/B CLKBUF1_22/Y NAND3X1_527/Y gnd vdd DFFPOSX1
XFILL_5_3 gnd vdd FILL
XNAND3X1_135 AOI21X1_96/C OAI21X1_129/Y NOR3X1_39/Y gnd INVX1_96/A vdd NAND3X1
XXNOR2X1_174 NOR2X1_261/Y XNOR2X1_174/B gnd XNOR2X1_174/Y vdd XNOR2X1
XINVX1_551 INVX1_551/A gnd INVX1_551/Y vdd INVX1
XBUFX2_136 gnd gnd BUFX2_136/Y vdd BUFX2
XCLKBUF1_13 BUFX4_2/Y gnd CLKBUF1_13/Y vdd CLKBUF1
XOAI21X1_153 OAI21X1_153/A XNOR2X1_79/B OAI21X1_153/C gnd NAND3X1_164/C vdd OAI21X1
XNOR2X1_186 BUFX2_176/A NOR2X1_186/B gnd NOR2X1_186/Y vdd NOR2X1
XXNOR2X1_96 XNOR2X1_96/A XNOR2X1_96/B gnd OR2X2_101/A vdd XNOR2X1
XNAND2X1_267 INVX2_50/Y XNOR2X1_122/A gnd XNOR2X1_123/B vdd NAND2X1
XNOR3X1_66 NOR3X1_66/A INVX2_63/Y NOR3X1_66/C gnd NOR3X1_66/Y vdd NOR3X1
XFILL_35_9_0 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XINVX1_515 bloque_bytes[59] gnd INVX1_515/Y vdd INVX1
XBUFX2_100 gnd gnd BUFX2_100/Y vdd BUFX2
XDFFPOSX1_333 INVX1_381/A CLKBUF1_45/Y OR2X2_147/Y gnd vdd DFFPOSX1
XXNOR2X1_60 AOI21X1_93/C XNOR2X1_60/B gnd OR2X2_69/A vdd XNOR2X1
XXNOR2X1_138 XNOR2X1_138/A OR2X2_119/Y gnd INVX1_175/A vdd XNOR2X1
XOAI21X1_117 AND2X2_41/Y NOR2X1_82/Y INVX1_80/A gnd OAI21X1_117/Y vdd OAI21X1
XNAND2X1_231 NAND2X1_231/A NAND2X1_231/B gnd AOI21X1_153/C vdd NAND2X1
XNOR2X1_150 gnd AND2X2_82/B gnd NOR2X1_150/Y vdd NOR2X1
XNOR3X1_30 INVX1_34/Y NOR3X1_30/B NOR3X1_30/C gnd NOR2X1_43/B vdd NOR3X1
XDFFPOSX1_297 XNOR2X1_170/B CLKBUF1_11/Y AOI21X1_385/C gnd vdd DFFPOSX1
XINVX1_479 INVX1_479/A gnd INVX1_479/Y vdd INVX1
XXNOR2X1_24 NAND2X1_60/Y NAND3X1_42/C gnd OR2X2_37/A vdd XNOR2X1
XXNOR2X1_102 XNOR2X1_101/Y OR2X2_87/Y gnd INVX1_131/A vdd XNOR2X1
XXOR2X1_294 XOR2X1_294/A BUFX2_237/A gnd INVX1_583/A vdd XOR2X1
XNOR2X1_114 OR2X2_77/A OR2X2_77/B gnd NOR2X1_114/Y vdd NOR2X1
XNAND2X1_195 NAND2X1_195/A NAND2X1_195/B gnd XNOR2X1_88/A vdd NAND2X1
XAOI21X1_93 INVX2_29/Y AOI21X1_93/B AOI21X1_93/C gnd AOI21X1_93/Y vdd AOI21X1
XOR2X2_82 gnd OR2X2_82/B gnd OR2X2_82/Y vdd OR2X2
XDFFPOSX1_261 INVX1_210/A CLKBUF1_17/Y INVX1_517/Y gnd vdd DFFPOSX1
XOAI21X1_622 AND2X2_187/Y NOR2X1_430/Y INVX1_545/A gnd OR2X2_149/A vdd OAI21X1
XFILL_19_2_0 gnd vdd FILL
XXOR2X1_258 XOR2X1_258/A BUFX2_221/A gnd NOR2X1_319/B vdd XOR2X1
XINVX1_443 INVX1_443/A gnd INVX1_443/Y vdd INVX1
XFILL_17_4_1 gnd vdd FILL
XBUFX2_96 gnd gnd BUFX2_96/Y vdd BUFX2
XAOI21X1_395 AOI21X1_395/A AOI21X1_395/B NAND3X1_535/C gnd NOR2X1_448/A vdd AOI21X1
XNAND2X1_159 gnd OR2X2_59/B gnd AOI21X1_98/A vdd NAND2X1
XAOI21X1_57 INVX2_20/Y AOI21X1_57/B AOI21X1_57/C gnd NAND3X1_75/A vdd AOI21X1
XOR2X2_46 OR2X2_46/A OR2X2_46/B gnd OR2X2_46/Y vdd OR2X2
XDFFPOSX1_225 XOR2X1_131/B CLKBUF1_6/Y OR2X2_149/B gnd vdd DFFPOSX1
XOAI21X1_586 NOR3X1_95/C INVX1_492/A BUFX4_32/Y gnd NOR2X1_405/B vdd OAI21X1
XINVX1_407 INVX1_407/A gnd INVX1_407/Y vdd INVX1
XBUFX2_60 gnd gnd BUFX2_60/Y vdd BUFX2
XNAND2X1_700 OAI21X1_632/Y NAND2X1_699/Y gnd NAND2X1_700/Y vdd NAND2X1
XXOR2X1_222 AND2X2_121/Y BUFX2_205/A gnd NOR2X1_271/B vdd XOR2X1
XFILL_7_0_1 gnd vdd FILL
XNAND2X1_123 INVX2_27/Y NAND3X1_110/C gnd XNOR2X1_53/A vdd NAND2X1
XAOI21X1_359 bloque_bytes[77] INVX2_86/Y INVX1_533/A gnd AOI21X1_359/Y vdd AOI21X1
XAOI21X1_21 INVX2_11/Y XNOR2X1_5/A XNOR2X1_6/A gnd NAND3X1_21/A vdd AOI21X1
XNAND3X1_532 INVX1_590/A NAND2X1_705/Y OR2X2_155/Y gnd NAND3X1_533/A vdd NAND3X1
XDFFPOSX1_189 INVX1_101/A CLKBUF1_16/Y bloque_bytes[19] gnd vdd DFFPOSX1
XDFFPOSX1_1 BUFX4_8/A CLKBUF1_28/Y NOR2X1_17/Y gnd vdd DFFPOSX1
XOR2X2_10 gnd AND2X2_9/B gnd OR2X2_10/Y vdd OR2X2
XXOR2X1_186 XOR2X1_186/A BUFX2_185/A gnd NOR2X1_223/B vdd XOR2X1
XINVX1_371 INVX1_371/A gnd INVX1_371/Y vdd INVX1
XOAI21X1_550 NOR3X1_85/A INVX1_456/A OAI21X1_556/B gnd NOR2X1_350/A vdd OAI21X1
XNAND2X1_664 INVX1_559/Y AOI21X1_371/Y gnd NAND2X1_664/Y vdd NAND2X1
XBUFX2_24 BUFX2_24/A gnd hash[23] vdd BUFX2
XFILL_31_1 gnd vdd FILL
XNAND2X1_84 OR2X2_28/A OR2X2_28/B gnd AOI21X1_52/A vdd NAND2X1
XOAI21X1_69 OAI21X1_69/A OAI21X1_69/B AND2X2_24/B gnd XNOR2X1_36/A vdd OAI21X1
XAOI21X1_323 AND2X2_159/B NOR2X1_384/A OAI21X1_567/Y gnd DFFPOSX1_60/D vdd AOI21X1
XNAND3X1_496 NOR2X1_387/Y NOR2X1_388/Y NOR3X1_89/Y gnd NOR3X1_90/C vdd NAND3X1
XFILL_16_7_0 gnd vdd FILL
XDFFPOSX1_153 XOR2X1_41/B CLKBUF1_29/Y bloque_bytes[63] gnd vdd DFFPOSX1
XDFFPOSX1_87 INVX2_80/A CLKBUF1_15/Y DFFPOSX1_87/D gnd vdd DFFPOSX1
XFILL_14_9_1 gnd vdd FILL
XINVX1_335 INVX1_335/A gnd INVX1_335/Y vdd INVX1
XOAI21X1_514 gnd NOR2X1_327/B INVX1_419/Y gnd NAND3X1_451/B vdd OAI21X1
XXOR2X1_150 XOR2X1_150/A XOR2X1_150/B gnd BUFX2_178/A vdd XOR2X1
XNAND2X1_628 INVX1_480/A AND2X2_172/Y gnd NAND2X1_628/Y vdd NAND2X1
XBUFX2_2 BUFX2_2/A gnd hash[1] vdd BUFX2
XAOI21X1_287 AOI21X1_287/A AOI21X1_287/B INVX1_389/Y gnd AOI21X1_288/A vdd AOI21X1
XNAND2X1_48 AND2X2_12/B AND2X2_12/A gnd OAI21X1_35/B vdd NAND2X1
XOAI21X1_33 AND2X2_11/Y NOR2X1_32/Y INVX1_25/Y gnd NAND3X1_35/A vdd OAI21X1
XDFFPOSX1_51 OR2X2_143/B CLKBUF1_30/Y NOR2X1_374/Y gnd vdd DFFPOSX1
XFILL_24_4_1 gnd vdd FILL
XFILL_26_2_0 gnd vdd FILL
XNAND3X1_460 INVX1_432/Y INVX1_431/A OAI21X1_525/Y gnd AND2X2_149/B vdd NAND3X1
XDFFPOSX1_117 INVX1_592/A CLKBUF1_25/Y bloque_bytes[91] gnd vdd DFFPOSX1
XFILL_4_5_1 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XINVX1_299 INVX1_299/A gnd INVX1_299/Y vdd INVX1
XOAI21X1_478 BUFX2_219/A INVX1_385/A INVX1_386/A gnd INVX1_388/A vdd OAI21X1
XXOR2X1_94 XOR2X1_94/A gnd gnd OR2X2_82/B vdd XOR2X1
XXOR2X1_114 BUFX2_161/A gnd gnd OR2X2_98/B vdd XOR2X1
XNAND2X1_592 INVX1_454/Y NOR2X1_347/Y gnd NAND3X1_475/C vdd NAND2X1
XNAND2X1_12 INVX1_6/A INVX2_9/Y gnd NAND3X1_2/B vdd NAND2X1
XNAND3X1_424 INVX1_382/A NAND2X1_517/Y INVX2_69/Y gnd OAI21X1_474/C vdd NAND3X1
XAOI21X1_251 INVX1_312/A NAND3X1_375/Y INVX1_307/Y gnd NOR2X1_256/B vdd AOI21X1
XDFFPOSX1_15 BUFX2_14/A CLKBUF1_48/Y NOR3X1_14/Y gnd vdd DFFPOSX1
XNAND3X1_89 OAI21X1_84/Y OAI21X1_87/Y NAND3X1_89/C gnd NAND3X1_89/Y vdd NAND3X1
XAND2X2_194 gnd gnd gnd NOR3X1_98/C vdd AND2X2
XXOR2X1_58 XOR2X1_58/A BUFX2_253/A gnd XOR2X1_58/Y vdd XOR2X1
XINVX1_263 INVX1_263/A gnd INVX1_263/Y vdd INVX1
XOAI21X1_442 NOR3X1_73/C OAI21X1_442/B INVX1_351/A gnd NOR2X1_281/A vdd OAI21X1
XOR2X2_141 OR2X2_141/A bloque_bytes[7] gnd OR2X2_141/Y vdd OR2X2
XNAND2X1_556 INVX1_420/A NAND2X1_555/Y gnd INVX1_418/A vdd NAND2X1
XAOI21X1_215 NAND2X1_350/A AOI21X1_215/B INVX1_218/Y gnd AOI21X1_216/A vdd AOI21X1
XNAND3X1_388 INVX1_327/Y INVX1_328/Y INVX1_329/Y gnd NAND3X1_388/Y vdd NAND3X1
XINVX1_227 INVX1_227/A gnd INVX1_227/Y vdd INVX1
XOAI21X1_406 BUFX2_204/A XOR2X1_212/Y INVX1_311/Y gnd NAND3X1_378/B vdd OAI21X1
XXOR2X1_22 OR2X2_28/A gnd gnd XOR2X1_22/Y vdd XOR2X1
XNAND3X1_53 NAND3X1_51/A NAND3X1_53/B NAND3X1_53/C gnd AOI21X1_41/A vdd NAND3X1
XAND2X2_158 BUFX4_33/Y AND2X2_158/B gnd AND2X2_158/Y vdd AND2X2
XFILL_23_7_0 gnd vdd FILL
XOR2X2_105 gnd OR2X2_105/B gnd OR2X2_105/Y vdd OR2X2
XNAND2X1_520 INVX1_381/Y NOR2X1_303/Y gnd AOI21X1_285/B vdd NAND2X1
XNOR2X1_439 INVX1_584/A XOR2X1_289/Y gnd NOR2X1_439/Y vdd NOR2X1
XFILL_3_8_0 gnd vdd FILL
XAOI21X1_179 NAND3X1_259/B OR2X2_114/Y INVX1_166/A gnd NOR2X1_163/A vdd AOI21X1
XFILL_21_9_1 gnd vdd FILL
XNAND2X1_1 target[7] NOR2X1_1/B gnd INVX1_1/A vdd NAND2X1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XNAND3X1_352 INVX1_274/A NAND3X1_352/B NAND3X1_352/C gnd AOI21X1_241/A vdd NAND3X1
XINVX1_191 INVX1_191/A gnd INVX1_191/Y vdd INVX1
XNOR2X1_403 INVX1_480/Y INVX2_77/Y gnd NOR2X1_403/Y vdd NOR2X1
XFILL_18_3 gnd vdd FILL
XOAI21X1_370 gnd NOR2X1_228/B INVX1_265/Y gnd AOI21X1_238/A vdd OAI21X1
XFILL_33_2_0 gnd vdd FILL
XAND2X2_122 AND2X2_122/A INVX1_301/Y gnd NOR3X1_70/A vdd AND2X2
XNAND3X1_17 NAND3X1_17/A NAND3X1_17/B NAND3X1_16/Y gnd AOI21X1_17/A vdd NAND3X1
XFILL_31_4_1 gnd vdd FILL
XNAND2X1_484 INVX1_349/A NOR2X1_282/Y gnd NAND3X1_404/C vdd NAND2X1
XNAND3X1_316 INVX1_212/A AOI21X1_212/A AOI21X1_212/B gnd NAND2X1_360/A vdd NAND3X1
XAND2X2_95 BUFX2_171/A OR2X2_124/B gnd AND2X2_95/Y vdd AND2X2
XAOI21X1_143 NAND2X1_232/Y OR2X2_90/Y INVX1_133/A gnd NOR2X1_133/A vdd AOI21X1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XINVX1_155 INVX1_155/A gnd INVX1_155/Y vdd INVX1
XOAI21X1_334 OAI21X1_334/A INVX1_242/A INVX1_241/Y gnd AND2X2_109/A vdd OAI21X1
XNOR2X1_367 BUFX4_16/Y INVX2_76/Y gnd NOR2X1_367/Y vdd NOR2X1
XNAND2X1_448 AOI21X1_257/A AOI21X1_257/B gnd XOR2X1_224/B vdd NAND2X1
XAOI21X1_107 NAND2X1_175/Y OR2X2_66/Y INVX1_100/A gnd NOR2X1_103/A vdd AOI21X1
XNAND3X1_280 INVX1_178/A NAND3X1_281/B OR2X2_123/Y gnd AOI21X1_192/B vdd NAND3X1
XAND2X2_59 OR2X2_76/A OR2X2_76/B gnd AND2X2_59/Y vdd AND2X2
XOAI21X1_298 AOI21X1_210/Y INVX1_202/A INVX1_205/A gnd OAI21X1_298/Y vdd OAI21X1
XINVX1_119 OR2X2_80/Y gnd INVX1_119/Y vdd INVX1
XNAND2X1_412 XOR2X1_206/B NOR2X1_232/Y gnd NAND2X1_412/Y vdd NAND2X1
XNOR2X1_331 BUFX2_229/A NOR2X1_331/B gnd NOR2X1_331/Y vdd NOR2X1
XAND2X2_23 OR2X2_28/A OR2X2_28/B gnd AND2X2_23/Y vdd AND2X2
XNAND3X1_244 INVX1_156/A NAND3X1_245/B OR2X2_107/Y gnd AOI21X1_168/B vdd NAND3X1
XNOR2X1_98 gnd OR2X2_65/B gnd NOR3X1_41/B vdd NOR2X1
XFILL_30_7_0 gnd vdd FILL
XBUFX2_245 BUFX2_245/A gnd BUFX2_245/Y vdd BUFX2
XFILL_28_9_1 gnd vdd FILL
XINVX2_83 INVX2_83/A gnd INVX2_83/Y vdd INVX2
XOAI21X1_262 NOR2X1_167/A INVX1_174/Y INVX1_175/Y gnd OAI21X1_262/Y vdd OAI21X1
XNOR2X1_295 BUFX2_217/A XOR2X1_240/Y gnd NOR2X1_295/Y vdd NOR2X1
.ends

