module modulo_area ( gnd, vdd, inicio, bloque_bytes, clk, reset, target, terminado, hash);

input gnd, vdd;
input inicio;
input clk;
input reset;
output terminado;
input [95:0] bloque_bytes;
input [7:0] target;
output [23:0] hash;

CLKBUF1 CLKBUF1_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf7) );
CLKBUF1 CLKBUF1_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf6) );
CLKBUF1 CLKBUF1_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
CLKBUF1 CLKBUF1_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
CLKBUF1 CLKBUF1_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
CLKBUF1 CLKBUF1_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
CLKBUF1 CLKBUF1_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
CLKBUF1 CLKBUF1_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_2200_), .Y(_2200__bF_buf4) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_2200_), .Y(_2200__bF_buf3) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_2200_), .Y(_2200__bF_buf2) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_2200_), .Y(_2200__bF_buf1) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_2200_), .Y(_2200__bF_buf0) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf5) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf4) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf3) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf2) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf1) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(reset_bF_buf0) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_29_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .Y(_30_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .Y(_31_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_22_), .Y(_32_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(micro_ucr_hash1_hash_23_), .C(_32_), .D(target[6]), .Y(_33_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_23_), .Y(_34_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .Y(_35_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(target[7]), .C(micro_ucr_hash1_hash_22_), .D(_35_), .Y(_36_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_36_), .Y(_37_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_21_), .Y(_38_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_20_), .Y(_39_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(target[5]), .C(_39_), .D(target[4]), .Y(_40_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .Y(_41_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .Y(_42_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(micro_ucr_hash1_hash_21_), .C(micro_ucr_hash1_hash_20_), .D(_42_), .Y(_43_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_43_), .C(_37_), .Y(_44_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .Y(_45_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_18_), .Y(_46_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(micro_ucr_hash1_hash_19_), .C(_46_), .D(target[2]), .Y(_47_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_19_), .Y(_48_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .Y(_49_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(target[3]), .C(micro_ucr_hash1_hash_18_), .D(_49_), .Y(_50_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_50_), .Y(_51_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .Y(_52_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_17_), .Y(_53_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_16_), .Y(_54_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(target[1]), .C(_54_), .D(target[0]), .Y(_55_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_17_), .B(_52_), .C(_55_), .Y(_56_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(_48_), .Y(_57_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(_48_), .Y(_58_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(_46_), .Y(_59_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_59_), .C(_57_), .Y(_60_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_51_), .C(_60_), .Y(_61_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_21_), .B(_41_), .C(_40_), .Y(_62_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .B(_34_), .Y(_63_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .B(_34_), .Y(_64_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .B(_32_), .Y(_65_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_65_), .C(_63_), .Y(_66_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_37_), .C(_66_), .Y(_67_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_44_), .C(_67_), .Y(_68_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .B(micro_ucr_hash1_hash_15_), .Y(_69_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(target[6]), .B(micro_ucr_hash1_hash_14_), .Y(_70_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_70_), .Y(_71_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_13_), .Y(_72_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_12_), .Y(_73_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(target[5]), .C(target[4]), .D(_73_), .Y(_74_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(micro_ucr_hash1_hash_13_), .C(_42_), .D(micro_ucr_hash1_hash_12_), .Y(_75_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .Y(_76_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_71_), .Y(_77_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(micro_ucr_hash1_hash_11_), .C(_49_), .D(micro_ucr_hash1_hash_10_), .Y(_78_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_11_), .Y(_79_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_10_), .Y(_80_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(target[3]), .C(target[2]), .D(_80_), .Y(_81_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_81_), .Y(_82_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_9_), .Y(_83_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_8_), .Y(_84_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(target[1]), .C(target[0]), .D(_84_), .Y(_85_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(micro_ucr_hash1_hash_9_), .C(_85_), .Y(_86_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(_79_), .Y(_87_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(target[2]), .B(_80_), .Y(_88_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(target[3]), .B(_79_), .Y(_89_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_88_), .C(_87_), .Y(_90_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_82_), .C(_90_), .Y(_91_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .B(_72_), .Y(_92_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(target[4]), .B(_73_), .Y(_93_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(target[5]), .B(_72_), .Y(_94_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_93_), .C(_92_), .Y(_95_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_hash_15_), .Y(_96_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .B(_96_), .Y(_97_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(target[7]), .B(_96_), .Y(_98_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(micro_ucr_hash1_hash_14_), .Y(_99_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_98_), .C(_97_), .Y(_100_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_71_), .C(_100_), .Y(_1_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_77_), .C(_1_), .Y(_2_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(target[7]), .C(micro_ucr_hash1_hash_22_), .D(_35_), .Y(_3_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(micro_ucr_hash1_hash_23_), .C(_32_), .D(target[6]), .Y(_4_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_3_), .B(_4_), .Y(_5_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_43_), .Y(_6_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_6_), .Y(_7_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_70_), .Y(_8_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_75_), .Y(_9_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(_8_), .Y(_10_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(target[3]), .C(target[2]), .D(_80_), .Y(_11_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(micro_ucr_hash1_hash_11_), .C(_49_), .D(micro_ucr_hash1_hash_10_), .Y(_12_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_12_), .Y(_13_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(target[1]), .B(_83_), .Y(_14_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .Y(_15_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(micro_ucr_hash1_hash_9_), .C(_15_), .D(micro_ucr_hash1_hash_8_), .Y(_16_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(target[0]), .B(_84_), .Y(_17_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_17_), .C(_16_), .Y(_18_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_18_), .Y(_19_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(target[3]), .C(micro_ucr_hash1_hash_18_), .D(_49_), .Y(_20_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(micro_ucr_hash1_hash_19_), .C(_46_), .D(target[2]), .Y(_21_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_20_), .B(_21_), .Y(_22_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(micro_ucr_hash1_hash_17_), .C(micro_ucr_hash1_hash_16_), .D(_15_), .Y(_23_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(target[1]), .C(_54_), .D(target[0]), .Y(_24_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_24_), .Y(_25_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_25_), .Y(_26_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(_26_), .C(_19_), .D(_10_), .Y(_27_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_68_), .C(_2_), .Y(_28_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_28_), .C(_30_), .Y(_0_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(hash[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(terminado) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0_), .Q(_101_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__4_), .B(gnd), .Y(micro_ucr_hash1_a_1__0_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__5_), .B(gnd), .Y(micro_ucr_hash1_a_1__1_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__6_), .B(gnd), .Y(micro_ucr_hash1_a_1__2_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__7_), .B(gnd), .Y(micro_ucr_hash1_a_1__3_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_0__4_), .B(gnd), .Y(micro_ucr_hash1_a_1__4_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_0__5_), .B(vdd), .Y(micro_ucr_hash1_a_1__5_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_0__6_), .B(vdd), .Y(micro_ucr_hash1_a_1__6_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_0__7_), .B(vdd), .Y(micro_ucr_hash1_a_1__7_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[80]), .Y(_103_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__0_), .Y(_104_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_103_), .Y(micro_ucr_hash1_b_2__4_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_104_), .Y(_105_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__1_), .Y(_106_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__1_), .Y(_107_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[81]), .B(_107_), .C(_106_), .Y(_108_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[81]), .Y(_109_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__1_), .Y(_110_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__1_), .Y(_111_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_110_), .C(_109_), .Y(_112_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_108_), .Y(_113_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_105_), .Y(micro_ucr_hash1_b_2__5_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_112_), .C(_105_), .Y(_114_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_110_), .C(_111_), .Y(_115_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[82]), .Y(_116_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__2_), .Y(_117_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__2_), .Y(_118_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_117_), .C(_118_), .Y(_119_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__2_), .Y(_120_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__2_), .Y(_121_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_120_), .C(bloque_bytes[82]), .Y(_122_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_122_), .C(_115_), .Y(_123_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[82]), .B(_121_), .C(_120_), .Y(_124_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_117_), .C(_116_), .Y(_125_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_108_), .C(_124_), .Y(_126_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_123_), .Y(_127_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_114_), .Y(micro_ucr_hash1_b_2__6_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_125_), .C(_115_), .Y(_128_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_122_), .C(_108_), .Y(_129_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_129_), .Y(_130_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_114_), .C(_128_), .Y(_131_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[83]), .Y(_132_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__3_), .Y(_133_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__3_), .Y(_134_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_133_), .C(_132_), .Y(_135_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__3_), .Y(_136_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_0__3_), .Y(_137_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[83]), .B(_137_), .C(_136_), .Y(_138_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_138_), .C(_124_), .Y(_139_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_132_), .B(_137_), .C(_136_), .Y(_140_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_133_), .C(bloque_bytes[83]), .Y(_141_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_140_), .C(_119_), .Y(_142_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_142_), .Y(_102_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_102_), .Y(micro_ucr_hash1_b_2__7_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_2__4_), .B(gnd), .Y(micro_ucr_hash1_a_2__0_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_2__5_), .B(gnd), .Y(micro_ucr_hash1_a_2__1_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_2__6_), .B(gnd), .Y(micro_ucr_hash1_a_2__2_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_2__7_), .B(gnd), .Y(micro_ucr_hash1_a_2__3_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[72]), .Y(_212_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__0_), .Y(_213_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_213_), .B(_212_), .Y(micro_ucr_hash1_b_3__4_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_213_), .Y(_214_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__1_), .Y(_215_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__1_), .Y(_216_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[73]), .B(_216_), .C(_215_), .Y(_217_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[73]), .Y(_218_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__1_), .Y(_219_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__1_), .Y(_220_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_219_), .C(_218_), .Y(_221_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_217_), .Y(_222_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_214_), .Y(micro_ucr_hash1_b_3__5_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_221_), .C(_214_), .Y(_223_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_219_), .C(_220_), .Y(_224_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[74]), .Y(_225_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__2_), .Y(_226_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__2_), .Y(_227_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_226_), .C(_227_), .Y(_228_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__2_), .Y(_229_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__2_), .Y(_230_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_229_), .C(bloque_bytes[74]), .Y(_231_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_231_), .C(_224_), .Y(_232_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[74]), .B(_230_), .C(_229_), .Y(_233_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_226_), .C(_225_), .Y(_234_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_217_), .C(_233_), .Y(_235_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_232_), .Y(_236_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_223_), .Y(micro_ucr_hash1_b_3__6_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_234_), .C(_224_), .Y(_237_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_231_), .C(_217_), .Y(_238_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_238_), .Y(_239_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_223_), .C(_237_), .Y(_240_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[75]), .Y(_241_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__3_), .Y(_242_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__3_), .Y(_243_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_242_), .C(_241_), .Y(_244_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__3_), .Y(_245_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_1__3_), .Y(_246_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[75]), .B(_246_), .C(_245_), .Y(_247_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_247_), .C(_233_), .Y(_248_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_246_), .C(_245_), .Y(_249_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_242_), .C(bloque_bytes[75]), .Y(_250_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_249_), .C(_228_), .Y(_251_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_251_), .Y(_143_) );
XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_143_), .Y(micro_ucr_hash1_b_3__7_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[76]), .Y(_144_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__4_), .B(micro_ucr_hash1_a_1__4_), .Y(_145_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__4_), .B(micro_ucr_hash1_a_1__4_), .Y(_146_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_146_), .C(_145_), .Y(_147_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__4_), .B(micro_ucr_hash1_a_1__4_), .Y(_148_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__4_), .B(micro_ucr_hash1_a_1__4_), .Y(_149_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_148_), .C(bloque_bytes[76]), .Y(_150_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_147_), .C(_150_), .Y(_151_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_245_), .C(bloque_bytes[75]), .Y(_152_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_148_), .C(_144_), .Y(_153_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[76]), .B(_146_), .C(_145_), .Y(_154_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_154_), .C(_152_), .Y(_155_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_151_), .Y(_156_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(_251_), .Y(_157_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_231_), .B(_228_), .Y(_158_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_158_), .C(_248_), .Y(_159_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_223_), .C(_159_), .Y(_160_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_160_), .Y(_161_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_156_), .Y(micro_ucr_hash1_c_2__4_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_151_), .B(_155_), .Y(_162_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_162_), .C(_151_), .Y(_163_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[77]), .Y(_164_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__5_), .B(micro_ucr_hash1_a_1__5_), .Y(_165_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__5_), .B(micro_ucr_hash1_a_1__5_), .Y(_166_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_166_), .C(_165_), .Y(_167_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__5_), .B(micro_ucr_hash1_a_1__5_), .Y(_168_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__5_), .B(micro_ucr_hash1_a_1__5_), .Y(_169_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_168_), .C(bloque_bytes[77]), .Y(_170_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_170_), .C(_167_), .Y(_171_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_145_), .C(bloque_bytes[76]), .Y(_172_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[77]), .B(_166_), .C(_165_), .Y(_173_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_168_), .C(_164_), .Y(_174_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_173_), .C(_172_), .Y(_175_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_175_), .Y(_176_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(_176_), .Y(_177_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_177_), .Y(micro_ucr_hash1_c_2__5_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_175_), .C(_162_), .Y(_178_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_178_), .C(_160_), .Y(_179_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_173_), .Y(_180_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_172_), .Y(_181_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_181_), .Y(_182_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_172_), .B(_180_), .C(_151_), .Y(_183_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_182_), .Y(_184_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[78]), .Y(_185_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__6_), .B(micro_ucr_hash1_a_1__6_), .Y(_186_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_185_), .Y(_187_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_186_), .Y(_188_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_187_), .Y(_189_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_173_), .Y(_190_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_189_), .Y(_191_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_190_), .Y(_192_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_179_), .C(_192_), .Y(_193_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_156_), .Y(_194_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_194_), .C(_184_), .Y(_195_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_192_), .Y(_196_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_195_), .Y(_197_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_197_), .Y(micro_ucr_hash1_c_2__6_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_237_), .Y(_198_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_157_), .B(_198_), .C(_248_), .Y(_199_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_213_), .C(_222_), .Y(_200_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_236_), .C(_143_), .Y(_201_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_201_), .C(_194_), .Y(_202_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_151_), .C(_181_), .Y(_203_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_203_), .C(_196_), .Y(_204_) );
XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__7_), .B(bloque_bytes[79]), .Y(_205_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(micro_ucr_hash1_a_1__7_), .Y(_206_) );
XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_187_), .Y(_207_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_207_), .C(_204_), .Y(_208_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_190_), .Y(_209_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_207_), .Y(_210_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_209_), .C(_210_), .Y(_211_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_211_), .Y(micro_ucr_hash1_c_2__7_) );
XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__4_), .B(gnd), .Y(micro_ucr_hash1_a_3__0_) );
XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__5_), .B(gnd), .Y(micro_ucr_hash1_a_3__1_) );
XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__6_), .B(gnd), .Y(micro_ucr_hash1_a_3__2_) );
XOR2X1 XOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__7_), .B(gnd), .Y(micro_ucr_hash1_a_3__3_) );
XOR2X1 XOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_2__4_), .B(micro_ucr_hash1_b_2__4_), .Y(micro_ucr_hash1_a_3__4_) );
XOR2X1 XOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_2__5_), .B(micro_ucr_hash1_b_2__5_), .Y(micro_ucr_hash1_a_3__5_) );
XOR2X1 XOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_2__6_), .B(micro_ucr_hash1_b_2__6_), .Y(micro_ucr_hash1_a_3__6_) );
XOR2X1 XOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_2__7_), .B(micro_ucr_hash1_b_2__7_), .Y(micro_ucr_hash1_a_3__7_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[64]), .Y(_253_) );
XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__0_), .Y(_254_) );
XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_253_), .Y(micro_ucr_hash1_b_4__4_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_253_), .B(_254_), .Y(_255_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__1_), .Y(_256_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__1_), .Y(_257_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[65]), .B(_257_), .C(_256_), .Y(_258_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[65]), .Y(_259_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__1_), .Y(_260_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__1_), .Y(_261_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_260_), .C(_259_), .Y(_262_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_258_), .Y(_263_) );
XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_255_), .Y(micro_ucr_hash1_b_4__5_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_262_), .C(_255_), .Y(_264_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_260_), .C(_261_), .Y(_265_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[66]), .Y(_266_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__2_), .Y(_267_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__2_), .Y(_268_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_267_), .C(_268_), .Y(_269_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__2_), .Y(_270_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__2_), .Y(_271_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_270_), .C(bloque_bytes[66]), .Y(_272_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_272_), .C(_265_), .Y(_273_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[66]), .B(_271_), .C(_270_), .Y(_274_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_267_), .C(_266_), .Y(_275_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_258_), .C(_274_), .Y(_276_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_273_), .Y(_277_) );
XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_277_), .B(_264_), .Y(micro_ucr_hash1_b_4__6_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_275_), .C(_265_), .Y(_278_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_272_), .C(_258_), .Y(_279_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_279_), .Y(_280_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_264_), .C(_278_), .Y(_281_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[67]), .Y(_282_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__3_), .Y(_283_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__3_), .Y(_284_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_283_), .C(_282_), .Y(_285_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__3_), .Y(_286_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_2__3_), .Y(_287_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[67]), .B(_287_), .C(_286_), .Y(_288_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_288_), .C(_274_), .Y(_289_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_287_), .C(_286_), .Y(_290_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_283_), .C(bloque_bytes[67]), .Y(_291_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_290_), .C(_269_), .Y(_292_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_292_), .Y(_252_) );
XOR2X1 XOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_252_), .Y(micro_ucr_hash1_b_4__7_) );
XOR2X1 XOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_4__4_), .B(gnd), .Y(micro_ucr_hash1_a_4__0_) );
XOR2X1 XOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_4__5_), .B(gnd), .Y(micro_ucr_hash1_a_4__1_) );
XOR2X1 XOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_4__6_), .B(gnd), .Y(micro_ucr_hash1_a_4__2_) );
XOR2X1 XOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_4__7_), .B(gnd), .Y(micro_ucr_hash1_a_4__3_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[56]), .Y(_362_) );
XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__0_), .Y(_363_) );
XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_362_), .Y(micro_ucr_hash1_b_5__4_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_363_), .Y(_364_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__1_), .Y(_365_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__1_), .Y(_366_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[57]), .B(_366_), .C(_365_), .Y(_367_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[57]), .Y(_368_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__1_), .Y(_369_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__1_), .Y(_370_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_369_), .C(_368_), .Y(_371_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_367_), .Y(_372_) );
XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_364_), .Y(micro_ucr_hash1_b_5__5_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_367_), .B(_371_), .C(_364_), .Y(_373_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_368_), .B(_369_), .C(_370_), .Y(_374_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[58]), .Y(_375_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__2_), .Y(_376_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__2_), .Y(_377_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_376_), .C(_377_), .Y(_378_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__2_), .Y(_379_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__2_), .Y(_380_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_379_), .C(bloque_bytes[58]), .Y(_381_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_381_), .C(_374_), .Y(_382_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[58]), .B(_380_), .C(_379_), .Y(_383_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_376_), .C(_375_), .Y(_384_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_367_), .C(_383_), .Y(_385_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_382_), .Y(_386_) );
XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_386_), .B(_373_), .Y(micro_ucr_hash1_b_5__6_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_384_), .C(_374_), .Y(_387_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_381_), .C(_367_), .Y(_388_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_388_), .Y(_389_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_373_), .C(_387_), .Y(_390_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[59]), .Y(_391_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__3_), .Y(_392_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__3_), .Y(_393_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_392_), .C(_391_), .Y(_394_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__3_), .Y(_395_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_3__3_), .Y(_396_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[59]), .B(_396_), .C(_395_), .Y(_397_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_397_), .C(_383_), .Y(_398_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_391_), .B(_396_), .C(_395_), .Y(_399_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_392_), .C(bloque_bytes[59]), .Y(_400_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_400_), .B(_399_), .C(_378_), .Y(_401_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_401_), .Y(_293_) );
XOR2X1 XOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_293_), .Y(micro_ucr_hash1_b_5__7_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[60]), .Y(_294_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__4_), .B(micro_ucr_hash1_a_3__4_), .Y(_295_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__4_), .B(micro_ucr_hash1_a_3__4_), .Y(_296_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_296_), .C(_295_), .Y(_297_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__4_), .B(micro_ucr_hash1_a_3__4_), .Y(_298_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__4_), .B(micro_ucr_hash1_a_3__4_), .Y(_299_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_298_), .C(bloque_bytes[60]), .Y(_300_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_297_), .C(_300_), .Y(_301_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_395_), .C(bloque_bytes[59]), .Y(_302_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_298_), .C(_294_), .Y(_303_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[60]), .B(_296_), .C(_295_), .Y(_304_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_304_), .C(_302_), .Y(_305_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_305_), .B(_301_), .Y(_306_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(_401_), .Y(_307_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_378_), .Y(_308_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_308_), .C(_398_), .Y(_309_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_373_), .C(_309_), .Y(_310_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_310_), .Y(_311_) );
XNOR2X1 XNOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_306_), .Y(micro_ucr_hash1_c_4__4_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_305_), .Y(_312_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_312_), .C(_301_), .Y(_313_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[61]), .Y(_314_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__5_), .B(micro_ucr_hash1_a_3__5_), .Y(_315_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__5_), .B(micro_ucr_hash1_a_3__5_), .Y(_316_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_316_), .C(_315_), .Y(_317_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__5_), .B(micro_ucr_hash1_a_3__5_), .Y(_318_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__5_), .B(micro_ucr_hash1_a_3__5_), .Y(_319_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_318_), .C(bloque_bytes[61]), .Y(_320_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_320_), .C(_317_), .Y(_321_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_295_), .C(bloque_bytes[60]), .Y(_322_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[61]), .B(_316_), .C(_315_), .Y(_323_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_318_), .C(_314_), .Y(_324_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_323_), .C(_322_), .Y(_325_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_325_), .Y(_326_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(_326_), .Y(_327_) );
XNOR2X1 XNOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_327_), .Y(micro_ucr_hash1_c_4__5_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_325_), .C(_312_), .Y(_328_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_328_), .C(_310_), .Y(_329_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_323_), .Y(_330_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_322_), .Y(_331_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_331_), .Y(_332_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_330_), .C(_301_), .Y(_333_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_332_), .Y(_334_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[62]), .Y(_335_) );
XNOR2X1 XNOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__6_), .B(micro_ucr_hash1_a_3__6_), .Y(_336_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_335_), .Y(_337_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_335_), .B(_336_), .Y(_338_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_337_), .Y(_339_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_323_), .Y(_340_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_339_), .Y(_341_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_340_), .Y(_342_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_329_), .C(_342_), .Y(_343_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_306_), .Y(_344_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_344_), .C(_334_), .Y(_345_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_342_), .Y(_346_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_345_), .Y(_347_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_347_), .Y(micro_ucr_hash1_c_4__6_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_387_), .Y(_348_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_348_), .C(_398_), .Y(_349_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_363_), .C(_372_), .Y(_350_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_386_), .C(_293_), .Y(_351_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_351_), .C(_344_), .Y(_352_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_301_), .C(_331_), .Y(_353_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_353_), .C(_346_), .Y(_354_) );
XOR2X1 XOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__7_), .B(bloque_bytes[63]), .Y(_355_) );
XNOR2X1 XNOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(micro_ucr_hash1_a_3__7_), .Y(_356_) );
XNOR2X1 XNOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_356_), .B(_337_), .Y(_357_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_357_), .C(_354_), .Y(_358_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_340_), .Y(_359_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_357_), .Y(_360_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_359_), .C(_360_), .Y(_361_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_361_), .Y(micro_ucr_hash1_c_4__7_) );
XOR2X1 XOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__4_), .B(gnd), .Y(micro_ucr_hash1_a_5__0_) );
XOR2X1 XOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__5_), .B(gnd), .Y(micro_ucr_hash1_a_5__1_) );
XOR2X1 XOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__6_), .B(gnd), .Y(micro_ucr_hash1_a_5__2_) );
XOR2X1 XOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__7_), .B(gnd), .Y(micro_ucr_hash1_a_5__3_) );
XOR2X1 XOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_4__4_), .B(micro_ucr_hash1_b_4__4_), .Y(micro_ucr_hash1_a_5__4_) );
XOR2X1 XOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_4__5_), .B(micro_ucr_hash1_b_4__5_), .Y(micro_ucr_hash1_a_5__5_) );
XOR2X1 XOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_4__6_), .B(micro_ucr_hash1_b_4__6_), .Y(micro_ucr_hash1_a_5__6_) );
XOR2X1 XOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_4__7_), .B(micro_ucr_hash1_b_4__7_), .Y(micro_ucr_hash1_a_5__7_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[48]), .Y(_403_) );
XNOR2X1 XNOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__0_), .Y(_404_) );
XNOR2X1 XNOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_403_), .Y(micro_ucr_hash1_b_6__4_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_404_), .Y(_405_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__1_), .Y(_406_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__1_), .Y(_407_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[49]), .B(_407_), .C(_406_), .Y(_408_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[49]), .Y(_409_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__1_), .Y(_410_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__1_), .Y(_411_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_410_), .C(_409_), .Y(_412_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_408_), .Y(_413_) );
XNOR2X1 XNOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_405_), .Y(micro_ucr_hash1_b_6__5_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_412_), .C(_405_), .Y(_414_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_410_), .C(_411_), .Y(_415_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[50]), .Y(_416_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__2_), .Y(_417_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__2_), .Y(_418_) );
NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_417_), .C(_418_), .Y(_419_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__2_), .Y(_420_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__2_), .Y(_421_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_420_), .C(bloque_bytes[50]), .Y(_422_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_422_), .C(_415_), .Y(_423_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[50]), .B(_421_), .C(_420_), .Y(_424_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_417_), .C(_416_), .Y(_425_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_408_), .C(_424_), .Y(_426_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_426_), .B(_423_), .Y(_427_) );
XNOR2X1 XNOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_427_), .B(_414_), .Y(micro_ucr_hash1_b_6__6_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_425_), .C(_415_), .Y(_428_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_422_), .C(_408_), .Y(_429_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_429_), .Y(_430_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_414_), .C(_428_), .Y(_431_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[51]), .Y(_432_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__3_), .Y(_433_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__3_), .Y(_434_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_433_), .C(_432_), .Y(_435_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__3_), .Y(_436_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_4__3_), .Y(_437_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[51]), .B(_437_), .C(_436_), .Y(_438_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_438_), .C(_424_), .Y(_439_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_437_), .C(_436_), .Y(_440_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_433_), .C(bloque_bytes[51]), .Y(_441_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_440_), .C(_419_), .Y(_442_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_442_), .Y(_402_) );
XOR2X1 XOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_402_), .Y(micro_ucr_hash1_b_6__7_) );
XOR2X1 XOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_6__4_), .B(gnd), .Y(micro_ucr_hash1_a_6__0_) );
XOR2X1 XOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_6__5_), .B(gnd), .Y(micro_ucr_hash1_a_6__1_) );
XOR2X1 XOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_6__6_), .B(gnd), .Y(micro_ucr_hash1_a_6__2_) );
XOR2X1 XOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_6__7_), .B(gnd), .Y(micro_ucr_hash1_a_6__3_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[40]), .Y(_512_) );
XNOR2X1 XNOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__0_), .Y(_513_) );
XNOR2X1 XNOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_512_), .Y(micro_ucr_hash1_b_7__4_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_513_), .Y(_514_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__1_), .Y(_515_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__1_), .Y(_516_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[41]), .B(_516_), .C(_515_), .Y(_517_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[41]), .Y(_518_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__1_), .Y(_519_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__1_), .Y(_520_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_519_), .C(_518_), .Y(_521_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_517_), .Y(_522_) );
XNOR2X1 XNOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_514_), .Y(micro_ucr_hash1_b_7__5_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(_521_), .C(_514_), .Y(_523_) );
NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_518_), .B(_519_), .C(_520_), .Y(_524_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[42]), .Y(_525_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__2_), .Y(_526_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__2_), .Y(_527_) );
NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_526_), .C(_527_), .Y(_528_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__2_), .Y(_529_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__2_), .Y(_530_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_530_), .B(_529_), .C(bloque_bytes[42]), .Y(_531_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_531_), .C(_524_), .Y(_532_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[42]), .B(_530_), .C(_529_), .Y(_533_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_527_), .B(_526_), .C(_525_), .Y(_534_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_517_), .C(_533_), .Y(_535_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_535_), .B(_532_), .Y(_536_) );
XNOR2X1 XNOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_523_), .Y(micro_ucr_hash1_b_7__6_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_533_), .B(_534_), .C(_524_), .Y(_537_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_528_), .B(_531_), .C(_517_), .Y(_538_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_538_), .Y(_539_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_523_), .C(_537_), .Y(_540_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[43]), .Y(_541_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__3_), .Y(_542_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__3_), .Y(_543_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_542_), .C(_541_), .Y(_544_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__3_), .Y(_545_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_5__3_), .Y(_546_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[43]), .B(_546_), .C(_545_), .Y(_547_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_547_), .C(_533_), .Y(_548_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_541_), .B(_546_), .C(_545_), .Y(_549_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_542_), .C(bloque_bytes[43]), .Y(_550_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_549_), .C(_528_), .Y(_551_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_551_), .Y(_443_) );
XOR2X1 XOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_443_), .Y(micro_ucr_hash1_b_7__7_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[44]), .Y(_444_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__4_), .B(micro_ucr_hash1_a_5__4_), .Y(_445_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__4_), .B(micro_ucr_hash1_a_5__4_), .Y(_446_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_446_), .C(_445_), .Y(_447_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__4_), .B(micro_ucr_hash1_a_5__4_), .Y(_448_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__4_), .B(micro_ucr_hash1_a_5__4_), .Y(_449_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_448_), .C(bloque_bytes[44]), .Y(_450_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_447_), .C(_450_), .Y(_451_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_546_), .B(_545_), .C(bloque_bytes[43]), .Y(_452_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_448_), .C(_444_), .Y(_453_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[44]), .B(_446_), .C(_445_), .Y(_454_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_454_), .C(_452_), .Y(_455_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_451_), .Y(_456_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(_551_), .Y(_457_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_528_), .Y(_458_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_524_), .B(_458_), .C(_548_), .Y(_459_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_523_), .C(_459_), .Y(_460_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_460_), .Y(_461_) );
XNOR2X1 XNOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_456_), .Y(micro_ucr_hash1_c_6__4_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_455_), .Y(_462_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_462_), .C(_451_), .Y(_463_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[45]), .Y(_464_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__5_), .B(micro_ucr_hash1_a_5__5_), .Y(_465_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__5_), .B(micro_ucr_hash1_a_5__5_), .Y(_466_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_466_), .C(_465_), .Y(_467_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__5_), .B(micro_ucr_hash1_a_5__5_), .Y(_468_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__5_), .B(micro_ucr_hash1_a_5__5_), .Y(_469_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_468_), .C(bloque_bytes[45]), .Y(_470_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_470_), .C(_467_), .Y(_471_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_446_), .B(_445_), .C(bloque_bytes[44]), .Y(_472_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[45]), .B(_466_), .C(_465_), .Y(_473_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_468_), .C(_464_), .Y(_474_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_473_), .C(_472_), .Y(_475_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_475_), .Y(_476_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(_476_), .Y(_477_) );
XNOR2X1 XNOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_477_), .Y(micro_ucr_hash1_c_6__5_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_471_), .B(_475_), .C(_462_), .Y(_478_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_478_), .C(_460_), .Y(_479_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_473_), .Y(_480_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_472_), .Y(_481_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_481_), .Y(_482_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_480_), .C(_451_), .Y(_483_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_482_), .Y(_484_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[46]), .Y(_485_) );
XNOR2X1 XNOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__6_), .B(micro_ucr_hash1_a_5__6_), .Y(_486_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_485_), .Y(_487_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_486_), .Y(_488_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_487_), .Y(_489_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_473_), .Y(_490_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_473_), .B(_489_), .Y(_491_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_490_), .Y(_492_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_479_), .C(_492_), .Y(_493_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_456_), .Y(_494_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_494_), .C(_484_), .Y(_495_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_492_), .Y(_496_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_496_), .B(_495_), .Y(_497_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_497_), .Y(micro_ucr_hash1_c_6__6_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_537_), .Y(_498_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_498_), .C(_548_), .Y(_499_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_513_), .C(_522_), .Y(_500_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_536_), .C(_443_), .Y(_501_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_499_), .B(_501_), .C(_494_), .Y(_502_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_477_), .B(_451_), .C(_481_), .Y(_503_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_503_), .C(_496_), .Y(_504_) );
XOR2X1 XOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__7_), .B(bloque_bytes[47]), .Y(_505_) );
XNOR2X1 XNOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_505_), .B(micro_ucr_hash1_a_5__7_), .Y(_506_) );
XNOR2X1 XNOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_487_), .Y(_507_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_507_), .C(_504_), .Y(_508_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_490_), .Y(_509_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_507_), .Y(_510_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_509_), .C(_510_), .Y(_511_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_511_), .Y(micro_ucr_hash1_c_6__7_) );
XOR2X1 XOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__4_), .B(gnd), .Y(micro_ucr_hash1_a_7__0_) );
XOR2X1 XOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__5_), .B(gnd), .Y(micro_ucr_hash1_a_7__1_) );
XOR2X1 XOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__6_), .B(gnd), .Y(micro_ucr_hash1_a_7__2_) );
XOR2X1 XOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__7_), .B(gnd), .Y(micro_ucr_hash1_a_7__3_) );
XOR2X1 XOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_6__4_), .B(micro_ucr_hash1_b_6__4_), .Y(micro_ucr_hash1_a_7__4_) );
XOR2X1 XOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_6__5_), .B(micro_ucr_hash1_b_6__5_), .Y(micro_ucr_hash1_a_7__5_) );
XOR2X1 XOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_6__6_), .B(micro_ucr_hash1_b_6__6_), .Y(micro_ucr_hash1_a_7__6_) );
XOR2X1 XOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_6__7_), .B(micro_ucr_hash1_b_6__7_), .Y(micro_ucr_hash1_a_7__7_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[32]), .Y(_553_) );
XNOR2X1 XNOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__0_), .Y(_554_) );
XNOR2X1 XNOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_554_), .B(_553_), .Y(micro_ucr_hash1_b_8__4_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_554_), .Y(_555_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__1_), .Y(_556_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__1_), .Y(_557_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[33]), .B(_557_), .C(_556_), .Y(_558_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[33]), .Y(_559_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__1_), .Y(_560_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__1_), .Y(_561_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_560_), .C(_559_), .Y(_562_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_562_), .B(_558_), .Y(_563_) );
XNOR2X1 XNOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_563_), .B(_555_), .Y(micro_ucr_hash1_b_8__5_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_562_), .C(_555_), .Y(_564_) );
NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_559_), .B(_560_), .C(_561_), .Y(_565_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[34]), .Y(_566_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__2_), .Y(_567_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__2_), .Y(_568_) );
NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_566_), .B(_567_), .C(_568_), .Y(_569_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__2_), .Y(_570_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__2_), .Y(_571_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_570_), .C(bloque_bytes[34]), .Y(_572_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_572_), .C(_565_), .Y(_573_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[34]), .B(_571_), .C(_570_), .Y(_574_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_568_), .B(_567_), .C(_566_), .Y(_575_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_575_), .B(_558_), .C(_574_), .Y(_576_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_573_), .Y(_577_) );
XNOR2X1 XNOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_564_), .Y(micro_ucr_hash1_b_8__6_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_575_), .C(_565_), .Y(_578_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_569_), .B(_572_), .C(_558_), .Y(_579_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_578_), .B(_579_), .Y(_580_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_564_), .C(_578_), .Y(_581_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[35]), .Y(_582_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__3_), .Y(_583_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__3_), .Y(_584_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_583_), .C(_582_), .Y(_585_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__3_), .Y(_586_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_6__3_), .Y(_587_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[35]), .B(_587_), .C(_586_), .Y(_588_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_585_), .B(_588_), .C(_574_), .Y(_589_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_587_), .C(_586_), .Y(_590_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_584_), .B(_583_), .C(bloque_bytes[35]), .Y(_591_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_591_), .B(_590_), .C(_569_), .Y(_592_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_589_), .B(_592_), .Y(_552_) );
XOR2X1 XOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_552_), .Y(micro_ucr_hash1_b_8__7_) );
XOR2X1 XOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_8__4_), .B(gnd), .Y(micro_ucr_hash1_a_8__0_) );
XOR2X1 XOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_8__5_), .B(gnd), .Y(micro_ucr_hash1_a_8__1_) );
XOR2X1 XOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_8__6_), .B(gnd), .Y(micro_ucr_hash1_a_8__2_) );
XOR2X1 XOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_8__7_), .B(gnd), .Y(micro_ucr_hash1_a_8__3_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[24]), .Y(_662_) );
XNOR2X1 XNOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__0_), .Y(_663_) );
XNOR2X1 XNOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_662_), .Y(micro_ucr_hash1_b_9__4_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_663_), .Y(_664_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__1_), .Y(_665_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__1_), .Y(_666_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[25]), .B(_666_), .C(_665_), .Y(_667_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[25]), .Y(_668_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__1_), .Y(_669_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__1_), .Y(_670_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_670_), .B(_669_), .C(_668_), .Y(_671_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_671_), .B(_667_), .Y(_672_) );
XNOR2X1 XNOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_664_), .Y(micro_ucr_hash1_b_9__5_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_667_), .B(_671_), .C(_664_), .Y(_673_) );
NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_669_), .C(_670_), .Y(_674_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[26]), .Y(_675_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__2_), .Y(_676_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__2_), .Y(_677_) );
NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_675_), .B(_676_), .C(_677_), .Y(_678_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__2_), .Y(_679_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__2_), .Y(_680_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_680_), .B(_679_), .C(bloque_bytes[26]), .Y(_681_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_681_), .C(_674_), .Y(_682_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[26]), .B(_680_), .C(_679_), .Y(_683_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_677_), .B(_676_), .C(_675_), .Y(_684_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_667_), .C(_683_), .Y(_685_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_682_), .Y(_686_) );
XNOR2X1 XNOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_686_), .B(_673_), .Y(micro_ucr_hash1_b_9__6_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_683_), .B(_684_), .C(_674_), .Y(_687_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_681_), .C(_667_), .Y(_688_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_688_), .Y(_689_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_673_), .C(_687_), .Y(_690_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[27]), .Y(_691_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__3_), .Y(_692_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__3_), .Y(_693_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_692_), .C(_691_), .Y(_694_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__3_), .Y(_695_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_7__3_), .Y(_696_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[27]), .B(_696_), .C(_695_), .Y(_697_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_697_), .C(_683_), .Y(_698_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_691_), .B(_696_), .C(_695_), .Y(_699_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_692_), .C(bloque_bytes[27]), .Y(_700_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_699_), .C(_678_), .Y(_701_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_698_), .B(_701_), .Y(_593_) );
XOR2X1 XOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(_593_), .Y(micro_ucr_hash1_b_9__7_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[28]), .Y(_594_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__4_), .B(micro_ucr_hash1_a_7__4_), .Y(_595_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__4_), .B(micro_ucr_hash1_a_7__4_), .Y(_596_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_596_), .C(_595_), .Y(_597_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__4_), .B(micro_ucr_hash1_a_7__4_), .Y(_598_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__4_), .B(micro_ucr_hash1_a_7__4_), .Y(_599_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(_598_), .C(bloque_bytes[28]), .Y(_600_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_694_), .B(_597_), .C(_600_), .Y(_601_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_695_), .C(bloque_bytes[27]), .Y(_602_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(_598_), .C(_594_), .Y(_603_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[28]), .B(_596_), .C(_595_), .Y(_604_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_604_), .C(_602_), .Y(_605_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_605_), .B(_601_), .Y(_606_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(_701_), .Y(_607_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_681_), .B(_678_), .Y(_608_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_674_), .B(_608_), .C(_698_), .Y(_609_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_673_), .C(_609_), .Y(_610_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_610_), .Y(_611_) );
XNOR2X1 XNOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_606_), .Y(micro_ucr_hash1_c_8__4_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_601_), .B(_605_), .Y(_612_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_612_), .C(_601_), .Y(_613_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[29]), .Y(_614_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__5_), .B(micro_ucr_hash1_a_7__5_), .Y(_615_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__5_), .B(micro_ucr_hash1_a_7__5_), .Y(_616_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_616_), .C(_615_), .Y(_617_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__5_), .B(micro_ucr_hash1_a_7__5_), .Y(_618_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__5_), .B(micro_ucr_hash1_a_7__5_), .Y(_619_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_618_), .C(bloque_bytes[29]), .Y(_620_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_620_), .C(_617_), .Y(_621_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_595_), .C(bloque_bytes[28]), .Y(_622_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[29]), .B(_616_), .C(_615_), .Y(_623_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_618_), .C(_614_), .Y(_624_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_623_), .C(_622_), .Y(_625_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_625_), .Y(_626_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(_626_), .Y(_627_) );
XNOR2X1 XNOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_613_), .B(_627_), .Y(micro_ucr_hash1_c_8__5_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_621_), .B(_625_), .C(_612_), .Y(_628_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_628_), .C(_610_), .Y(_629_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_624_), .B(_623_), .Y(_630_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_630_), .B(_622_), .Y(_631_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_631_), .Y(_632_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_622_), .B(_630_), .C(_601_), .Y(_633_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_633_), .B(_632_), .Y(_634_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[30]), .Y(_635_) );
XNOR2X1 XNOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__6_), .B(micro_ucr_hash1_a_7__6_), .Y(_636_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_636_), .B(_635_), .Y(_637_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_636_), .Y(_638_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_637_), .Y(_639_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_639_), .B(_623_), .Y(_640_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(_639_), .Y(_641_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_640_), .Y(_642_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_634_), .B(_629_), .C(_642_), .Y(_643_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_626_), .B(_606_), .Y(_644_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_644_), .C(_634_), .Y(_645_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(_642_), .Y(_646_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_646_), .B(_645_), .Y(_647_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_647_), .Y(micro_ucr_hash1_c_8__6_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_687_), .Y(_648_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_648_), .C(_698_), .Y(_649_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_662_), .B(_663_), .C(_672_), .Y(_650_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_686_), .C(_593_), .Y(_651_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_649_), .B(_651_), .C(_644_), .Y(_652_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_601_), .C(_631_), .Y(_653_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_652_), .B(_653_), .C(_646_), .Y(_654_) );
XOR2X1 XOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__7_), .B(bloque_bytes[31]), .Y(_655_) );
XNOR2X1 XNOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(micro_ucr_hash1_a_7__7_), .Y(_656_) );
XNOR2X1 XNOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_656_), .B(_637_), .Y(_657_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_640_), .B(_657_), .C(_654_), .Y(_658_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_640_), .Y(_659_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_657_), .Y(_660_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_643_), .B(_659_), .C(_660_), .Y(_661_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_661_), .Y(micro_ucr_hash1_c_8__7_) );
XOR2X1 XOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__4_), .B(gnd), .Y(micro_ucr_hash1_a_9__0_) );
XOR2X1 XOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__5_), .B(gnd), .Y(micro_ucr_hash1_a_9__1_) );
XOR2X1 XOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__6_), .B(gnd), .Y(micro_ucr_hash1_a_9__2_) );
XOR2X1 XOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__7_), .B(gnd), .Y(micro_ucr_hash1_a_9__3_) );
XOR2X1 XOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_8__4_), .B(micro_ucr_hash1_b_8__4_), .Y(micro_ucr_hash1_a_9__4_) );
XOR2X1 XOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_8__5_), .B(micro_ucr_hash1_b_8__5_), .Y(micro_ucr_hash1_a_9__5_) );
XOR2X1 XOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_8__6_), .B(micro_ucr_hash1_b_8__6_), .Y(micro_ucr_hash1_a_9__6_) );
XOR2X1 XOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_8__7_), .B(micro_ucr_hash1_b_8__7_), .Y(micro_ucr_hash1_a_9__7_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[16]), .Y(_703_) );
XNOR2X1 XNOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__0_), .Y(_704_) );
XNOR2X1 XNOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_703_), .Y(micro_ucr_hash1_b_10__4_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_704_), .Y(_705_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__1_), .Y(_706_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__1_), .Y(_707_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[17]), .B(_707_), .C(_706_), .Y(_708_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[17]), .Y(_709_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__1_), .Y(_710_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__1_), .Y(_711_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_710_), .C(_709_), .Y(_712_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_712_), .B(_708_), .Y(_713_) );
XNOR2X1 XNOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_705_), .Y(micro_ucr_hash1_b_10__5_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_712_), .C(_705_), .Y(_714_) );
NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_710_), .C(_711_), .Y(_715_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[18]), .Y(_716_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__2_), .Y(_717_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__2_), .Y(_718_) );
NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_717_), .C(_718_), .Y(_719_) );
OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__2_), .Y(_720_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__2_), .Y(_721_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_721_), .B(_720_), .C(bloque_bytes[18]), .Y(_722_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_722_), .C(_715_), .Y(_723_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[18]), .B(_721_), .C(_720_), .Y(_724_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_717_), .C(_716_), .Y(_725_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(_725_), .B(_708_), .C(_724_), .Y(_726_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_723_), .Y(_727_) );
XNOR2X1 XNOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_714_), .Y(micro_ucr_hash1_b_10__6_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_725_), .C(_715_), .Y(_728_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_722_), .C(_708_), .Y(_729_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_728_), .B(_729_), .Y(_730_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_730_), .B(_714_), .C(_728_), .Y(_731_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[19]), .Y(_732_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__3_), .Y(_733_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__3_), .Y(_734_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_733_), .C(_732_), .Y(_735_) );
OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__3_), .Y(_736_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_8__3_), .Y(_737_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[19]), .B(_737_), .C(_736_), .Y(_738_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_735_), .B(_738_), .C(_724_), .Y(_739_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_737_), .C(_736_), .Y(_740_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_733_), .C(bloque_bytes[19]), .Y(_741_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_740_), .C(_719_), .Y(_742_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_742_), .Y(_702_) );
XOR2X1 XOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_731_), .B(_702_), .Y(micro_ucr_hash1_b_10__7_) );
XOR2X1 XOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_10__4_), .B(gnd), .Y(micro_ucr_hash1_a_10__0_) );
XOR2X1 XOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_10__5_), .B(gnd), .Y(micro_ucr_hash1_a_10__1_) );
XOR2X1 XOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_10__6_), .B(gnd), .Y(micro_ucr_hash1_a_10__2_) );
XOR2X1 XOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_10__7_), .B(gnd), .Y(micro_ucr_hash1_a_10__3_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[8]), .Y(_812_) );
XNOR2X1 XNOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__0_), .Y(_813_) );
XNOR2X1 XNOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_813_), .B(_812_), .Y(micro_ucr_hash1_b_11__4_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_813_), .Y(_814_) );
OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__1_), .Y(_815_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__1_), .Y(_816_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[9]), .B(_816_), .C(_815_), .Y(_817_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[9]), .Y(_818_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__1_), .Y(_819_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__1_), .Y(_820_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_820_), .B(_819_), .C(_818_), .Y(_821_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_821_), .B(_817_), .Y(_822_) );
XNOR2X1 XNOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_822_), .B(_814_), .Y(micro_ucr_hash1_b_11__5_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_817_), .B(_821_), .C(_814_), .Y(_823_) );
NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_819_), .C(_820_), .Y(_824_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[10]), .Y(_825_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__2_), .Y(_826_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__2_), .Y(_827_) );
NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_826_), .C(_827_), .Y(_828_) );
OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__2_), .Y(_829_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__2_), .Y(_830_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_830_), .B(_829_), .C(bloque_bytes[10]), .Y(_831_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_828_), .B(_831_), .C(_824_), .Y(_832_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[10]), .B(_830_), .C(_829_), .Y(_833_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_827_), .B(_826_), .C(_825_), .Y(_834_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_834_), .B(_817_), .C(_833_), .Y(_835_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_835_), .B(_832_), .Y(_836_) );
XNOR2X1 XNOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_836_), .B(_823_), .Y(micro_ucr_hash1_b_11__6_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_833_), .B(_834_), .C(_824_), .Y(_837_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_828_), .B(_831_), .C(_817_), .Y(_838_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_837_), .B(_838_), .Y(_839_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_823_), .C(_837_), .Y(_840_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[11]), .Y(_841_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__3_), .Y(_842_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__3_), .Y(_843_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_842_), .C(_841_), .Y(_844_) );
OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__3_), .Y(_845_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_9__3_), .Y(_846_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[11]), .B(_846_), .C(_845_), .Y(_847_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_847_), .C(_833_), .Y(_848_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_841_), .B(_846_), .C(_845_), .Y(_849_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_842_), .C(bloque_bytes[11]), .Y(_850_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_850_), .B(_849_), .C(_828_), .Y(_851_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_848_), .B(_851_), .Y(_743_) );
XOR2X1 XOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_743_), .Y(micro_ucr_hash1_b_11__7_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[12]), .Y(_744_) );
OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__4_), .B(micro_ucr_hash1_a_9__4_), .Y(_745_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__4_), .B(micro_ucr_hash1_a_9__4_), .Y(_746_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(_744_), .B(_746_), .C(_745_), .Y(_747_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__4_), .B(micro_ucr_hash1_a_9__4_), .Y(_748_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__4_), .B(micro_ucr_hash1_a_9__4_), .Y(_749_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_748_), .C(bloque_bytes[12]), .Y(_750_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_747_), .C(_750_), .Y(_751_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_845_), .C(bloque_bytes[11]), .Y(_752_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_749_), .B(_748_), .C(_744_), .Y(_753_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[12]), .B(_746_), .C(_745_), .Y(_754_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_754_), .C(_752_), .Y(_755_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_751_), .Y(_756_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(_851_), .Y(_757_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_831_), .B(_828_), .Y(_758_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_758_), .C(_848_), .Y(_759_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_839_), .B(_823_), .C(_759_), .Y(_760_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_760_), .Y(_761_) );
XNOR2X1 XNOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_756_), .Y(micro_ucr_hash1_c_10__4_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_751_), .B(_755_), .Y(_762_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_762_), .C(_751_), .Y(_763_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[13]), .Y(_764_) );
OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__5_), .B(micro_ucr_hash1_a_9__5_), .Y(_765_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__5_), .B(micro_ucr_hash1_a_9__5_), .Y(_766_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(_766_), .C(_765_), .Y(_767_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__5_), .B(micro_ucr_hash1_a_9__5_), .Y(_768_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__5_), .B(micro_ucr_hash1_a_9__5_), .Y(_769_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_768_), .C(bloque_bytes[13]), .Y(_770_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_753_), .B(_770_), .C(_767_), .Y(_771_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_746_), .B(_745_), .C(bloque_bytes[12]), .Y(_772_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[13]), .B(_766_), .C(_765_), .Y(_773_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_768_), .C(_764_), .Y(_774_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_774_), .B(_773_), .C(_772_), .Y(_775_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_775_), .Y(_776_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(_776_), .Y(_777_) );
XNOR2X1 XNOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_777_), .Y(micro_ucr_hash1_c_10__5_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_771_), .B(_775_), .C(_762_), .Y(_778_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_778_), .C(_760_), .Y(_779_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_774_), .B(_773_), .Y(_780_) );
OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_780_), .B(_772_), .Y(_781_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_781_), .Y(_782_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_780_), .C(_751_), .Y(_783_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_782_), .Y(_784_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[14]), .Y(_785_) );
XNOR2X1 XNOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__6_), .B(micro_ucr_hash1_a_9__6_), .Y(_786_) );
OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_785_), .Y(_787_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_786_), .Y(_788_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_787_), .Y(_789_) );
OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_773_), .Y(_790_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_773_), .B(_789_), .Y(_791_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_791_), .B(_790_), .Y(_792_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_784_), .B(_779_), .C(_792_), .Y(_793_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_776_), .B(_756_), .Y(_794_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_761_), .B(_794_), .C(_784_), .Y(_795_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_792_), .Y(_796_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_795_), .Y(_797_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_797_), .Y(micro_ucr_hash1_c_10__6_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(_837_), .Y(_798_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_757_), .B(_798_), .C(_848_), .Y(_799_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_813_), .C(_822_), .Y(_800_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_836_), .C(_743_), .Y(_801_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_799_), .B(_801_), .C(_794_), .Y(_802_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_777_), .B(_751_), .C(_781_), .Y(_803_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_803_), .C(_796_), .Y(_804_) );
XOR2X1 XOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__7_), .B(bloque_bytes[15]), .Y(_805_) );
XNOR2X1 XNOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(micro_ucr_hash1_a_9__7_), .Y(_806_) );
XNOR2X1 XNOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_787_), .Y(_807_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_807_), .C(_804_), .Y(_808_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(_790_), .Y(_809_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_807_), .Y(_810_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_809_), .C(_810_), .Y(_811_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_808_), .B(_811_), .Y(micro_ucr_hash1_c_10__7_) );
XOR2X1 XOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__4_), .B(gnd), .Y(micro_ucr_hash1_a_11__0_) );
XOR2X1 XOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__5_), .B(gnd), .Y(micro_ucr_hash1_a_11__1_) );
XOR2X1 XOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__6_), .B(gnd), .Y(micro_ucr_hash1_a_11__2_) );
XOR2X1 XOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__7_), .B(gnd), .Y(micro_ucr_hash1_a_11__3_) );
XOR2X1 XOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_10__4_), .B(micro_ucr_hash1_b_10__4_), .Y(micro_ucr_hash1_a_11__4_) );
XOR2X1 XOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_10__5_), .B(micro_ucr_hash1_b_10__5_), .Y(micro_ucr_hash1_a_11__5_) );
XOR2X1 XOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_10__6_), .B(micro_ucr_hash1_b_10__6_), .Y(micro_ucr_hash1_a_11__6_) );
XOR2X1 XOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_10__7_), .B(micro_ucr_hash1_b_10__7_), .Y(micro_ucr_hash1_a_11__7_) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[0]), .Y(_853_) );
XNOR2X1 XNOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__0_), .Y(_854_) );
XNOR2X1 XNOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_854_), .B(_853_), .Y(micro_ucr_hash1_b_12__4_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_854_), .Y(_855_) );
OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__1_), .Y(_856_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__1_), .Y(_857_) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[1]), .B(_857_), .C(_856_), .Y(_858_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[1]), .Y(_859_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__1_), .Y(_860_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__1_), .Y(_861_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_861_), .B(_860_), .C(_859_), .Y(_862_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_858_), .Y(_863_) );
XNOR2X1 XNOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_863_), .B(_855_), .Y(micro_ucr_hash1_b_12__5_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_862_), .C(_855_), .Y(_864_) );
NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_859_), .B(_860_), .C(_861_), .Y(_865_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[2]), .Y(_866_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__2_), .Y(_867_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__2_), .Y(_868_) );
NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_866_), .B(_867_), .C(_868_), .Y(_869_) );
OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__2_), .Y(_870_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__2_), .Y(_871_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_871_), .B(_870_), .C(bloque_bytes[2]), .Y(_872_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_872_), .C(_865_), .Y(_873_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[2]), .B(_871_), .C(_870_), .Y(_874_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_867_), .C(_866_), .Y(_875_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_875_), .B(_858_), .C(_874_), .Y(_876_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_876_), .B(_873_), .Y(_877_) );
XNOR2X1 XNOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_877_), .B(_864_), .Y(micro_ucr_hash1_b_12__6_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_874_), .B(_875_), .C(_865_), .Y(_878_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_872_), .C(_858_), .Y(_879_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_878_), .B(_879_), .Y(_880_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_880_), .B(_864_), .C(_878_), .Y(_881_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[3]), .Y(_882_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__3_), .Y(_883_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__3_), .Y(_884_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_884_), .B(_883_), .C(_882_), .Y(_885_) );
OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__3_), .Y(_886_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_10__3_), .Y(_887_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[3]), .B(_887_), .C(_886_), .Y(_888_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_885_), .B(_888_), .C(_874_), .Y(_889_) );
NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_882_), .B(_887_), .C(_886_), .Y(_890_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_884_), .B(_883_), .C(bloque_bytes[3]), .Y(_891_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_890_), .C(_869_), .Y(_892_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_889_), .B(_892_), .Y(_852_) );
XOR2X1 XOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_852_), .Y(micro_ucr_hash1_b_12__7_) );
XOR2X1 XOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_12__4_), .B(gnd), .Y(micro_ucr_hash1_a_12__0_) );
XOR2X1 XOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_12__5_), .B(gnd), .Y(micro_ucr_hash1_a_12__1_) );
XOR2X1 XOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_12__6_), .B(gnd), .Y(micro_ucr_hash1_a_12__2_) );
XOR2X1 XOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_12__7_), .B(gnd), .Y(micro_ucr_hash1_a_12__3_) );
INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_24_), .Y(_962_) );
XNOR2X1 XNOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__0_), .Y(_963_) );
XNOR2X1 XNOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_963_), .B(_962_), .Y(micro_ucr_hash1_b_13__4_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_963_), .Y(_964_) );
OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__1_), .Y(_965_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__1_), .Y(_966_) );
NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_25_), .B(_966_), .C(_965_), .Y(_967_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_25_), .Y(_968_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__1_), .Y(_969_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__1_), .Y(_970_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_970_), .B(_969_), .C(_968_), .Y(_971_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_967_), .Y(_972_) );
XNOR2X1 XNOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_964_), .Y(micro_ucr_hash1_b_13__5_) );
NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_967_), .B(_971_), .C(_964_), .Y(_973_) );
NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_969_), .C(_970_), .Y(_974_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_26_), .Y(_975_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__2_), .Y(_976_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__2_), .Y(_977_) );
NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_976_), .C(_977_), .Y(_978_) );
OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__2_), .Y(_979_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__2_), .Y(_980_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_980_), .B(_979_), .C(entrada_hash1_nonce_26_), .Y(_981_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_981_), .C(_974_), .Y(_982_) );
NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_26_), .B(_980_), .C(_979_), .Y(_983_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_977_), .B(_976_), .C(_975_), .Y(_984_) );
NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_984_), .B(_967_), .C(_983_), .Y(_985_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_985_), .B(_982_), .Y(_986_) );
XNOR2X1 XNOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_986_), .B(_973_), .Y(micro_ucr_hash1_b_13__6_) );
NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_983_), .B(_984_), .C(_974_), .Y(_987_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_978_), .B(_981_), .C(_967_), .Y(_988_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_987_), .B(_988_), .Y(_989_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_973_), .C(_987_), .Y(_990_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_27_), .Y(_991_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__3_), .Y(_992_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__3_), .Y(_993_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_992_), .C(_991_), .Y(_994_) );
OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__3_), .Y(_995_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_11__3_), .Y(_996_) );
NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_27_), .B(_996_), .C(_995_), .Y(_997_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_997_), .C(_983_), .Y(_998_) );
NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_991_), .B(_996_), .C(_995_), .Y(_999_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_992_), .C(entrada_hash1_nonce_27_), .Y(_1000_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_999_), .C(_978_), .Y(_1001_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_1001_), .Y(_893_) );
XOR2X1 XOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_893_), .Y(micro_ucr_hash1_b_13__7_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_28_), .Y(_894_) );
OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__4_), .B(micro_ucr_hash1_a_11__4_), .Y(_895_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__4_), .B(micro_ucr_hash1_a_11__4_), .Y(_896_) );
NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_896_), .C(_895_), .Y(_897_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__4_), .B(micro_ucr_hash1_a_11__4_), .Y(_898_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__4_), .B(micro_ucr_hash1_a_11__4_), .Y(_899_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_899_), .B(_898_), .C(entrada_hash1_nonce_28_), .Y(_900_) );
NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_994_), .B(_897_), .C(_900_), .Y(_901_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_995_), .C(entrada_hash1_nonce_27_), .Y(_902_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_899_), .B(_898_), .C(_894_), .Y(_903_) );
NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_28_), .B(_896_), .C(_895_), .Y(_904_) );
NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_904_), .C(_902_), .Y(_905_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_901_), .Y(_906_) );
INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .Y(_907_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_981_), .B(_978_), .Y(_908_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_974_), .B(_908_), .C(_998_), .Y(_909_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_973_), .C(_909_), .Y(_910_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_910_), .Y(_911_) );
XNOR2X1 XNOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_906_), .Y(micro_ucr_hash1_c_12__4_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_905_), .Y(_912_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_912_), .C(_901_), .Y(_913_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_29_), .Y(_914_) );
OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__5_), .B(micro_ucr_hash1_a_11__5_), .Y(_915_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__5_), .B(micro_ucr_hash1_a_11__5_), .Y(_916_) );
NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_916_), .C(_915_), .Y(_917_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__5_), .B(micro_ucr_hash1_a_11__5_), .Y(_918_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__5_), .B(micro_ucr_hash1_a_11__5_), .Y(_919_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_918_), .C(entrada_hash1_nonce_29_), .Y(_920_) );
NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_920_), .C(_917_), .Y(_921_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_896_), .B(_895_), .C(entrada_hash1_nonce_28_), .Y(_922_) );
NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_29_), .B(_916_), .C(_915_), .Y(_923_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_918_), .C(_914_), .Y(_924_) );
NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_923_), .C(_922_), .Y(_925_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_921_), .B(_925_), .Y(_926_) );
INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(_926_), .Y(_927_) );
XNOR2X1 XNOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_913_), .B(_927_), .Y(micro_ucr_hash1_c_12__5_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_921_), .B(_925_), .C(_912_), .Y(_928_) );
NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_928_), .C(_910_), .Y(_929_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_923_), .Y(_930_) );
OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_930_), .B(_922_), .Y(_931_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_931_), .Y(_932_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_930_), .C(_901_), .Y(_933_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_933_), .B(_932_), .Y(_934_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_30_), .Y(_935_) );
XNOR2X1 XNOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__6_), .B(micro_ucr_hash1_a_11__6_), .Y(_936_) );
OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_935_), .Y(_937_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_936_), .Y(_938_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_937_), .Y(_939_) );
OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(_923_), .Y(_940_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_923_), .B(_939_), .Y(_941_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_940_), .Y(_942_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_929_), .C(_942_), .Y(_943_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_926_), .B(_906_), .Y(_944_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_944_), .C(_934_), .Y(_945_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_942_), .Y(_946_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_946_), .B(_945_), .Y(_947_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_943_), .B(_947_), .Y(micro_ucr_hash1_c_12__6_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_987_), .Y(_948_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_948_), .C(_998_), .Y(_949_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_963_), .C(_972_), .Y(_950_) );
NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(_950_), .B(_986_), .C(_893_), .Y(_951_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_951_), .C(_944_), .Y(_952_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_927_), .B(_901_), .C(_931_), .Y(_953_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_952_), .B(_953_), .C(_946_), .Y(_954_) );
XOR2X1 XOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__7_), .B(entrada_hash1_nonce_31_), .Y(_955_) );
XNOR2X1 XNOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(micro_ucr_hash1_a_11__7_), .Y(_956_) );
XNOR2X1 XNOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_956_), .B(_937_), .Y(_957_) );
NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_940_), .B(_957_), .C(_954_), .Y(_958_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_940_), .Y(_959_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_957_), .Y(_960_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_943_), .B(_959_), .C(_960_), .Y(_961_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_958_), .B(_961_), .Y(micro_ucr_hash1_c_12__7_) );
XOR2X1 XOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__4_), .B(gnd), .Y(micro_ucr_hash1_a_13__0_) );
XOR2X1 XOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__5_), .B(gnd), .Y(micro_ucr_hash1_a_13__1_) );
XOR2X1 XOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__6_), .B(gnd), .Y(micro_ucr_hash1_a_13__2_) );
XOR2X1 XOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__7_), .B(gnd), .Y(micro_ucr_hash1_a_13__3_) );
XOR2X1 XOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_12__4_), .B(micro_ucr_hash1_b_12__4_), .Y(micro_ucr_hash1_a_13__4_) );
XOR2X1 XOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_12__5_), .B(micro_ucr_hash1_b_12__5_), .Y(micro_ucr_hash1_a_13__5_) );
XOR2X1 XOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_12__6_), .B(micro_ucr_hash1_b_12__6_), .Y(micro_ucr_hash1_a_13__6_) );
XOR2X1 XOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_12__7_), .B(micro_ucr_hash1_b_12__7_), .Y(micro_ucr_hash1_a_13__7_) );
INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_16_), .Y(_1003_) );
XNOR2X1 XNOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__0_), .Y(_1004_) );
XNOR2X1 XNOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .B(_1003_), .Y(micro_ucr_hash1_b_14__4_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .B(_1004_), .Y(_1005_) );
OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__1_), .Y(_1006_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__1_), .Y(_1007_) );
NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_17_), .B(_1007_), .C(_1006_), .Y(_1008_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_17_), .Y(_1009_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__1_), .Y(_1010_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__1_), .Y(_1011_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1010_), .C(_1009_), .Y(_1012_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1012_), .B(_1008_), .Y(_1013_) );
XNOR2X1 XNOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1013_), .B(_1005_), .Y(micro_ucr_hash1_b_14__5_) );
NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1008_), .B(_1012_), .C(_1005_), .Y(_1014_) );
NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_1009_), .B(_1010_), .C(_1011_), .Y(_1015_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_18_), .Y(_1016_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__2_), .Y(_1017_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__2_), .Y(_1018_) );
NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_1016_), .B(_1017_), .C(_1018_), .Y(_1019_) );
OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__2_), .Y(_1020_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__2_), .Y(_1021_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1021_), .B(_1020_), .C(entrada_hash1_nonce_18_), .Y(_1022_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1022_), .C(_1015_), .Y(_1023_) );
NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_18_), .B(_1021_), .C(_1020_), .Y(_1024_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .B(_1017_), .C(_1016_), .Y(_1025_) );
NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1025_), .B(_1008_), .C(_1024_), .Y(_1026_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1026_), .B(_1023_), .Y(_1027_) );
XNOR2X1 XNOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1027_), .B(_1014_), .Y(micro_ucr_hash1_b_14__6_) );
NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1024_), .B(_1025_), .C(_1015_), .Y(_1028_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1022_), .C(_1008_), .Y(_1029_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1028_), .B(_1029_), .Y(_1030_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_1014_), .C(_1028_), .Y(_1031_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_19_), .Y(_1032_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__3_), .Y(_1033_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__3_), .Y(_1034_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1034_), .B(_1033_), .C(_1032_), .Y(_1035_) );
OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__3_), .Y(_1036_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_12__3_), .Y(_1037_) );
NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_19_), .B(_1037_), .C(_1036_), .Y(_1038_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1038_), .C(_1024_), .Y(_1039_) );
NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1032_), .B(_1037_), .C(_1036_), .Y(_1040_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1034_), .B(_1033_), .C(entrada_hash1_nonce_19_), .Y(_1041_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .B(_1040_), .C(_1019_), .Y(_1042_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1039_), .B(_1042_), .Y(_1002_) );
XOR2X1 XOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1031_), .B(_1002_), .Y(micro_ucr_hash1_b_14__7_) );
XOR2X1 XOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_14__4_), .B(gnd), .Y(micro_ucr_hash1_a_14__0_) );
XOR2X1 XOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_14__5_), .B(gnd), .Y(micro_ucr_hash1_a_14__1_) );
XOR2X1 XOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_14__6_), .B(gnd), .Y(micro_ucr_hash1_a_14__2_) );
XOR2X1 XOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_14__7_), .B(gnd), .Y(micro_ucr_hash1_a_14__3_) );
INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_8_), .Y(_1112_) );
XNOR2X1 XNOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__0_), .Y(_1113_) );
XNOR2X1 XNOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1113_), .B(_1112_), .Y(micro_ucr_hash1_b_15__4_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .B(_1113_), .Y(_1114_) );
OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__1_), .Y(_1115_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__1_), .Y(_1116_) );
NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_9_), .B(_1116_), .C(_1115_), .Y(_1117_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_9_), .Y(_1118_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__1_), .Y(_1119_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__1_), .Y(_1120_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1120_), .B(_1119_), .C(_1118_), .Y(_1121_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1117_), .Y(_1122_) );
XNOR2X1 XNOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_1114_), .Y(micro_ucr_hash1_b_15__5_) );
NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1117_), .B(_1121_), .C(_1114_), .Y(_1123_) );
NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_1118_), .B(_1119_), .C(_1120_), .Y(_1124_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_10_), .Y(_1125_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__2_), .Y(_1126_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__2_), .Y(_1127_) );
NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_1125_), .B(_1126_), .C(_1127_), .Y(_1128_) );
OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__2_), .Y(_1129_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__2_), .Y(_1130_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1130_), .B(_1129_), .C(entrada_hash1_nonce_10_), .Y(_1131_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_1131_), .C(_1124_), .Y(_1132_) );
NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_10_), .B(_1130_), .C(_1129_), .Y(_1133_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1127_), .B(_1126_), .C(_1125_), .Y(_1134_) );
NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1134_), .B(_1117_), .C(_1133_), .Y(_1135_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_1132_), .Y(_1136_) );
XNOR2X1 XNOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1136_), .B(_1123_), .Y(micro_ucr_hash1_b_15__6_) );
NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1133_), .B(_1134_), .C(_1124_), .Y(_1137_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_1131_), .C(_1117_), .Y(_1138_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1138_), .Y(_1139_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1139_), .B(_1123_), .C(_1137_), .Y(_1140_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_11_), .Y(_1141_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__3_), .Y(_1142_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__3_), .Y(_1143_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(_1142_), .C(_1141_), .Y(_1144_) );
OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__3_), .Y(_1145_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_13__3_), .Y(_1146_) );
NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_11_), .B(_1146_), .C(_1145_), .Y(_1147_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_1147_), .C(_1133_), .Y(_1148_) );
NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1146_), .C(_1145_), .Y(_1149_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1143_), .B(_1142_), .C(entrada_hash1_nonce_11_), .Y(_1150_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1150_), .B(_1149_), .C(_1128_), .Y(_1151_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1148_), .B(_1151_), .Y(_1043_) );
XOR2X1 XOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1043_), .Y(micro_ucr_hash1_b_15__7_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_12_), .Y(_1044_) );
OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__4_), .B(micro_ucr_hash1_a_13__4_), .Y(_1045_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__4_), .B(micro_ucr_hash1_a_13__4_), .Y(_1046_) );
NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1044_), .B(_1046_), .C(_1045_), .Y(_1047_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__4_), .B(micro_ucr_hash1_a_13__4_), .Y(_1048_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__4_), .B(micro_ucr_hash1_a_13__4_), .Y(_1049_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1048_), .C(entrada_hash1_nonce_12_), .Y(_1050_) );
NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_1047_), .C(_1050_), .Y(_1051_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1146_), .B(_1145_), .C(entrada_hash1_nonce_11_), .Y(_1052_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1049_), .B(_1048_), .C(_1044_), .Y(_1053_) );
NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_12_), .B(_1046_), .C(_1045_), .Y(_1054_) );
NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .B(_1054_), .C(_1052_), .Y(_1055_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1051_), .Y(_1056_) );
INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .Y(_1057_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1131_), .B(_1128_), .Y(_1058_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1124_), .B(_1058_), .C(_1148_), .Y(_1059_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1139_), .B(_1123_), .C(_1059_), .Y(_1060_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1060_), .Y(_1061_) );
XNOR2X1 XNOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_1056_), .Y(micro_ucr_hash1_c_14__4_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_1055_), .Y(_1062_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_1062_), .C(_1051_), .Y(_1063_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_13_), .Y(_1064_) );
OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__5_), .B(micro_ucr_hash1_a_13__5_), .Y(_1065_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__5_), .B(micro_ucr_hash1_a_13__5_), .Y(_1066_) );
NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1064_), .B(_1066_), .C(_1065_), .Y(_1067_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__5_), .B(micro_ucr_hash1_a_13__5_), .Y(_1068_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__5_), .B(micro_ucr_hash1_a_13__5_), .Y(_1069_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1068_), .C(entrada_hash1_nonce_13_), .Y(_1070_) );
NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1053_), .B(_1070_), .C(_1067_), .Y(_1071_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1046_), .B(_1045_), .C(entrada_hash1_nonce_12_), .Y(_1072_) );
NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_13_), .B(_1066_), .C(_1065_), .Y(_1073_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1069_), .B(_1068_), .C(_1064_), .Y(_1074_) );
NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .B(_1073_), .C(_1072_), .Y(_1075_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .B(_1075_), .Y(_1076_) );
INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .Y(_1077_) );
XNOR2X1 XNOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1077_), .Y(micro_ucr_hash1_c_14__5_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1071_), .B(_1075_), .C(_1062_), .Y(_1078_) );
NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1078_), .C(_1060_), .Y(_1079_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1074_), .B(_1073_), .Y(_1080_) );
OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(_1072_), .Y(_1081_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .Y(_1082_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1080_), .C(_1051_), .Y(_1083_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1082_), .Y(_1084_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_14_), .Y(_1085_) );
XNOR2X1 XNOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__6_), .B(micro_ucr_hash1_a_13__6_), .Y(_1086_) );
OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_1086_), .B(_1085_), .Y(_1087_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1085_), .B(_1086_), .Y(_1088_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1088_), .B(_1087_), .Y(_1089_) );
OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1073_), .Y(_1090_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_1089_), .Y(_1091_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1091_), .B(_1090_), .Y(_1092_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1079_), .C(_1092_), .Y(_1093_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .B(_1056_), .Y(_1094_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1061_), .B(_1094_), .C(_1084_), .Y(_1095_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_1092_), .Y(_1096_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1095_), .Y(_1097_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(_1097_), .Y(micro_ucr_hash1_c_14__6_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .Y(_1098_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1057_), .B(_1098_), .C(_1148_), .Y(_1099_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .B(_1113_), .C(_1122_), .Y(_1100_) );
NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1100_), .B(_1136_), .C(_1043_), .Y(_1101_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1099_), .B(_1101_), .C(_1094_), .Y(_1102_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1077_), .B(_1051_), .C(_1081_), .Y(_1103_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1102_), .B(_1103_), .C(_1096_), .Y(_1104_) );
XOR2X1 XOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__7_), .B(entrada_hash1_nonce_15_), .Y(_1105_) );
XNOR2X1 XNOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1105_), .B(micro_ucr_hash1_a_13__7_), .Y(_1106_) );
XNOR2X1 XNOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1106_), .B(_1087_), .Y(_1107_) );
NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1107_), .C(_1104_), .Y(_1108_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .Y(_1109_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_1107_), .Y(_1110_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(_1109_), .C(_1110_), .Y(_1111_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1108_), .B(_1111_), .Y(micro_ucr_hash1_c_14__7_) );
XOR2X1 XOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__4_), .B(gnd), .Y(micro_ucr_hash1_a_15__0_) );
XOR2X1 XOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__5_), .B(gnd), .Y(micro_ucr_hash1_a_15__1_) );
XOR2X1 XOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__6_), .B(gnd), .Y(micro_ucr_hash1_a_15__2_) );
XOR2X1 XOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__7_), .B(gnd), .Y(micro_ucr_hash1_a_15__3_) );
XOR2X1 XOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_14__4_), .B(micro_ucr_hash1_b_14__4_), .Y(micro_ucr_hash1_a_15__4_) );
XOR2X1 XOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_14__5_), .B(micro_ucr_hash1_b_14__5_), .Y(micro_ucr_hash1_a_15__5_) );
XOR2X1 XOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_14__6_), .B(micro_ucr_hash1_b_14__6_), .Y(micro_ucr_hash1_a_15__6_) );
XOR2X1 XOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_14__7_), .B(micro_ucr_hash1_b_14__7_), .Y(micro_ucr_hash1_a_15__7_) );
INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_0_), .Y(_1153_) );
XNOR2X1 XNOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__0_), .Y(_1154_) );
XNOR2X1 XNOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1154_), .B(_1153_), .Y(micro_ucr_hash1_b_16__4_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1154_), .Y(_1155_) );
OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__1_), .Y(_1156_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__1_), .Y(_1157_) );
NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_1_), .B(_1157_), .C(_1156_), .Y(_1158_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_1_), .Y(_1159_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__1_), .Y(_1160_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__1_), .Y(_1161_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_1161_), .B(_1160_), .C(_1159_), .Y(_1162_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1162_), .B(_1158_), .Y(_1163_) );
XNOR2X1 XNOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1163_), .B(_1155_), .Y(micro_ucr_hash1_b_16__5_) );
NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1158_), .B(_1162_), .C(_1155_), .Y(_1164_) );
NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_1160_), .C(_1161_), .Y(_1165_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_2_), .Y(_1166_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__2_), .Y(_1167_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__2_), .Y(_1168_) );
NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_1166_), .B(_1167_), .C(_1168_), .Y(_1169_) );
OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__2_), .Y(_1170_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__2_), .Y(_1171_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1171_), .B(_1170_), .C(entrada_hash1_nonce_2_), .Y(_1172_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1172_), .C(_1165_), .Y(_1173_) );
NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_2_), .B(_1171_), .C(_1170_), .Y(_1174_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1168_), .B(_1167_), .C(_1166_), .Y(_1175_) );
NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(_1158_), .C(_1174_), .Y(_1176_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1176_), .B(_1173_), .Y(_1177_) );
XNOR2X1 XNOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_1164_), .Y(micro_ucr_hash1_b_16__6_) );
NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1174_), .B(_1175_), .C(_1165_), .Y(_1178_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1172_), .C(_1158_), .Y(_1179_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1178_), .B(_1179_), .Y(_1180_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1180_), .B(_1164_), .C(_1178_), .Y(_1181_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_3_), .Y(_1182_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__3_), .Y(_1183_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__3_), .Y(_1184_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(_1183_), .C(_1182_), .Y(_1185_) );
OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__3_), .Y(_1186_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_14__3_), .Y(_1187_) );
NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_3_), .B(_1187_), .C(_1186_), .Y(_1188_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(_1188_), .C(_1174_), .Y(_1189_) );
NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1182_), .B(_1187_), .C(_1186_), .Y(_1190_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(_1183_), .C(entrada_hash1_nonce_3_), .Y(_1191_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1191_), .B(_1190_), .C(_1169_), .Y(_1192_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1189_), .B(_1192_), .Y(_1152_) );
XOR2X1 XOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(_1152_), .Y(micro_ucr_hash1_b_16__7_) );
XOR2X1 XOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_16__4_), .B(gnd), .Y(micro_ucr_hash1_a_16__0_) );
XOR2X1 XOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_16__5_), .B(gnd), .Y(micro_ucr_hash1_a_16__1_) );
XOR2X1 XOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_16__6_), .B(gnd), .Y(micro_ucr_hash1_a_16__2_) );
XOR2X1 XOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_16__7_), .B(gnd), .Y(micro_ucr_hash1_a_16__3_) );
INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__0_), .Y(_1262_) );
XNOR2X1 XNOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__0_), .Y(_1263_) );
XNOR2X1 XNOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1263_), .B(_1262_), .Y(micro_ucr_hash1_b_17__4_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .B(_1263_), .Y(_1264_) );
OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__1_), .Y(_1265_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__1_), .Y(_1266_) );
NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__1_), .B(_1266_), .C(_1265_), .Y(_1267_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__1_), .Y(_1268_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__1_), .Y(_1269_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__1_), .Y(_1270_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1270_), .B(_1269_), .C(_1268_), .Y(_1271_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1271_), .B(_1267_), .Y(_1272_) );
XNOR2X1 XNOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1272_), .B(_1264_), .Y(micro_ucr_hash1_b_17__5_) );
NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1271_), .C(_1264_), .Y(_1273_) );
NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_1269_), .C(_1270_), .Y(_1274_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__2_), .Y(_1275_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__2_), .Y(_1276_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__2_), .Y(_1277_) );
NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_1275_), .B(_1276_), .C(_1277_), .Y(_1278_) );
OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__2_), .Y(_1279_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__2_), .Y(_1280_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1279_), .C(micro_ucr_hash1_W_16__2_), .Y(_1281_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .B(_1281_), .C(_1274_), .Y(_1282_) );
NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__2_), .B(_1280_), .C(_1279_), .Y(_1283_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1277_), .B(_1276_), .C(_1275_), .Y(_1284_) );
NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .B(_1267_), .C(_1283_), .Y(_1285_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1285_), .B(_1282_), .Y(_1286_) );
XNOR2X1 XNOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1273_), .Y(micro_ucr_hash1_b_17__6_) );
NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(_1284_), .C(_1274_), .Y(_1287_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .B(_1281_), .C(_1267_), .Y(_1288_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1287_), .B(_1288_), .Y(_1289_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1273_), .C(_1287_), .Y(_1290_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__3_), .Y(_1291_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__3_), .Y(_1292_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__3_), .Y(_1293_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1293_), .B(_1292_), .C(_1291_), .Y(_1294_) );
OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__3_), .Y(_1295_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_15__3_), .Y(_1296_) );
NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__3_), .B(_1296_), .C(_1295_), .Y(_1297_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_1297_), .C(_1283_), .Y(_1298_) );
NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1291_), .B(_1296_), .C(_1295_), .Y(_1299_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1293_), .B(_1292_), .C(micro_ucr_hash1_W_16__3_), .Y(_1300_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1300_), .B(_1299_), .C(_1278_), .Y(_1301_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1298_), .B(_1301_), .Y(_1193_) );
XOR2X1 XOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1290_), .B(_1193_), .Y(micro_ucr_hash1_b_17__7_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__4_), .Y(_1194_) );
OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__4_), .B(micro_ucr_hash1_a_15__4_), .Y(_1195_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__4_), .B(micro_ucr_hash1_a_15__4_), .Y(_1196_) );
NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1194_), .B(_1196_), .C(_1195_), .Y(_1197_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__4_), .B(micro_ucr_hash1_a_15__4_), .Y(_1198_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__4_), .B(micro_ucr_hash1_a_15__4_), .Y(_1199_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .B(_1198_), .C(micro_ucr_hash1_W_16__4_), .Y(_1200_) );
NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_1197_), .C(_1200_), .Y(_1201_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1296_), .B(_1295_), .C(micro_ucr_hash1_W_16__3_), .Y(_1202_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1199_), .B(_1198_), .C(_1194_), .Y(_1203_) );
NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__4_), .B(_1196_), .C(_1195_), .Y(_1204_) );
NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(_1204_), .C(_1202_), .Y(_1205_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1201_), .Y(_1206_) );
INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(_1301_), .Y(_1207_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1281_), .B(_1278_), .Y(_1208_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1274_), .B(_1208_), .C(_1298_), .Y(_1209_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1273_), .C(_1209_), .Y(_1210_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1210_), .Y(_1211_) );
XNOR2X1 XNOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1211_), .B(_1206_), .Y(micro_ucr_hash1_c_16__4_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(_1205_), .Y(_1212_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1211_), .B(_1212_), .C(_1201_), .Y(_1213_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__5_), .Y(_1214_) );
OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__5_), .B(micro_ucr_hash1_a_15__5_), .Y(_1215_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__5_), .B(micro_ucr_hash1_a_15__5_), .Y(_1216_) );
NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1214_), .B(_1216_), .C(_1215_), .Y(_1217_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__5_), .B(micro_ucr_hash1_a_15__5_), .Y(_1218_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__5_), .B(micro_ucr_hash1_a_15__5_), .Y(_1219_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1219_), .B(_1218_), .C(micro_ucr_hash1_W_16__5_), .Y(_1220_) );
NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(_1220_), .C(_1217_), .Y(_1221_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1196_), .B(_1195_), .C(micro_ucr_hash1_W_16__4_), .Y(_1222_) );
NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__5_), .B(_1216_), .C(_1215_), .Y(_1223_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1219_), .B(_1218_), .C(_1214_), .Y(_1224_) );
NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .B(_1223_), .C(_1222_), .Y(_1225_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .B(_1225_), .Y(_1226_) );
INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .Y(_1227_) );
XNOR2X1 XNOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1213_), .B(_1227_), .Y(micro_ucr_hash1_c_16__5_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .B(_1225_), .C(_1212_), .Y(_1228_) );
NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1228_), .C(_1210_), .Y(_1229_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .B(_1223_), .Y(_1230_) );
OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_1230_), .B(_1222_), .Y(_1231_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(_1231_), .Y(_1232_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .B(_1230_), .C(_1201_), .Y(_1233_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1233_), .B(_1232_), .Y(_1234_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__6_), .Y(_1235_) );
XNOR2X1 XNOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__6_), .B(micro_ucr_hash1_a_15__6_), .Y(_1236_) );
OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_1235_), .Y(_1237_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1235_), .B(_1236_), .Y(_1238_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1238_), .B(_1237_), .Y(_1239_) );
OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_1239_), .B(_1223_), .Y(_1240_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1239_), .Y(_1241_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_1240_), .Y(_1242_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1234_), .B(_1229_), .C(_1242_), .Y(_1243_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1226_), .B(_1206_), .Y(_1244_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1211_), .B(_1244_), .C(_1234_), .Y(_1245_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(_1242_), .Y(_1246_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1246_), .B(_1245_), .Y(_1247_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1243_), .B(_1247_), .Y(micro_ucr_hash1_c_16__6_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(_1287_), .Y(_1248_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1207_), .B(_1248_), .C(_1298_), .Y(_1249_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .B(_1263_), .C(_1272_), .Y(_1250_) );
NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1250_), .B(_1286_), .C(_1193_), .Y(_1251_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1249_), .B(_1251_), .C(_1244_), .Y(_1252_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1227_), .B(_1201_), .C(_1231_), .Y(_1253_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1252_), .B(_1253_), .C(_1246_), .Y(_1254_) );
XOR2X1 XOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__7_), .B(micro_ucr_hash1_W_16__7_), .Y(_1255_) );
XNOR2X1 XNOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1255_), .B(micro_ucr_hash1_a_15__7_), .Y(_1256_) );
XNOR2X1 XNOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1256_), .B(_1237_), .Y(_1257_) );
NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .B(_1257_), .C(_1254_), .Y(_1258_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .Y(_1259_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(_1257_), .Y(_1260_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1243_), .B(_1259_), .C(_1260_), .Y(_1261_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1258_), .B(_1261_), .Y(micro_ucr_hash1_c_16__7_) );
XOR2X1 XOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__4_), .B(gnd), .Y(micro_ucr_hash1_a_17__0_) );
XOR2X1 XOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__5_), .B(gnd), .Y(micro_ucr_hash1_a_17__1_) );
XOR2X1 XOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__6_), .B(gnd), .Y(micro_ucr_hash1_a_17__2_) );
XOR2X1 XOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__7_), .B(gnd), .Y(micro_ucr_hash1_a_17__3_) );
XOR2X1 XOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_16__4_), .B(micro_ucr_hash1_b_16__4_), .Y(micro_ucr_hash1_a_17__4_) );
XOR2X1 XOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_16__5_), .B(micro_ucr_hash1_b_16__5_), .Y(micro_ucr_hash1_a_17__5_) );
XOR2X1 XOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_16__6_), .B(micro_ucr_hash1_b_16__6_), .Y(micro_ucr_hash1_a_17__6_) );
XOR2X1 XOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_16__7_), .B(micro_ucr_hash1_b_16__7_), .Y(micro_ucr_hash1_a_17__7_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_17__0_), .Y(_1302_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_16__0_), .Y(_1303_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(_1303_), .Y(_1304_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_16__0_), .C(micro_ucr_hash1_W_17__0_), .Y(_1305_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1305_), .B(_1304_), .Y(micro_ucr_hash1_b_18__4_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_16__1_), .C(micro_ucr_hash1_W_17__1_), .Y(_1306_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_17__1_), .Y(_1307_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_16__1_), .Y(_1308_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(_1308_), .Y(_1309_) );
NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .B(_1304_), .C(_1309_), .Y(_1310_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .B(_1302_), .Y(_1311_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_1306_), .Y(_1312_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(_1307_), .Y(_1313_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1313_), .B(_1312_), .C(_1311_), .Y(_1314_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_1310_), .Y(micro_ucr_hash1_b_18__5_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_16__2_), .C(micro_ucr_hash1_W_17__2_), .Y(_1315_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_17__2_), .Y(_1316_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_16__2_), .Y(_1317_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(_1317_), .Y(_1318_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1315_), .B(_1318_), .Y(_1319_) );
NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1315_), .B(_1318_), .C(_1312_), .Y(_1320_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .B(_1319_), .C(_1320_), .Y(_1321_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_1319_), .Y(_1322_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1311_), .B(_1313_), .C(_1306_), .Y(_1323_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1323_), .B(_1322_), .Y(_1324_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_1324_), .Y(micro_ucr_hash1_b_18__6_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_17__3_), .Y(_1325_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_16__3_), .C(_1325_), .Y(_1326_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_16__3_), .Y(_1327_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_17__3_), .B(_1327_), .Y(_1328_) );
NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1315_), .B(_1326_), .C(_1328_), .Y(_1329_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(_1315_), .Y(_1330_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_16__3_), .C(micro_ucr_hash1_W_17__3_), .Y(_1331_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_1327_), .Y(_1332_) );
NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1331_), .B(_1332_), .C(_1330_), .Y(_1333_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1329_), .B(_1333_), .Y(_1334_) );
XNOR2X1 XNOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_1334_), .Y(micro_ucr_hash1_b_18__7_) );
XOR2X1 XOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_18__4_), .B(gnd), .Y(micro_ucr_hash1_a_18__0_) );
XOR2X1 XOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_18__5_), .B(gnd), .Y(micro_ucr_hash1_a_18__1_) );
XOR2X1 XOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_18__6_), .B(gnd), .Y(micro_ucr_hash1_a_18__2_) );
XOR2X1 XOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_18__7_), .B(gnd), .Y(micro_ucr_hash1_a_18__3_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__0_), .Y(_1391_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__0_), .Y(_1392_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_1392_), .Y(_1393_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__0_), .C(micro_ucr_hash1_W_18__0_), .Y(_1394_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1394_), .B(_1393_), .Y(micro_ucr_hash1_b_19__4_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__1_), .C(micro_ucr_hash1_W_18__1_), .Y(_1395_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__1_), .Y(_1396_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__1_), .Y(_1397_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1396_), .B(_1397_), .Y(_1398_) );
NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_1393_), .C(_1398_), .Y(_1399_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_1392_), .B(_1391_), .Y(_1400_) );
INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .Y(_1401_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_1397_), .B(_1396_), .Y(_1402_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .B(_1401_), .C(_1400_), .Y(_1403_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_1403_), .B(_1399_), .Y(micro_ucr_hash1_b_19__5_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__2_), .C(micro_ucr_hash1_W_18__2_), .Y(_1404_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__2_), .Y(_1405_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__2_), .Y(_1406_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1405_), .B(_1406_), .Y(_1407_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1404_), .B(_1407_), .Y(_1408_) );
NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1404_), .B(_1407_), .C(_1401_), .Y(_1409_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1399_), .B(_1408_), .C(_1409_), .Y(_1410_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .Y(_1411_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1400_), .B(_1402_), .C(_1395_), .Y(_1412_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .B(_1411_), .Y(_1413_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1410_), .B(_1413_), .Y(micro_ucr_hash1_b_19__6_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__3_), .Y(_1414_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__3_), .C(_1414_), .Y(_1415_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__3_), .Y(_1416_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__3_), .B(_1416_), .Y(_1417_) );
NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1404_), .B(_1415_), .C(_1417_), .Y(_1418_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(_1404_), .Y(_1419_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__3_), .C(micro_ucr_hash1_W_18__3_), .Y(_1420_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_1416_), .Y(_1421_) );
NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1421_), .C(_1419_), .Y(_1422_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(_1422_), .Y(_1423_) );
XNOR2X1 XNOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1410_), .B(_1423_), .Y(micro_ucr_hash1_b_19__7_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .Y(_1424_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__4_), .B(micro_ucr_hash1_a_17__4_), .C(micro_ucr_hash1_W_18__4_), .Y(_1425_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__4_), .Y(_1426_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_17__4_), .Y(_1427_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__4_), .Y(_1428_) );
NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1426_), .B(_1427_), .C(_1428_), .Y(_1429_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1425_), .B(_1429_), .C(_1424_), .Y(_1335_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__4_), .B(micro_ucr_hash1_a_17__4_), .C(_1428_), .Y(_1336_) );
NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__4_), .B(_1426_), .C(_1427_), .Y(_1337_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1337_), .C(_1420_), .Y(_1338_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1338_), .B(_1335_), .Y(_1339_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1421_), .C(_1419_), .Y(_1340_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_1409_), .C(_1422_), .Y(_1341_) );
NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_1399_), .B(_1408_), .C(_1340_), .Y(_1342_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_1342_), .Y(_1343_) );
XNOR2X1 XNOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1339_), .Y(micro_ucr_hash1_c_18__4_) );
NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1425_), .B(_1429_), .C(_1424_), .Y(_1344_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1335_), .C(_1344_), .Y(_1345_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__5_), .Y(_1346_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__5_), .B(micro_ucr_hash1_a_17__5_), .C(_1346_), .Y(_1347_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__5_), .B(micro_ucr_hash1_a_17__5_), .Y(_1348_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__5_), .B(_1348_), .Y(_1349_) );
NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1425_), .B(_1347_), .C(_1349_), .Y(_1350_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(_1425_), .Y(_1351_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(_1348_), .Y(_1352_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__5_), .B(micro_ucr_hash1_a_17__5_), .C(micro_ucr_hash1_W_18__5_), .Y(_1353_) );
NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1353_), .B(_1352_), .C(_1351_), .Y(_1354_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_1354_), .Y(_1355_) );
XOR2X1 XOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_1355_), .Y(micro_ucr_hash1_c_18__5_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_17__2_), .C(_1405_), .Y(_1356_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__2_), .B(_1406_), .Y(_1357_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1356_), .B(_1357_), .C(_1395_), .Y(_1358_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .Y(_1359_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(_1358_), .C(_1359_), .Y(_1360_) );
NOR3X1 NOR3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_1400_), .B(_1401_), .C(_1402_), .Y(_1361_) );
NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1411_), .B(_1418_), .C(_1361_), .Y(_1362_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1355_), .B(_1339_), .Y(_1363_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1360_), .B(_1362_), .C(_1363_), .Y(_1364_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .B(_1353_), .C(_1344_), .D(_1425_), .Y(_1365_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(_1352_), .Y(_1366_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__6_), .B(micro_ucr_hash1_a_17__6_), .C(micro_ucr_hash1_W_18__6_), .Y(_1367_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_18__6_), .Y(_1368_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__6_), .B(micro_ucr_hash1_a_17__6_), .Y(_1369_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1368_), .B(_1369_), .Y(_1370_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .B(_1370_), .Y(_1371_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(_1371_), .Y(_1372_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .Y(_1373_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(_1371_), .Y(_1374_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1374_), .B(_1373_), .Y(_1375_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(_1375_), .Y(_1376_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1364_), .B(_1365_), .C(_1376_), .Y(_1377_) );
NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1336_), .C(_1337_), .Y(_1378_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1378_), .B(_1344_), .Y(_1379_) );
AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1350_), .B(_1354_), .C(_1379_), .Y(_1380_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_1342_), .C(_1380_), .Y(_1381_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(_1365_), .Y(_1382_) );
NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1382_), .B(_1375_), .C(_1381_), .Y(_1383_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .B(_1383_), .Y(micro_ucr_hash1_c_18__6_) );
AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1382_), .B(_1381_), .C(_1375_), .Y(_1384_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__7_), .B(micro_ucr_hash1_a_17__7_), .Y(_1385_) );
XNOR2X1 XNOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1385_), .B(micro_ucr_hash1_W_18__7_), .Y(_1386_) );
XNOR2X1 XNOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1386_), .B(_1367_), .Y(_1387_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1384_), .B(_1372_), .C(_1387_), .Y(_1388_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(_1387_), .Y(_1389_) );
NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1373_), .B(_1389_), .C(_1377_), .Y(_1390_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1388_), .B(_1390_), .Y(micro_ucr_hash1_c_18__7_) );
XOR2X1 XOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__4_), .B(gnd), .Y(micro_ucr_hash1_a_19__0_) );
XOR2X1 XOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__5_), .B(gnd), .Y(micro_ucr_hash1_a_19__1_) );
XOR2X1 XOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__6_), .B(gnd), .Y(micro_ucr_hash1_a_19__2_) );
XOR2X1 XOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__7_), .B(gnd), .Y(micro_ucr_hash1_a_19__3_) );
XOR2X1 XOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_18__4_), .B(micro_ucr_hash1_b_18__4_), .Y(micro_ucr_hash1_a_19__4_) );
XOR2X1 XOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_18__5_), .B(micro_ucr_hash1_b_18__5_), .Y(micro_ucr_hash1_a_19__5_) );
XOR2X1 XOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_18__6_), .B(micro_ucr_hash1_b_18__6_), .Y(micro_ucr_hash1_a_19__6_) );
XOR2X1 XOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_18__7_), .B(micro_ucr_hash1_b_18__7_), .Y(micro_ucr_hash1_a_19__7_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_19__0_), .Y(_1430_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_18__0_), .Y(_1431_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1430_), .B(_1431_), .Y(_1432_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_18__0_), .C(micro_ucr_hash1_W_19__0_), .Y(_1433_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1433_), .B(_1432_), .Y(micro_ucr_hash1_b_20__4_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_18__1_), .C(micro_ucr_hash1_W_19__1_), .Y(_1434_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_19__1_), .Y(_1435_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_18__1_), .Y(_1436_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1435_), .B(_1436_), .Y(_1437_) );
NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1432_), .C(_1437_), .Y(_1438_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_1431_), .B(_1430_), .Y(_1439_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .Y(_1440_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_1435_), .Y(_1441_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1441_), .B(_1440_), .C(_1439_), .Y(_1442_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_1442_), .B(_1438_), .Y(micro_ucr_hash1_b_20__5_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_18__2_), .C(micro_ucr_hash1_W_19__2_), .Y(_1443_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_19__2_), .Y(_1444_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_18__2_), .Y(_1445_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1444_), .B(_1445_), .Y(_1446_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .B(_1446_), .Y(_1447_) );
NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .B(_1446_), .C(_1440_), .Y(_1448_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1438_), .B(_1447_), .C(_1448_), .Y(_1449_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .Y(_1450_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(_1441_), .C(_1434_), .Y(_1451_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1451_), .B(_1450_), .Y(_1452_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .B(_1452_), .Y(micro_ucr_hash1_b_20__6_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_19__3_), .Y(_1453_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_18__3_), .C(_1453_), .Y(_1454_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_18__3_), .Y(_1455_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_19__3_), .B(_1455_), .Y(_1456_) );
NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .B(_1454_), .C(_1456_), .Y(_1457_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(_1443_), .Y(_1458_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_18__3_), .C(micro_ucr_hash1_W_19__3_), .Y(_1459_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1455_), .Y(_1460_) );
NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .B(_1460_), .C(_1458_), .Y(_1461_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1457_), .B(_1461_), .Y(_1462_) );
XNOR2X1 XNOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .B(_1462_), .Y(micro_ucr_hash1_b_20__7_) );
XOR2X1 XOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_20__4_), .B(gnd), .Y(micro_ucr_hash1_a_20__0_) );
XOR2X1 XOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_20__5_), .B(gnd), .Y(micro_ucr_hash1_a_20__1_) );
XOR2X1 XOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_20__6_), .B(gnd), .Y(micro_ucr_hash1_a_20__2_) );
XOR2X1 XOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_20__7_), .B(gnd), .Y(micro_ucr_hash1_a_20__3_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__0_), .Y(_1519_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__0_), .Y(_1520_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1519_), .B(_1520_), .Y(_1521_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__0_), .C(micro_ucr_hash1_W_20__0_), .Y(_1522_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1522_), .B(_1521_), .Y(micro_ucr_hash1_b_21__4_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__1_), .C(micro_ucr_hash1_W_20__1_), .Y(_1523_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__1_), .Y(_1524_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__1_), .Y(_1525_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1525_), .Y(_1526_) );
NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .B(_1521_), .C(_1526_), .Y(_1527_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(_1520_), .B(_1519_), .Y(_1528_) );
INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .Y(_1529_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_1525_), .B(_1524_), .Y(_1530_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1530_), .B(_1529_), .C(_1528_), .Y(_1531_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_1531_), .B(_1527_), .Y(micro_ucr_hash1_b_21__5_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__2_), .C(micro_ucr_hash1_W_20__2_), .Y(_1532_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__2_), .Y(_1533_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__2_), .Y(_1534_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1533_), .B(_1534_), .Y(_1535_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_1535_), .Y(_1536_) );
NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_1535_), .C(_1529_), .Y(_1537_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1536_), .C(_1537_), .Y(_1538_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(_1536_), .Y(_1539_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1530_), .C(_1523_), .Y(_1540_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1540_), .B(_1539_), .Y(_1541_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1541_), .Y(micro_ucr_hash1_b_21__6_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__3_), .Y(_1542_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__3_), .C(_1542_), .Y(_1543_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__3_), .Y(_1544_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__3_), .B(_1544_), .Y(_1545_) );
NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .B(_1543_), .C(_1545_), .Y(_1546_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(_1532_), .Y(_1547_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__3_), .C(micro_ucr_hash1_W_20__3_), .Y(_1548_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .B(_1544_), .Y(_1549_) );
NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_1549_), .C(_1547_), .Y(_1550_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1546_), .B(_1550_), .Y(_1551_) );
XNOR2X1 XNOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1551_), .Y(micro_ucr_hash1_b_21__7_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .Y(_1552_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__4_), .B(micro_ucr_hash1_a_19__4_), .C(micro_ucr_hash1_W_20__4_), .Y(_1553_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__4_), .Y(_1554_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_19__4_), .Y(_1555_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__4_), .Y(_1556_) );
NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1554_), .B(_1555_), .C(_1556_), .Y(_1557_) );
AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1557_), .C(_1552_), .Y(_1463_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__4_), .B(micro_ucr_hash1_a_19__4_), .C(_1556_), .Y(_1464_) );
NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__4_), .B(_1554_), .C(_1555_), .Y(_1465_) );
AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1465_), .C(_1548_), .Y(_1466_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1466_), .B(_1463_), .Y(_1467_) );
AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_1549_), .C(_1547_), .Y(_1468_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_1537_), .C(_1550_), .Y(_1469_) );
NOR3X1 NOR3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_1527_), .B(_1536_), .C(_1468_), .Y(_1470_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_1470_), .Y(_1471_) );
XNOR2X1 XNOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_1467_), .Y(micro_ucr_hash1_c_20__4_) );
NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1557_), .C(_1552_), .Y(_1472_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1471_), .B(_1463_), .C(_1472_), .Y(_1473_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__5_), .Y(_1474_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__5_), .B(micro_ucr_hash1_a_19__5_), .C(_1474_), .Y(_1475_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__5_), .B(micro_ucr_hash1_a_19__5_), .Y(_1476_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__5_), .B(_1476_), .Y(_1477_) );
NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1475_), .C(_1477_), .Y(_1478_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .Y(_1479_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1474_), .B(_1476_), .Y(_1480_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__5_), .B(micro_ucr_hash1_a_19__5_), .C(micro_ucr_hash1_W_20__5_), .Y(_1481_) );
NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1481_), .B(_1480_), .C(_1479_), .Y(_1482_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .B(_1482_), .Y(_1483_) );
XOR2X1 XOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(_1483_), .Y(micro_ucr_hash1_c_20__5_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_19__2_), .C(_1533_), .Y(_1484_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__2_), .B(_1534_), .Y(_1485_) );
AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .B(_1485_), .C(_1523_), .Y(_1486_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(_1550_), .Y(_1487_) );
AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1546_), .B(_1486_), .C(_1487_), .Y(_1488_) );
NOR3X1 NOR3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_1528_), .B(_1529_), .C(_1530_), .Y(_1489_) );
NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1539_), .B(_1546_), .C(_1489_), .Y(_1490_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1483_), .B(_1467_), .Y(_1491_) );
AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_1488_), .B(_1490_), .C(_1491_), .Y(_1492_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .B(_1481_), .C(_1472_), .D(_1553_), .Y(_1493_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(_1480_), .Y(_1494_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__6_), .B(micro_ucr_hash1_a_19__6_), .C(micro_ucr_hash1_W_20__6_), .Y(_1495_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_20__6_), .Y(_1496_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__6_), .B(micro_ucr_hash1_a_19__6_), .Y(_1497_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1496_), .B(_1497_), .Y(_1498_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(_1498_), .Y(_1499_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .B(_1499_), .Y(_1500_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .Y(_1501_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .B(_1499_), .Y(_1502_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1502_), .B(_1501_), .Y(_1503_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(_1503_), .Y(_1504_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1492_), .B(_1493_), .C(_1504_), .Y(_1505_) );
NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_1464_), .C(_1465_), .Y(_1506_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1506_), .B(_1472_), .Y(_1507_) );
AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1478_), .B(_1482_), .C(_1507_), .Y(_1508_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1469_), .B(_1470_), .C(_1508_), .Y(_1509_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .Y(_1510_) );
NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1510_), .B(_1503_), .C(_1509_), .Y(_1511_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_1505_), .B(_1511_), .Y(micro_ucr_hash1_c_20__6_) );
AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1510_), .B(_1509_), .C(_1503_), .Y(_1512_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__7_), .B(micro_ucr_hash1_a_19__7_), .Y(_1513_) );
XNOR2X1 XNOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1513_), .B(micro_ucr_hash1_W_20__7_), .Y(_1514_) );
XNOR2X1 XNOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1514_), .B(_1495_), .Y(_1515_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1512_), .B(_1500_), .C(_1515_), .Y(_1516_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(_1515_), .Y(_1517_) );
NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1501_), .B(_1517_), .C(_1505_), .Y(_1518_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1516_), .B(_1518_), .Y(micro_ucr_hash1_c_20__7_) );
XOR2X1 XOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__4_), .B(gnd), .Y(micro_ucr_hash1_a_21__0_) );
XOR2X1 XOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__5_), .B(gnd), .Y(micro_ucr_hash1_a_21__1_) );
XOR2X1 XOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__6_), .B(gnd), .Y(micro_ucr_hash1_a_21__2_) );
XOR2X1 XOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__7_), .B(gnd), .Y(micro_ucr_hash1_a_21__3_) );
XOR2X1 XOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_20__4_), .B(micro_ucr_hash1_b_20__4_), .Y(micro_ucr_hash1_a_21__4_) );
XOR2X1 XOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_20__5_), .B(micro_ucr_hash1_b_20__5_), .Y(micro_ucr_hash1_a_21__5_) );
XOR2X1 XOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_20__6_), .B(micro_ucr_hash1_b_20__6_), .Y(micro_ucr_hash1_a_21__6_) );
XOR2X1 XOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_20__7_), .B(micro_ucr_hash1_b_20__7_), .Y(micro_ucr_hash1_a_21__7_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_21__0_), .Y(_1558_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_20__0_), .Y(_1559_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1558_), .B(_1559_), .Y(_1560_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_20__0_), .C(micro_ucr_hash1_W_21__0_), .Y(_1561_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1561_), .B(_1560_), .Y(micro_ucr_hash1_b_22__4_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_20__1_), .C(micro_ucr_hash1_W_21__1_), .Y(_1562_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_21__1_), .Y(_1563_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_20__1_), .Y(_1564_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1563_), .B(_1564_), .Y(_1565_) );
NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .B(_1560_), .C(_1565_), .Y(_1566_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(_1558_), .Y(_1567_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .Y(_1568_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_1564_), .B(_1563_), .Y(_1569_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(_1568_), .C(_1567_), .Y(_1570_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_1570_), .B(_1566_), .Y(micro_ucr_hash1_b_22__5_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_20__2_), .C(micro_ucr_hash1_W_21__2_), .Y(_1571_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_21__2_), .Y(_1572_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_20__2_), .Y(_1573_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1572_), .B(_1573_), .Y(_1574_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .B(_1574_), .Y(_1575_) );
NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .B(_1574_), .C(_1568_), .Y(_1576_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1566_), .B(_1575_), .C(_1576_), .Y(_1577_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(_1575_), .Y(_1578_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1567_), .B(_1569_), .C(_1562_), .Y(_1579_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1579_), .B(_1578_), .Y(_1580_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .B(_1580_), .Y(micro_ucr_hash1_b_22__6_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_21__3_), .Y(_1581_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_20__3_), .C(_1581_), .Y(_1582_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_20__3_), .Y(_1583_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_21__3_), .B(_1583_), .Y(_1584_) );
NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .B(_1582_), .C(_1584_), .Y(_1585_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(_1571_), .Y(_1586_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_20__3_), .C(micro_ucr_hash1_W_21__3_), .Y(_1587_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1581_), .B(_1583_), .Y(_1588_) );
NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .B(_1588_), .C(_1586_), .Y(_1589_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .B(_1589_), .Y(_1590_) );
XNOR2X1 XNOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1577_), .B(_1590_), .Y(micro_ucr_hash1_b_22__7_) );
XOR2X1 XOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_22__4_), .B(gnd), .Y(micro_ucr_hash1_a_22__0_) );
XOR2X1 XOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_22__5_), .B(gnd), .Y(micro_ucr_hash1_a_22__1_) );
XOR2X1 XOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_22__6_), .B(gnd), .Y(micro_ucr_hash1_a_22__2_) );
XOR2X1 XOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_22__7_), .B(gnd), .Y(micro_ucr_hash1_a_22__3_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__0_), .Y(_1647_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__0_), .Y(_1648_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1647_), .B(_1648_), .Y(_1649_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__0_), .C(micro_ucr_hash1_W_22__0_), .Y(_1650_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1650_), .B(_1649_), .Y(micro_ucr_hash1_b_23__4_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__1_), .C(micro_ucr_hash1_W_22__1_), .Y(_1651_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__1_), .Y(_1652_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__1_), .Y(_1653_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1652_), .B(_1653_), .Y(_1654_) );
NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .B(_1649_), .C(_1654_), .Y(_1655_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_1648_), .B(_1647_), .Y(_1656_) );
INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(_1651_), .Y(_1657_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_1652_), .Y(_1658_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1658_), .B(_1657_), .C(_1656_), .Y(_1659_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_1659_), .B(_1655_), .Y(micro_ucr_hash1_b_23__5_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__2_), .C(micro_ucr_hash1_W_22__2_), .Y(_1660_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__2_), .Y(_1661_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__2_), .Y(_1662_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1661_), .B(_1662_), .Y(_1663_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1663_), .Y(_1664_) );
NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1663_), .C(_1657_), .Y(_1665_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1664_), .C(_1665_), .Y(_1666_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(_1664_), .Y(_1667_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1656_), .B(_1658_), .C(_1651_), .Y(_1668_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1668_), .B(_1667_), .Y(_1669_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1669_), .Y(micro_ucr_hash1_b_23__6_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__3_), .Y(_1670_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__3_), .C(_1670_), .Y(_1671_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__3_), .Y(_1672_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__3_), .B(_1672_), .Y(_1673_) );
NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .B(_1671_), .C(_1673_), .Y(_1674_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(_1660_), .Y(_1675_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__3_), .C(micro_ucr_hash1_W_22__3_), .Y(_1676_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1670_), .B(_1672_), .Y(_1677_) );
NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_1676_), .B(_1677_), .C(_1675_), .Y(_1678_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_1674_), .B(_1678_), .Y(_1679_) );
XNOR2X1 XNOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1666_), .B(_1679_), .Y(micro_ucr_hash1_b_23__7_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(_1676_), .Y(_1680_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__4_), .B(micro_ucr_hash1_a_21__4_), .C(micro_ucr_hash1_W_22__4_), .Y(_1681_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__4_), .Y(_1682_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_21__4_), .Y(_1683_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__4_), .Y(_1684_) );
NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(_1682_), .B(_1683_), .C(_1684_), .Y(_1685_) );
AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .B(_1685_), .C(_1680_), .Y(_1591_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__4_), .B(micro_ucr_hash1_a_21__4_), .C(_1684_), .Y(_1592_) );
NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__4_), .B(_1682_), .C(_1683_), .Y(_1593_) );
AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1592_), .B(_1593_), .C(_1676_), .Y(_1594_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1594_), .B(_1591_), .Y(_1595_) );
AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1676_), .B(_1677_), .C(_1675_), .Y(_1596_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1596_), .B(_1665_), .C(_1678_), .Y(_1597_) );
NOR3X1 NOR3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_1655_), .B(_1664_), .C(_1596_), .Y(_1598_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1597_), .B(_1598_), .Y(_1599_) );
XNOR2X1 XNOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .B(_1595_), .Y(micro_ucr_hash1_c_22__4_) );
NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .B(_1685_), .C(_1680_), .Y(_1600_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1599_), .B(_1591_), .C(_1600_), .Y(_1601_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__5_), .Y(_1602_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__5_), .B(micro_ucr_hash1_a_21__5_), .C(_1602_), .Y(_1603_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__5_), .B(micro_ucr_hash1_a_21__5_), .Y(_1604_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__5_), .B(_1604_), .Y(_1605_) );
NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .B(_1603_), .C(_1605_), .Y(_1606_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(_1681_), .Y(_1607_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .B(_1604_), .Y(_1608_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__5_), .B(micro_ucr_hash1_a_21__5_), .C(micro_ucr_hash1_W_22__5_), .Y(_1609_) );
NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(_1609_), .B(_1608_), .C(_1607_), .Y(_1610_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .B(_1610_), .Y(_1611_) );
XOR2X1 XOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1601_), .B(_1611_), .Y(micro_ucr_hash1_c_22__5_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_21__2_), .C(_1661_), .Y(_1612_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__2_), .B(_1662_), .Y(_1613_) );
AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1612_), .B(_1613_), .C(_1651_), .Y(_1614_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(_1678_), .Y(_1615_) );
AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_1674_), .B(_1614_), .C(_1615_), .Y(_1616_) );
NOR3X1 NOR3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_1656_), .B(_1657_), .C(_1658_), .Y(_1617_) );
NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1667_), .B(_1674_), .C(_1617_), .Y(_1618_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(_1595_), .Y(_1619_) );
AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1616_), .B(_1618_), .C(_1619_), .Y(_1620_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_1609_), .C(_1600_), .D(_1681_), .Y(_1621_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .Y(_1622_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__6_), .B(micro_ucr_hash1_a_21__6_), .C(micro_ucr_hash1_W_22__6_), .Y(_1623_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_22__6_), .Y(_1624_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__6_), .B(micro_ucr_hash1_a_21__6_), .Y(_1625_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_1624_), .B(_1625_), .Y(_1626_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_1623_), .B(_1626_), .Y(_1627_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1622_), .B(_1627_), .Y(_1628_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(_1628_), .Y(_1629_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_1622_), .B(_1627_), .Y(_1630_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_1630_), .B(_1629_), .Y(_1631_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .Y(_1632_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1620_), .B(_1621_), .C(_1632_), .Y(_1633_) );
NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1676_), .B(_1592_), .C(_1593_), .Y(_1634_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1634_), .B(_1600_), .Y(_1635_) );
AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_1606_), .B(_1610_), .C(_1635_), .Y(_1636_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_1597_), .B(_1598_), .C(_1636_), .Y(_1637_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(_1621_), .Y(_1638_) );
NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1638_), .B(_1631_), .C(_1637_), .Y(_1639_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_1633_), .B(_1639_), .Y(micro_ucr_hash1_c_22__6_) );
AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1638_), .B(_1637_), .C(_1631_), .Y(_1640_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__7_), .B(micro_ucr_hash1_a_21__7_), .Y(_1641_) );
XNOR2X1 XNOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1641_), .B(micro_ucr_hash1_W_22__7_), .Y(_1642_) );
XNOR2X1 XNOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1642_), .B(_1623_), .Y(_1643_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1640_), .B(_1628_), .C(_1643_), .Y(_1644_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .Y(_1645_) );
NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_1629_), .B(_1645_), .C(_1633_), .Y(_1646_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1644_), .B(_1646_), .Y(micro_ucr_hash1_c_22__7_) );
XOR2X1 XOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__4_), .B(gnd), .Y(micro_ucr_hash1_a_23__0_) );
XOR2X1 XOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__5_), .B(gnd), .Y(micro_ucr_hash1_a_23__1_) );
XOR2X1 XOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__6_), .B(gnd), .Y(micro_ucr_hash1_a_23__2_) );
XOR2X1 XOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__7_), .B(gnd), .Y(micro_ucr_hash1_a_23__3_) );
XOR2X1 XOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_22__4_), .B(micro_ucr_hash1_b_22__4_), .Y(micro_ucr_hash1_a_23__4_) );
XOR2X1 XOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_22__5_), .B(micro_ucr_hash1_b_22__5_), .Y(micro_ucr_hash1_a_23__5_) );
XOR2X1 XOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_22__6_), .B(micro_ucr_hash1_b_22__6_), .Y(micro_ucr_hash1_a_23__6_) );
XOR2X1 XOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_22__7_), .B(micro_ucr_hash1_b_22__7_), .Y(micro_ucr_hash1_a_23__7_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_23__0_), .Y(_1686_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_22__0_), .Y(_1687_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1686_), .B(_1687_), .Y(_1688_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_22__0_), .C(micro_ucr_hash1_W_23__0_), .Y(_1689_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1689_), .B(_1688_), .Y(micro_ucr_hash1_b_24__4_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_22__1_), .C(micro_ucr_hash1_W_23__1_), .Y(_1690_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_23__1_), .Y(_1691_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_22__1_), .Y(_1692_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_1691_), .B(_1692_), .Y(_1693_) );
NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1690_), .B(_1688_), .C(_1693_), .Y(_1694_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_1687_), .B(_1686_), .Y(_1695_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(_1690_), .Y(_1696_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_1692_), .B(_1691_), .Y(_1697_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1697_), .B(_1696_), .C(_1695_), .Y(_1698_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_1698_), .B(_1694_), .Y(micro_ucr_hash1_b_24__5_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_22__2_), .C(micro_ucr_hash1_W_23__2_), .Y(_1699_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_23__2_), .Y(_1700_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_22__2_), .Y(_1701_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1700_), .B(_1701_), .Y(_1702_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .B(_1702_), .Y(_1703_) );
NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .B(_1702_), .C(_1696_), .Y(_1704_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1694_), .B(_1703_), .C(_1704_), .Y(_1705_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(_1703_), .Y(_1706_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1695_), .B(_1697_), .C(_1690_), .Y(_1707_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1707_), .B(_1706_), .Y(_1708_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .B(_1708_), .Y(micro_ucr_hash1_b_24__6_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_23__3_), .Y(_1709_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_22__3_), .C(_1709_), .Y(_1710_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_22__3_), .Y(_1711_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_23__3_), .B(_1711_), .Y(_1712_) );
NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .B(_1710_), .C(_1712_), .Y(_1713_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(_1699_), .Y(_1714_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_22__3_), .C(micro_ucr_hash1_W_23__3_), .Y(_1715_) );
NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1709_), .B(_1711_), .Y(_1716_) );
NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1715_), .B(_1716_), .C(_1714_), .Y(_1717_) );
NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_1713_), .B(_1717_), .Y(_1718_) );
XNOR2X1 XNOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1705_), .B(_1718_), .Y(micro_ucr_hash1_b_24__7_) );
XOR2X1 XOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_24__4_), .B(gnd), .Y(micro_ucr_hash1_a_24__0_) );
XOR2X1 XOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_24__5_), .B(gnd), .Y(micro_ucr_hash1_a_24__1_) );
XOR2X1 XOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_24__6_), .B(gnd), .Y(micro_ucr_hash1_a_24__2_) );
XOR2X1 XOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_24__7_), .B(gnd), .Y(micro_ucr_hash1_a_24__3_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__0_), .Y(_1775_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__0_), .Y(_1776_) );
NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1775_), .B(_1776_), .Y(_1777_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__0_), .C(micro_ucr_hash1_W_24__0_), .Y(_1778_) );
NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_1778_), .B(_1777_), .Y(micro_ucr_hash1_b_25__4_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__1_), .C(micro_ucr_hash1_W_24__1_), .Y(_1779_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__1_), .Y(_1780_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__1_), .Y(_1781_) );
NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_1780_), .B(_1781_), .Y(_1782_) );
NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1779_), .B(_1777_), .C(_1782_), .Y(_1783_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_1776_), .B(_1775_), .Y(_1784_) );
INVX2 INVX2_48 ( .gnd(gnd), .vdd(vdd), .A(_1779_), .Y(_1785_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_1781_), .B(_1780_), .Y(_1786_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_1786_), .B(_1785_), .C(_1784_), .Y(_1787_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_1787_), .B(_1783_), .Y(micro_ucr_hash1_b_25__5_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__2_), .C(micro_ucr_hash1_W_24__2_), .Y(_1788_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__2_), .Y(_1789_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__2_), .Y(_1790_) );
NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .B(_1790_), .Y(_1791_) );
NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_1788_), .B(_1791_), .Y(_1792_) );
NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_1788_), .B(_1791_), .C(_1785_), .Y(_1793_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_1783_), .B(_1792_), .C(_1793_), .Y(_1794_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .Y(_1795_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1784_), .B(_1786_), .C(_1779_), .Y(_1796_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1796_), .B(_1795_), .Y(_1797_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(_1797_), .Y(micro_ucr_hash1_b_25__6_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__3_), .Y(_1798_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__3_), .C(_1798_), .Y(_1799_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__3_), .Y(_1800_) );
NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__3_), .B(_1800_), .Y(_1801_) );
NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1788_), .B(_1799_), .C(_1801_), .Y(_1802_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(_1788_), .Y(_1803_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__3_), .C(micro_ucr_hash1_W_24__3_), .Y(_1804_) );
NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1798_), .B(_1800_), .Y(_1805_) );
NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1804_), .B(_1805_), .C(_1803_), .Y(_1806_) );
NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .B(_1806_), .Y(_1807_) );
XNOR2X1 XNOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(_1807_), .Y(micro_ucr_hash1_b_25__7_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(_1804_), .Y(_1808_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__4_), .B(micro_ucr_hash1_a_23__4_), .C(micro_ucr_hash1_W_24__4_), .Y(_1809_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__4_), .Y(_1810_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_23__4_), .Y(_1811_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__4_), .Y(_1812_) );
NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(_1810_), .B(_1811_), .C(_1812_), .Y(_1813_) );
AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1809_), .B(_1813_), .C(_1808_), .Y(_1719_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__4_), .B(micro_ucr_hash1_a_23__4_), .C(_1812_), .Y(_1720_) );
NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__4_), .B(_1810_), .C(_1811_), .Y(_1721_) );
AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1720_), .B(_1721_), .C(_1804_), .Y(_1722_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1722_), .B(_1719_), .Y(_1723_) );
AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_1804_), .B(_1805_), .C(_1803_), .Y(_1724_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_1793_), .C(_1806_), .Y(_1725_) );
NOR3X1 NOR3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_1783_), .B(_1792_), .C(_1724_), .Y(_1726_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .B(_1726_), .Y(_1727_) );
XNOR2X1 XNOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(_1723_), .Y(micro_ucr_hash1_c_24__4_) );
NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1809_), .B(_1813_), .C(_1808_), .Y(_1728_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_1727_), .B(_1719_), .C(_1728_), .Y(_1729_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__5_), .Y(_1730_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__5_), .B(micro_ucr_hash1_a_23__5_), .C(_1730_), .Y(_1731_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__5_), .B(micro_ucr_hash1_a_23__5_), .Y(_1732_) );
NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__5_), .B(_1732_), .Y(_1733_) );
NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1809_), .B(_1731_), .C(_1733_), .Y(_1734_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(_1809_), .Y(_1735_) );
NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_1730_), .B(_1732_), .Y(_1736_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__5_), .B(micro_ucr_hash1_a_23__5_), .C(micro_ucr_hash1_W_24__5_), .Y(_1737_) );
NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_1737_), .B(_1736_), .C(_1735_), .Y(_1738_) );
NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1734_), .B(_1738_), .Y(_1739_) );
XOR2X1 XOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1729_), .B(_1739_), .Y(micro_ucr_hash1_c_24__5_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_23__2_), .C(_1789_), .Y(_1740_) );
NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__2_), .B(_1790_), .Y(_1741_) );
AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1740_), .B(_1741_), .C(_1779_), .Y(_1742_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(_1806_), .Y(_1743_) );
AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1802_), .B(_1742_), .C(_1743_), .Y(_1744_) );
NOR3X1 NOR3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_1784_), .B(_1785_), .C(_1786_), .Y(_1745_) );
NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_1795_), .B(_1802_), .C(_1745_), .Y(_1746_) );
NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(_1723_), .Y(_1747_) );
AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_1744_), .B(_1746_), .C(_1747_), .Y(_1748_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_1737_), .C(_1728_), .D(_1809_), .Y(_1749_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .Y(_1750_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__6_), .B(micro_ucr_hash1_a_23__6_), .C(micro_ucr_hash1_W_24__6_), .Y(_1751_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__6_), .Y(_1752_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__6_), .B(micro_ucr_hash1_a_23__6_), .Y(_1753_) );
NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_1753_), .Y(_1754_) );
NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_1751_), .B(_1754_), .Y(_1755_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1750_), .B(_1755_), .Y(_1756_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(_1756_), .Y(_1757_) );
NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1750_), .B(_1755_), .Y(_1758_) );
NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_1758_), .B(_1757_), .Y(_1759_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(_1759_), .Y(_1760_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_1748_), .B(_1749_), .C(_1760_), .Y(_1761_) );
NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1804_), .B(_1720_), .C(_1721_), .Y(_1762_) );
NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1762_), .B(_1728_), .Y(_1763_) );
AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_1734_), .B(_1738_), .C(_1763_), .Y(_1764_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_1725_), .B(_1726_), .C(_1764_), .Y(_1765_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(_1749_), .Y(_1766_) );
NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1766_), .B(_1759_), .C(_1765_), .Y(_1767_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_1761_), .B(_1767_), .Y(micro_ucr_hash1_c_24__6_) );
AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_1766_), .B(_1765_), .C(_1759_), .Y(_1768_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__7_), .B(micro_ucr_hash1_a_23__7_), .Y(_1769_) );
XNOR2X1 XNOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1769_), .B(micro_ucr_hash1_W_24__7_), .Y(_1770_) );
XNOR2X1 XNOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1770_), .B(_1751_), .Y(_1771_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_1768_), .B(_1756_), .C(_1771_), .Y(_1772_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(_1771_), .Y(_1773_) );
NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1757_), .B(_1773_), .C(_1761_), .Y(_1774_) );
NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1772_), .B(_1774_), .Y(micro_ucr_hash1_c_24__7_) );
XOR2X1 XOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__4_), .B(gnd), .Y(micro_ucr_hash1_a_25__0_) );
XOR2X1 XOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__5_), .B(gnd), .Y(micro_ucr_hash1_a_25__1_) );
XOR2X1 XOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__6_), .B(gnd), .Y(micro_ucr_hash1_a_25__2_) );
XOR2X1 XOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__7_), .B(gnd), .Y(micro_ucr_hash1_a_25__3_) );
XOR2X1 XOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_24__4_), .B(micro_ucr_hash1_b_24__4_), .Y(micro_ucr_hash1_a_25__4_) );
XOR2X1 XOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_24__5_), .B(micro_ucr_hash1_b_24__5_), .Y(micro_ucr_hash1_a_25__5_) );
XOR2X1 XOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_24__6_), .B(micro_ucr_hash1_b_24__6_), .Y(micro_ucr_hash1_a_25__6_) );
XOR2X1 XOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_24__7_), .B(micro_ucr_hash1_b_24__7_), .Y(micro_ucr_hash1_a_25__7_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_25__0_), .Y(_1814_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_24__0_), .Y(_1815_) );
NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_1814_), .B(_1815_), .Y(_1816_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_24__0_), .C(micro_ucr_hash1_W_25__0_), .Y(_1817_) );
NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_1817_), .B(_1816_), .Y(micro_ucr_hash1_b_26__4_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_24__1_), .C(micro_ucr_hash1_W_25__1_), .Y(_1818_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_25__1_), .Y(_1819_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_24__1_), .Y(_1820_) );
NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_1819_), .B(_1820_), .Y(_1821_) );
NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .B(_1816_), .C(_1821_), .Y(_1822_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .B(_1814_), .Y(_1823_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .Y(_1824_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_1820_), .B(_1819_), .Y(_1825_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_1825_), .B(_1824_), .C(_1823_), .Y(_1826_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_1826_), .B(_1822_), .Y(micro_ucr_hash1_b_26__5_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_24__2_), .C(micro_ucr_hash1_W_25__2_), .Y(_1827_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_25__2_), .Y(_1828_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_24__2_), .Y(_1829_) );
NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_1828_), .B(_1829_), .Y(_1830_) );
NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_1830_), .Y(_1831_) );
NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_1830_), .C(_1824_), .Y(_1832_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_1822_), .B(_1831_), .C(_1832_), .Y(_1833_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(_1831_), .Y(_1834_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_1823_), .B(_1825_), .C(_1818_), .Y(_1835_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1835_), .B(_1834_), .Y(_1836_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(_1836_), .Y(micro_ucr_hash1_b_26__6_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_25__3_), .Y(_1837_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_24__3_), .C(_1837_), .Y(_1838_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_24__3_), .Y(_1839_) );
NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_25__3_), .B(_1839_), .Y(_1840_) );
NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_1838_), .C(_1840_), .Y(_1841_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .Y(_1842_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_24__3_), .C(micro_ucr_hash1_W_25__3_), .Y(_1843_) );
NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_1837_), .B(_1839_), .Y(_1844_) );
NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_1843_), .B(_1844_), .C(_1842_), .Y(_1845_) );
NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_1841_), .B(_1845_), .Y(_1846_) );
XNOR2X1 XNOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(_1846_), .Y(micro_ucr_hash1_b_26__7_) );
XOR2X1 XOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_26__4_), .B(gnd), .Y(micro_ucr_hash1_a_26__0_) );
XOR2X1 XOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_26__5_), .B(gnd), .Y(micro_ucr_hash1_a_26__1_) );
XOR2X1 XOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_26__6_), .B(gnd), .Y(micro_ucr_hash1_a_26__2_) );
XOR2X1 XOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_26__7_), .B(gnd), .Y(micro_ucr_hash1_a_26__3_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__0_), .Y(_1903_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__0_), .Y(_1904_) );
NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(_1903_), .B(_1904_), .Y(_1905_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__0_), .C(micro_ucr_hash1_W_26__0_), .Y(_1906_) );
NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_1906_), .B(_1905_), .Y(micro_ucr_hash1_b_27__4_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__1_), .C(micro_ucr_hash1_W_26__1_), .Y(_1907_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__1_), .Y(_1908_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__1_), .Y(_1909_) );
NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_1908_), .B(_1909_), .Y(_1910_) );
NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1907_), .B(_1905_), .C(_1910_), .Y(_1911_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_1904_), .B(_1903_), .Y(_1912_) );
INVX2 INVX2_49 ( .gnd(gnd), .vdd(vdd), .A(_1907_), .Y(_1913_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_1909_), .B(_1908_), .Y(_1914_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_1914_), .B(_1913_), .C(_1912_), .Y(_1915_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_1915_), .B(_1911_), .Y(micro_ucr_hash1_b_27__5_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__2_), .C(micro_ucr_hash1_W_26__2_), .Y(_1916_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__2_), .Y(_1917_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__2_), .Y(_1918_) );
NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_1917_), .B(_1918_), .Y(_1919_) );
NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_1919_), .Y(_1920_) );
NAND3X1 NAND3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_1919_), .C(_1913_), .Y(_1921_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_1911_), .B(_1920_), .C(_1921_), .Y(_1922_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(_1920_), .Y(_1923_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(_1914_), .C(_1907_), .Y(_1924_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1924_), .B(_1923_), .Y(_1925_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1922_), .B(_1925_), .Y(micro_ucr_hash1_b_27__6_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__3_), .Y(_1926_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__3_), .C(_1926_), .Y(_1927_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__3_), .Y(_1928_) );
NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__3_), .B(_1928_), .Y(_1929_) );
NAND3X1 NAND3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .B(_1927_), .C(_1929_), .Y(_1930_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(_1916_), .Y(_1931_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__3_), .C(micro_ucr_hash1_W_26__3_), .Y(_1932_) );
NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(_1928_), .Y(_1933_) );
NAND3X1 NAND3X1_279 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(_1933_), .C(_1931_), .Y(_1934_) );
NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_1934_), .Y(_1935_) );
XNOR2X1 XNOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1922_), .B(_1935_), .Y(micro_ucr_hash1_b_27__7_) );
INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .Y(_1936_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__4_), .B(micro_ucr_hash1_a_25__4_), .C(micro_ucr_hash1_W_26__4_), .Y(_1937_) );
INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__4_), .Y(_1938_) );
INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_25__4_), .Y(_1939_) );
INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__4_), .Y(_1940_) );
NAND3X1 NAND3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_1939_), .C(_1940_), .Y(_1941_) );
AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1937_), .B(_1941_), .C(_1936_), .Y(_1847_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__4_), .B(micro_ucr_hash1_a_25__4_), .C(_1940_), .Y(_1848_) );
NAND3X1 NAND3X1_281 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__4_), .B(_1938_), .C(_1939_), .Y(_1849_) );
AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_1849_), .C(_1932_), .Y(_1850_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1850_), .B(_1847_), .Y(_1851_) );
AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(_1933_), .C(_1931_), .Y(_1852_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_1852_), .B(_1921_), .C(_1934_), .Y(_1853_) );
NOR3X1 NOR3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_1911_), .B(_1920_), .C(_1852_), .Y(_1854_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .B(_1854_), .Y(_1855_) );
XNOR2X1 XNOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_1851_), .Y(micro_ucr_hash1_c_26__4_) );
NAND3X1 NAND3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1937_), .B(_1941_), .C(_1936_), .Y(_1856_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_1855_), .B(_1847_), .C(_1856_), .Y(_1857_) );
INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__5_), .Y(_1858_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__5_), .B(micro_ucr_hash1_a_25__5_), .C(_1858_), .Y(_1859_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__5_), .B(micro_ucr_hash1_a_25__5_), .Y(_1860_) );
NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__5_), .B(_1860_), .Y(_1861_) );
NAND3X1 NAND3X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1937_), .B(_1859_), .C(_1861_), .Y(_1862_) );
INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(_1937_), .Y(_1863_) );
NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_1858_), .B(_1860_), .Y(_1864_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__5_), .B(micro_ucr_hash1_a_25__5_), .C(micro_ucr_hash1_W_26__5_), .Y(_1865_) );
NAND3X1 NAND3X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1865_), .B(_1864_), .C(_1863_), .Y(_1866_) );
NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_1866_), .Y(_1867_) );
XOR2X1 XOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1857_), .B(_1867_), .Y(micro_ucr_hash1_c_26__5_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_25__2_), .C(_1917_), .Y(_1868_) );
NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__2_), .B(_1918_), .Y(_1869_) );
AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1868_), .B(_1869_), .C(_1907_), .Y(_1870_) );
INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(_1934_), .Y(_1871_) );
AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_1870_), .C(_1871_), .Y(_1872_) );
NOR3X1 NOR3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_1912_), .B(_1913_), .C(_1914_), .Y(_1873_) );
NAND3X1 NAND3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1923_), .B(_1930_), .C(_1873_), .Y(_1874_) );
NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1867_), .B(_1851_), .Y(_1875_) );
AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1872_), .B(_1874_), .C(_1875_), .Y(_1876_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1864_), .B(_1865_), .C(_1856_), .D(_1937_), .Y(_1877_) );
INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(_1864_), .Y(_1878_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__6_), .B(micro_ucr_hash1_a_25__6_), .C(micro_ucr_hash1_W_26__6_), .Y(_1879_) );
INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_26__6_), .Y(_1880_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__6_), .B(micro_ucr_hash1_a_25__6_), .Y(_1881_) );
NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_1880_), .B(_1881_), .Y(_1882_) );
NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_1879_), .B(_1882_), .Y(_1883_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1878_), .B(_1883_), .Y(_1884_) );
INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(_1884_), .Y(_1885_) );
NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_1878_), .B(_1883_), .Y(_1886_) );
NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_1886_), .B(_1885_), .Y(_1887_) );
INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(_1887_), .Y(_1888_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_1876_), .B(_1877_), .C(_1888_), .Y(_1889_) );
NAND3X1 NAND3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_1932_), .B(_1848_), .C(_1849_), .Y(_1890_) );
NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_1890_), .B(_1856_), .Y(_1891_) );
AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1862_), .B(_1866_), .C(_1891_), .Y(_1892_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_1853_), .B(_1854_), .C(_1892_), .Y(_1893_) );
INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(_1877_), .Y(_1894_) );
NAND3X1 NAND3X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(_1887_), .C(_1893_), .Y(_1895_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_1889_), .B(_1895_), .Y(micro_ucr_hash1_c_26__6_) );
AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1894_), .B(_1893_), .C(_1887_), .Y(_1896_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__7_), .B(micro_ucr_hash1_a_25__7_), .Y(_1897_) );
XNOR2X1 XNOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1897_), .B(micro_ucr_hash1_W_26__7_), .Y(_1898_) );
XNOR2X1 XNOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1898_), .B(_1879_), .Y(_1899_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .B(_1884_), .C(_1899_), .Y(_1900_) );
INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(_1899_), .Y(_1901_) );
NAND3X1 NAND3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1885_), .B(_1901_), .C(_1889_), .Y(_1902_) );
NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_1900_), .B(_1902_), .Y(micro_ucr_hash1_c_26__7_) );
XOR2X1 XOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__4_), .B(gnd), .Y(micro_ucr_hash1_a_27__0_) );
XOR2X1 XOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__5_), .B(gnd), .Y(micro_ucr_hash1_a_27__1_) );
XOR2X1 XOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__6_), .B(gnd), .Y(micro_ucr_hash1_a_27__2_) );
XOR2X1 XOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__7_), .B(gnd), .Y(micro_ucr_hash1_a_27__3_) );
XOR2X1 XOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_26__4_), .B(micro_ucr_hash1_b_26__4_), .Y(micro_ucr_hash1_a_27__4_) );
XOR2X1 XOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_26__5_), .B(micro_ucr_hash1_b_26__5_), .Y(micro_ucr_hash1_a_27__5_) );
XOR2X1 XOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_26__6_), .B(micro_ucr_hash1_b_26__6_), .Y(micro_ucr_hash1_a_27__6_) );
XOR2X1 XOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_26__7_), .B(micro_ucr_hash1_b_26__7_), .Y(micro_ucr_hash1_a_27__7_) );
INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_27__0_), .Y(_1942_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_26__0_), .Y(_1943_) );
NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_1942_), .B(_1943_), .Y(_1944_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_26__0_), .C(micro_ucr_hash1_W_27__0_), .Y(_1945_) );
NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1945_), .B(_1944_), .Y(micro_ucr_hash1_b_28__4_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_26__1_), .C(micro_ucr_hash1_W_27__1_), .Y(_1946_) );
INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_27__1_), .Y(_1947_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_26__1_), .Y(_1948_) );
NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(_1947_), .B(_1948_), .Y(_1949_) );
NAND3X1 NAND3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .B(_1944_), .C(_1949_), .Y(_1950_) );
AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_1943_), .B(_1942_), .Y(_1951_) );
INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(_1946_), .Y(_1952_) );
AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_1948_), .B(_1947_), .Y(_1953_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_1953_), .B(_1952_), .C(_1951_), .Y(_1954_) );
AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_1954_), .B(_1950_), .Y(micro_ucr_hash1_b_28__5_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_26__2_), .C(micro_ucr_hash1_W_27__2_), .Y(_1955_) );
INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_27__2_), .Y(_1956_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_26__2_), .Y(_1957_) );
NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(_1957_), .Y(_1958_) );
NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_1955_), .B(_1958_), .Y(_1959_) );
NAND3X1 NAND3X1_290 ( .gnd(gnd), .vdd(vdd), .A(_1955_), .B(_1958_), .C(_1952_), .Y(_1960_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_1950_), .B(_1959_), .C(_1960_), .Y(_1961_) );
INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(_1959_), .Y(_1962_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_1951_), .B(_1953_), .C(_1946_), .Y(_1963_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1963_), .B(_1962_), .Y(_1964_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1961_), .B(_1964_), .Y(micro_ucr_hash1_b_28__6_) );
INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_27__3_), .Y(_1965_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_26__3_), .C(_1965_), .Y(_1966_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_26__3_), .Y(_1967_) );
NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_27__3_), .B(_1967_), .Y(_1968_) );
NAND3X1 NAND3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_1955_), .B(_1966_), .C(_1968_), .Y(_1969_) );
INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(_1955_), .Y(_1970_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_26__3_), .C(micro_ucr_hash1_W_27__3_), .Y(_1971_) );
NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_1965_), .B(_1967_), .Y(_1972_) );
NAND3X1 NAND3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1972_), .C(_1970_), .Y(_1973_) );
NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_1969_), .B(_1973_), .Y(_1974_) );
XNOR2X1 XNOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1961_), .B(_1974_), .Y(micro_ucr_hash1_b_28__7_) );
XOR2X1 XOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_28__4_), .B(gnd), .Y(micro_ucr_hash1_a_28__0_) );
XOR2X1 XOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_28__5_), .B(gnd), .Y(micro_ucr_hash1_a_28__1_) );
XOR2X1 XOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_28__6_), .B(gnd), .Y(micro_ucr_hash1_a_28__2_) );
XOR2X1 XOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_28__7_), .B(gnd), .Y(micro_ucr_hash1_a_28__3_) );
INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__0_), .Y(_2031_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__0_), .Y(_2032_) );
NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_2031_), .B(_2032_), .Y(_2033_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__0_), .C(micro_ucr_hash1_W_28__0_), .Y(_2034_) );
NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_2034_), .B(_2033_), .Y(micro_ucr_hash1_b_29__4_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__1_), .C(micro_ucr_hash1_W_28__1_), .Y(_2035_) );
INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__1_), .Y(_2036_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__1_), .Y(_2037_) );
NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(_2037_), .Y(_2038_) );
NAND3X1 NAND3X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2035_), .B(_2033_), .C(_2038_), .Y(_2039_) );
AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_2032_), .B(_2031_), .Y(_2040_) );
INVX2 INVX2_50 ( .gnd(gnd), .vdd(vdd), .A(_2035_), .Y(_2041_) );
AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_2037_), .B(_2036_), .Y(_2042_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2042_), .B(_2041_), .C(_2040_), .Y(_2043_) );
AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_2043_), .B(_2039_), .Y(micro_ucr_hash1_b_29__5_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__2_), .C(micro_ucr_hash1_W_28__2_), .Y(_2044_) );
INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__2_), .Y(_2045_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__2_), .Y(_2046_) );
NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2045_), .B(_2046_), .Y(_2047_) );
NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .B(_2047_), .Y(_2048_) );
NAND3X1 NAND3X1_294 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .B(_2047_), .C(_2041_), .Y(_2049_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2039_), .B(_2048_), .C(_2049_), .Y(_2050_) );
INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(_2048_), .Y(_2051_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(_2042_), .C(_2035_), .Y(_2052_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_2052_), .B(_2051_), .Y(_2053_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_2050_), .B(_2053_), .Y(micro_ucr_hash1_b_29__6_) );
INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__3_), .Y(_2054_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__3_), .C(_2054_), .Y(_2055_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__3_), .Y(_2056_) );
NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__3_), .B(_2056_), .Y(_2057_) );
NAND3X1 NAND3X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .B(_2055_), .C(_2057_), .Y(_2058_) );
INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(_2044_), .Y(_2059_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__3_), .C(micro_ucr_hash1_W_28__3_), .Y(_2060_) );
NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_2054_), .B(_2056_), .Y(_2061_) );
NAND3X1 NAND3X1_296 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(_2061_), .C(_2059_), .Y(_2062_) );
NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_2058_), .B(_2062_), .Y(_2063_) );
XNOR2X1 XNOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_2050_), .B(_2063_), .Y(micro_ucr_hash1_b_29__7_) );
INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .Y(_2064_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__4_), .B(micro_ucr_hash1_a_27__4_), .C(micro_ucr_hash1_W_28__4_), .Y(_2065_) );
INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__4_), .Y(_2066_) );
INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_27__4_), .Y(_2067_) );
INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__4_), .Y(_2068_) );
NAND3X1 NAND3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2066_), .B(_2067_), .C(_2068_), .Y(_2069_) );
AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .B(_2069_), .C(_2064_), .Y(_1975_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__4_), .B(micro_ucr_hash1_a_27__4_), .C(_2068_), .Y(_1976_) );
NAND3X1 NAND3X1_298 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__4_), .B(_2066_), .C(_2067_), .Y(_1977_) );
AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1976_), .B(_1977_), .C(_2060_), .Y(_1978_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1978_), .B(_1975_), .Y(_1979_) );
AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(_2061_), .C(_2059_), .Y(_1980_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_1980_), .B(_2049_), .C(_2062_), .Y(_1981_) );
NOR3X1 NOR3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_2039_), .B(_2048_), .C(_1980_), .Y(_1982_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1981_), .B(_1982_), .Y(_1983_) );
XNOR2X1 XNOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .B(_1979_), .Y(micro_ucr_hash1_c_28__4_) );
NAND3X1 NAND3X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .B(_2069_), .C(_2064_), .Y(_1984_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_1983_), .B(_1975_), .C(_1984_), .Y(_1985_) );
INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__5_), .Y(_1986_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__5_), .B(micro_ucr_hash1_a_27__5_), .C(_1986_), .Y(_1987_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__5_), .B(micro_ucr_hash1_a_27__5_), .Y(_1988_) );
NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__5_), .B(_1988_), .Y(_1989_) );
NAND3X1 NAND3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .B(_1987_), .C(_1989_), .Y(_1990_) );
INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .Y(_1991_) );
NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_1986_), .B(_1988_), .Y(_1992_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__5_), .B(micro_ucr_hash1_a_27__5_), .C(micro_ucr_hash1_W_28__5_), .Y(_1993_) );
NAND3X1 NAND3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_1993_), .B(_1992_), .C(_1991_), .Y(_1994_) );
NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_1994_), .Y(_1995_) );
XOR2X1 XOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1985_), .B(_1995_), .Y(micro_ucr_hash1_c_28__5_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_27__2_), .C(_2045_), .Y(_1996_) );
NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__2_), .B(_2046_), .Y(_1997_) );
AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_1997_), .C(_2035_), .Y(_1998_) );
INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .Y(_1999_) );
AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_2058_), .B(_1998_), .C(_1999_), .Y(_2000_) );
NOR3X1 NOR3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(_2041_), .C(_2042_), .Y(_2001_) );
NAND3X1 NAND3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_2051_), .B(_2058_), .C(_2001_), .Y(_2002_) );
NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_1995_), .B(_1979_), .Y(_2003_) );
AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_2000_), .B(_2002_), .C(_2003_), .Y(_2004_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_1992_), .B(_1993_), .C(_1984_), .D(_2065_), .Y(_2005_) );
INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(_1992_), .Y(_2006_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__6_), .B(micro_ucr_hash1_a_27__6_), .C(micro_ucr_hash1_W_28__6_), .Y(_2007_) );
INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_28__6_), .Y(_2008_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__6_), .B(micro_ucr_hash1_a_27__6_), .Y(_2009_) );
NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_2008_), .B(_2009_), .Y(_2010_) );
NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_2007_), .B(_2010_), .Y(_2011_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(_2011_), .Y(_2012_) );
INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .Y(_2013_) );
NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .B(_2011_), .Y(_2014_) );
NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(_2013_), .Y(_2015_) );
INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(_2015_), .Y(_2016_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(_2005_), .C(_2016_), .Y(_2017_) );
NAND3X1 NAND3X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(_1976_), .C(_1977_), .Y(_2018_) );
NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2018_), .B(_1984_), .Y(_2019_) );
AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_1994_), .C(_2019_), .Y(_2020_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_1981_), .B(_1982_), .C(_2020_), .Y(_2021_) );
INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2022_) );
NAND3X1 NAND3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2022_), .B(_2015_), .C(_2021_), .Y(_2023_) );
AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_2017_), .B(_2023_), .Y(micro_ucr_hash1_c_28__6_) );
AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_2022_), .B(_2021_), .C(_2015_), .Y(_2024_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__7_), .B(micro_ucr_hash1_a_27__7_), .Y(_2025_) );
XNOR2X1 XNOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_2025_), .B(micro_ucr_hash1_W_28__7_), .Y(_2026_) );
XNOR2X1 XNOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_2026_), .B(_2007_), .Y(_2027_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(_2012_), .C(_2027_), .Y(_2028_) );
INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(_2027_), .Y(_2029_) );
NAND3X1 NAND3X1_305 ( .gnd(gnd), .vdd(vdd), .A(_2013_), .B(_2029_), .C(_2017_), .Y(_2030_) );
NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .B(_2030_), .Y(micro_ucr_hash1_c_28__7_) );
XOR2X1 XOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__4_), .B(gnd), .Y(micro_ucr_hash1_a_29__0_) );
XOR2X1 XOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__5_), .B(gnd), .Y(micro_ucr_hash1_a_29__1_) );
XOR2X1 XOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__6_), .B(gnd), .Y(micro_ucr_hash1_a_29__2_) );
XOR2X1 XOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__7_), .B(gnd), .Y(micro_ucr_hash1_a_29__3_) );
XOR2X1 XOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_28__4_), .B(micro_ucr_hash1_b_28__4_), .Y(micro_ucr_hash1_a_29__4_) );
XOR2X1 XOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_28__5_), .B(micro_ucr_hash1_b_28__5_), .Y(micro_ucr_hash1_a_29__5_) );
XOR2X1 XOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_28__6_), .B(micro_ucr_hash1_b_28__6_), .Y(micro_ucr_hash1_a_29__6_) );
XOR2X1 XOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_28__7_), .B(micro_ucr_hash1_b_28__7_), .Y(micro_ucr_hash1_a_29__7_) );
INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_29__0_), .Y(_2070_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_28__0_), .Y(_2071_) );
NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_2070_), .B(_2071_), .Y(_2072_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_28__0_), .C(micro_ucr_hash1_W_29__0_), .Y(_2073_) );
NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_2073_), .B(_2072_), .Y(micro_ucr_hash1_b_30__4_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_28__1_), .C(micro_ucr_hash1_W_29__1_), .Y(_2074_) );
INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_29__1_), .Y(_2075_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_28__1_), .Y(_2076_) );
NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2075_), .B(_2076_), .Y(_2077_) );
NAND3X1 NAND3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2074_), .B(_2072_), .C(_2077_), .Y(_2078_) );
AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_2071_), .B(_2070_), .Y(_2079_) );
INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(_2074_), .Y(_2080_) );
AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_2076_), .B(_2075_), .Y(_2081_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2081_), .B(_2080_), .C(_2079_), .Y(_2082_) );
AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_2082_), .B(_2078_), .Y(micro_ucr_hash1_b_30__5_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_28__2_), .C(micro_ucr_hash1_W_29__2_), .Y(_2083_) );
INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_29__2_), .Y(_2084_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_28__2_), .Y(_2085_) );
NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2084_), .B(_2085_), .Y(_2086_) );
NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2083_), .B(_2086_), .Y(_2087_) );
NAND3X1 NAND3X1_307 ( .gnd(gnd), .vdd(vdd), .A(_2083_), .B(_2086_), .C(_2080_), .Y(_2088_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .B(_2087_), .C(_2088_), .Y(_2089_) );
INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(_2087_), .Y(_2090_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_2079_), .B(_2081_), .C(_2074_), .Y(_2091_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_2091_), .B(_2090_), .Y(_2092_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .B(_2092_), .Y(micro_ucr_hash1_b_30__6_) );
INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_29__3_), .Y(_2093_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_28__3_), .C(_2093_), .Y(_2094_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_28__3_), .Y(_2095_) );
NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_29__3_), .B(_2095_), .Y(_2096_) );
NAND3X1 NAND3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_2083_), .B(_2094_), .C(_2096_), .Y(_2097_) );
INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(_2083_), .Y(_2098_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_28__3_), .C(micro_ucr_hash1_W_29__3_), .Y(_2099_) );
NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_2093_), .B(_2095_), .Y(_2100_) );
NAND3X1 NAND3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .B(_2100_), .C(_2098_), .Y(_2101_) );
NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2097_), .B(_2101_), .Y(_2102_) );
XNOR2X1 XNOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_2089_), .B(_2102_), .Y(micro_ucr_hash1_b_30__7_) );
INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__0_), .Y(_2159_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__0_), .Y(_2160_) );
NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2159_), .B(_2160_), .Y(_2161_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__0_), .C(micro_ucr_hash1_W_30__0_), .Y(_2162_) );
NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2162_), .B(_2161_), .Y(micro_ucr_hash1_b_31__4_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__1_), .C(micro_ucr_hash1_W_30__1_), .Y(_2163_) );
INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__1_), .Y(_2164_) );
NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__1_), .Y(_2165_) );
NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2164_), .B(_2165_), .Y(_2166_) );
NAND3X1 NAND3X1_310 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_2161_), .C(_2166_), .Y(_2167_) );
AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_2160_), .B(_2159_), .Y(_2168_) );
INVX2 INVX2_51 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .Y(_2169_) );
AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_2165_), .B(_2164_), .Y(_2170_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2170_), .B(_2169_), .C(_2168_), .Y(_2171_) );
AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_2171_), .B(_2167_), .Y(micro_ucr_hash1_b_31__5_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__2_), .C(micro_ucr_hash1_W_30__2_), .Y(_2172_) );
INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__2_), .Y(_2173_) );
NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__2_), .Y(_2174_) );
NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2173_), .B(_2174_), .Y(_2175_) );
NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_2172_), .B(_2175_), .Y(_2176_) );
NAND3X1 NAND3X1_311 ( .gnd(gnd), .vdd(vdd), .A(_2172_), .B(_2175_), .C(_2169_), .Y(_2177_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_2167_), .B(_2176_), .C(_2177_), .Y(_2178_) );
INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(_2176_), .Y(_2179_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_2168_), .B(_2170_), .C(_2163_), .Y(_2180_) );
NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_2180_), .B(_2179_), .Y(_2181_) );
NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_2178_), .B(_2181_), .Y(micro_ucr_hash1_b_31__6_) );
INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__3_), .Y(_2182_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__3_), .C(_2182_), .Y(_2183_) );
NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__3_), .Y(_2184_) );
NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__3_), .B(_2184_), .Y(_2185_) );
NAND3X1 NAND3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_2172_), .B(_2183_), .C(_2185_), .Y(_2186_) );
INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(_2172_), .Y(_2187_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__3_), .C(micro_ucr_hash1_W_30__3_), .Y(_2188_) );
NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2182_), .B(_2184_), .Y(_2189_) );
NAND3X1 NAND3X1_313 ( .gnd(gnd), .vdd(vdd), .A(_2188_), .B(_2189_), .C(_2187_), .Y(_2190_) );
NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2190_), .Y(_2191_) );
XNOR2X1 XNOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_2178_), .B(_2191_), .Y(micro_ucr_hash1_b_31__7_) );
INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(_2188_), .Y(_2192_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__4_), .B(micro_ucr_hash1_a_29__4_), .C(micro_ucr_hash1_W_30__4_), .Y(_2193_) );
INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__4_), .Y(_2194_) );
INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_29__4_), .Y(_2195_) );
INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__4_), .Y(_2196_) );
NAND3X1 NAND3X1_314 ( .gnd(gnd), .vdd(vdd), .A(_2194_), .B(_2195_), .C(_2196_), .Y(_2197_) );
AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .B(_2197_), .C(_2192_), .Y(_2103_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__4_), .B(micro_ucr_hash1_a_29__4_), .C(_2196_), .Y(_2104_) );
NAND3X1 NAND3X1_315 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__4_), .B(_2194_), .C(_2195_), .Y(_2105_) );
AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_2104_), .B(_2105_), .C(_2188_), .Y(_2106_) );
NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_2106_), .B(_2103_), .Y(_2107_) );
AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_2188_), .B(_2189_), .C(_2187_), .Y(_2108_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_2108_), .B(_2177_), .C(_2190_), .Y(_2109_) );
NOR3X1 NOR3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_2167_), .B(_2176_), .C(_2108_), .Y(_2110_) );
NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .B(_2110_), .Y(_2111_) );
XNOR2X1 XNOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(_2107_), .Y(micro_ucr_hash1_c_30__4_) );
NAND3X1 NAND3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .B(_2197_), .C(_2192_), .Y(_2112_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_2111_), .B(_2103_), .C(_2112_), .Y(_2113_) );
INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__5_), .Y(_2114_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__5_), .B(micro_ucr_hash1_a_29__5_), .C(_2114_), .Y(_2115_) );
NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__5_), .B(micro_ucr_hash1_a_29__5_), .Y(_2116_) );
NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__5_), .B(_2116_), .Y(_2117_) );
NAND3X1 NAND3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .B(_2115_), .C(_2117_), .Y(_2118_) );
INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .Y(_2119_) );
NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(_2114_), .B(_2116_), .Y(_2120_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__5_), .B(micro_ucr_hash1_a_29__5_), .C(micro_ucr_hash1_W_30__5_), .Y(_2121_) );
NAND3X1 NAND3X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2121_), .B(_2120_), .C(_2119_), .Y(_2122_) );
NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2118_), .B(_2122_), .Y(_2123_) );
XOR2X1 XOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_2113_), .B(_2123_), .Y(micro_ucr_hash1_c_30__5_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(micro_ucr_hash1_a_29__2_), .C(_2173_), .Y(_2124_) );
NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__2_), .B(_2174_), .Y(_2125_) );
AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_2124_), .B(_2125_), .C(_2163_), .Y(_2126_) );
INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(_2190_), .Y(_2127_) );
AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2126_), .C(_2127_), .Y(_2128_) );
NOR3X1 NOR3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_2168_), .B(_2169_), .C(_2170_), .Y(_2129_) );
NAND3X1 NAND3X1_319 ( .gnd(gnd), .vdd(vdd), .A(_2179_), .B(_2186_), .C(_2129_), .Y(_2130_) );
NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_2123_), .B(_2107_), .Y(_2131_) );
AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .B(_2130_), .C(_2131_), .Y(_2132_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .B(_2121_), .C(_2112_), .D(_2193_), .Y(_2133_) );
INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .Y(_2134_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__6_), .B(micro_ucr_hash1_a_29__6_), .C(micro_ucr_hash1_W_30__6_), .Y(_2135_) );
INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_30__6_), .Y(_2136_) );
NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__6_), .B(micro_ucr_hash1_a_29__6_), .Y(_2137_) );
NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_2136_), .B(_2137_), .Y(_2138_) );
NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2135_), .B(_2138_), .Y(_2139_) );
NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_2134_), .B(_2139_), .Y(_2140_) );
INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(_2140_), .Y(_2141_) );
NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_2134_), .B(_2139_), .Y(_2142_) );
NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_2142_), .B(_2141_), .Y(_2143_) );
INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .Y(_2144_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2132_), .B(_2133_), .C(_2144_), .Y(_2145_) );
NAND3X1 NAND3X1_320 ( .gnd(gnd), .vdd(vdd), .A(_2188_), .B(_2104_), .C(_2105_), .Y(_2146_) );
NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_2146_), .B(_2112_), .Y(_2147_) );
AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_2118_), .B(_2122_), .C(_2147_), .Y(_2148_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_2109_), .B(_2110_), .C(_2148_), .Y(_2149_) );
INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .Y(_2150_) );
NAND3X1 NAND3X1_321 ( .gnd(gnd), .vdd(vdd), .A(_2150_), .B(_2143_), .C(_2149_), .Y(_2151_) );
AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_2145_), .B(_2151_), .Y(micro_ucr_hash1_c_30__6_) );
AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_2150_), .B(_2149_), .C(_2143_), .Y(_2152_) );
NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__7_), .B(micro_ucr_hash1_a_29__7_), .Y(_2153_) );
XNOR2X1 XNOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .B(micro_ucr_hash1_W_30__7_), .Y(_2154_) );
XNOR2X1 XNOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_2154_), .B(_2135_), .Y(_2155_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_2152_), .B(_2140_), .C(_2155_), .Y(_2156_) );
INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(_2155_), .Y(_2157_) );
NAND3X1 NAND3X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2141_), .B(_2157_), .C(_2145_), .Y(_2158_) );
NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_2156_), .B(_2158_), .Y(micro_ucr_hash1_c_30__7_) );
XOR2X1 XOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__4_), .B(gnd), .Y(micro_ucr_hash1_a_31__0_) );
XOR2X1 XOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__5_), .B(gnd), .Y(micro_ucr_hash1_a_31__1_) );
XOR2X1 XOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__6_), .B(gnd), .Y(micro_ucr_hash1_a_31__2_) );
XOR2X1 XOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__7_), .B(gnd), .Y(micro_ucr_hash1_a_31__3_) );
XOR2X1 XOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_30__4_), .B(micro_ucr_hash1_b_30__4_), .Y(micro_ucr_hash1_a_31__4_) );
XOR2X1 XOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_30__5_), .B(micro_ucr_hash1_b_30__5_), .Y(micro_ucr_hash1_a_31__5_) );
XOR2X1 XOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_30__6_), .B(micro_ucr_hash1_b_30__6_), .Y(micro_ucr_hash1_a_31__6_) );
XOR2X1 XOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_c_30__7_), .B(micro_ucr_hash1_b_30__7_), .Y(micro_ucr_hash1_a_31__7_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .Y(_2200_) );
INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_0_), .Y(_2201_) );
NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf2), .B(_2201_), .Y(_2199__0_) );
AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(entrada_hash1_contadores_1_), .Y(_2199__1_) );
AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(entrada_hash1_contadores_2_), .Y(_2199__2_) );
INVX2 INVX2_52 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_3_), .Y(_2202_) );
NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf2), .B(_2202_), .Y(_2199__3_) );
INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_4_), .Y(_2203_) );
NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf4), .B(_2203_), .Y(_2199__4_) );
INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_5_), .Y(_2204_) );
NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf2), .B(_2204_), .Y(_2199__5_) );
AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .B(entrada_hash1_contadores_6_), .Y(_2199__6_) );
INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_7_), .Y(_2205_) );
NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf2), .B(_2205_), .Y(_2199__7_) );
AND2X2 AND2X2_127 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf4), .B(entrada_hash1_contadores_8_), .Y(_2199__8_) );
INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_9_), .Y(_2206_) );
NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf1), .B(_2206_), .Y(_2199__9_) );
AND2X2 AND2X2_128 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .B(entrada_hash1_contadores_10_), .Y(_2199__10_) );
AND2X2 AND2X2_129 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .B(entrada_hash1_contadores_11_), .Y(_2199__11_) );
INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_12_), .Y(_2207_) );
NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf4), .B(_2207_), .Y(_2199__12_) );
AND2X2 AND2X2_130 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .B(entrada_hash1_contadores_13_), .Y(_2199__13_) );
INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_14_), .Y(_2208_) );
NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf2), .B(_2208_), .Y(_2199__14_) );
INVX2 INVX2_53 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_15_), .Y(_2209_) );
NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf3), .B(_2209_), .Y(_2199__15_) );
INVX2 INVX2_54 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_16_), .Y(_2210_) );
NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf3), .B(_2210_), .Y(_2199__16_) );
AND2X2 AND2X2_131 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf1), .B(entrada_hash1_contadores_17_), .Y(_2199__17_) );
AND2X2 AND2X2_132 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .B(entrada_hash1_contadores_18_), .Y(_2199__18_) );
INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_19_), .Y(_2211_) );
NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf4), .B(_2211_), .Y(_2199__19_) );
INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_20_), .Y(_2212_) );
NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf2), .B(_2212_), .Y(_2199__20_) );
INVX2 INVX2_55 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_21_), .Y(_2213_) );
NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf4), .B(_2213_), .Y(_2199__21_) );
INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_22_), .Y(_2214_) );
NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf3), .B(_2214_), .Y(_2199__22_) );
INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_23_), .Y(_2215_) );
NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf3), .B(_2215_), .Y(_2199__23_) );
INVX2 INVX2_56 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_24_), .Y(_2216_) );
NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf4), .B(_2216_), .Y(_2199__24_) );
INVX2 INVX2_57 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_25_), .Y(_2217_) );
NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf1), .B(_2217_), .Y(_2199__25_) );
AND2X2 AND2X2_133 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf2), .B(entrada_hash1_contadores_26_), .Y(_2199__26_) );
INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_27_), .Y(_2218_) );
NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf0), .B(_2218_), .Y(_2199__27_) );
INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_28_), .Y(_2219_) );
NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf1), .B(_2219_), .Y(_2199__28_) );
INVX2 INVX2_58 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_29_), .Y(_2220_) );
NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf1), .B(_2220_), .Y(_2199__29_) );
INVX2 INVX2_59 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_30_), .Y(_2221_) );
NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf1), .B(_2221_), .Y(_2199__30_) );
INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_31_), .Y(_2222_) );
NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf0), .B(_2222_), .Y(_2199__31_) );
INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_2223_) );
NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(inicio), .B(_2223_), .Y(_2224_) );
NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_2201_), .B(_2224_), .Y(_2225_) );
INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(inicio), .Y(_2226_) );
NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_2226_), .Y(_2227_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_2227_), .B(entrada_hash1_contadores_0_), .C(reset_bF_buf1), .Y(_2228_) );
NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .B(_2228_), .Y(_2198__0_) );
NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_0_), .B(entrada_hash1_contadores_1_), .Y(_2229_) );
NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .B(_2224_), .Y(_2230_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2225_), .B(entrada_hash1_contadores_1_), .C(reset_bF_buf0), .Y(_2231_) );
NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_2230_), .B(_2231_), .Y(_2198__1_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_2230_), .B(entrada_hash1_contadores_2_), .C(reset_bF_buf0), .Y(_2232_) );
AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_2_), .B(_2230_), .C(_2232_), .Y(_2198__2_) );
NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_2_), .B(_2230_), .Y(_2233_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2233_), .B(_2202_), .C(reset_bF_buf1), .Y(_2234_) );
AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_2202_), .B(_2233_), .C(_2234_), .Y(_2198__3_) );
AND2X2 AND2X2_134 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_2_), .B(entrada_hash1_contadores_3_), .Y(_2235_) );
NAND3X1 NAND3X1_323 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_4_), .B(_2235_), .C(_2230_), .Y(_2236_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(_2236_), .Y(_2237_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_2233_), .B(_2202_), .C(_2203_), .Y(_2238_) );
NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf0), .B(_2238_), .Y(_2239_) );
NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_2237_), .B(_2239_), .Y(_2198__4_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_2237_), .B(entrada_hash1_contadores_5_), .C(reset_bF_buf2), .Y(_2240_) );
AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_5_), .B(_2237_), .C(_2240_), .Y(_2198__5_) );
AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_5_), .B(_2237_), .C(entrada_hash1_contadores_6_), .Y(_2241_) );
NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_5_), .B(entrada_hash1_contadores_6_), .Y(_2242_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2236_), .B(_2242_), .C(reset_bF_buf1), .Y(_2243_) );
NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_2243_), .B(_2241_), .Y(_2198__6_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2236_), .B(_2242_), .C(entrada_hash1_contadores_7_), .Y(_2244_) );
AND2X2 AND2X2_135 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_5_), .B(entrada_hash1_contadores_6_), .Y(_2245_) );
NAND3X1 NAND3X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2205_), .B(_2245_), .C(_2237_), .Y(_2246_) );
AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_2244_), .B(_2246_), .C(_2200__bF_buf4), .Y(_2198__7_) );
NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_4_), .B(entrada_hash1_contadores_7_), .Y(_2247_) );
NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .B(_2247_), .Y(_2248_) );
NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_2_), .B(entrada_hash1_contadores_3_), .Y(_2249_) );
NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_2249_), .B(_2242_), .Y(_2250_) );
NAND3X1 NAND3X1_325 ( .gnd(gnd), .vdd(vdd), .A(_2227_), .B(_2248_), .C(_2250_), .Y(_2251_) );
INVX2 INVX2_60 ( .gnd(gnd), .vdd(vdd), .A(_2251_), .Y(_2252_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2252_), .B(entrada_hash1_contadores_8_), .C(reset_bF_buf4), .Y(_2253_) );
AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_8_), .B(_2252_), .C(_2253_), .Y(_2198__8_) );
NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_8_), .B(_2252_), .Y(_2254_) );
NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_8_), .B(entrada_hash1_contadores_9_), .Y(_2255_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_2251_), .B(_2255_), .C(reset_bF_buf4), .Y(_2256_) );
AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_2206_), .B(_2254_), .C(_2256_), .Y(_2198__9_) );
NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .B(_2251_), .Y(_2257_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_2257_), .B(entrada_hash1_contadores_10_), .C(reset_bF_buf4), .Y(_2258_) );
AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_10_), .B(_2257_), .C(_2258_), .Y(_2198__10_) );
NAND3X1 NAND3X1_326 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_8_), .B(entrada_hash1_contadores_9_), .C(entrada_hash1_contadores_10_), .Y(_2259_) );
NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_2259_), .B(_2251_), .Y(_2260_) );
NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_11_), .B(_2260_), .Y(_2261_) );
NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_11_), .B(_2260_), .Y(_2262_) );
NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf4), .B(_2262_), .Y(_2263_) );
NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_2261_), .B(_2263_), .Y(_2198__11_) );
NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_2207_), .B(_2262_), .Y(_2264_) );
AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_11_), .B(_2260_), .C(entrada_hash1_contadores_12_), .Y(_2265_) );
NOR3X1 NOR3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf0), .B(_2265_), .C(_2264_), .Y(_2198__12_) );
INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(_2259_), .Y(_2266_) );
NAND3X1 NAND3X1_327 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_11_), .B(entrada_hash1_contadores_12_), .C(_2266_), .Y(_2267_) );
NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2267_), .B(_2251_), .Y(_2268_) );
NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_13_), .B(_2268_), .Y(_2269_) );
NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_13_), .B(_2268_), .Y(_2270_) );
NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf4), .B(_2270_), .Y(_2271_) );
NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_2269_), .B(_2271_), .Y(_2198__13_) );
NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2208_), .B(_2270_), .Y(_2272_) );
AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_13_), .B(_2268_), .C(entrada_hash1_contadores_14_), .Y(_2273_) );
NOR3X1 NOR3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf1), .B(_2273_), .C(_2272_), .Y(_2198__14_) );
NAND3X1 NAND3X1_328 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_10_), .B(entrada_hash1_contadores_11_), .C(entrada_hash1_contadores_12_), .Y(_2274_) );
INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(_2274_), .Y(_2275_) );
NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_13_), .B(entrada_hash1_contadores_14_), .Y(_2276_) );
NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .B(_2276_), .Y(_2277_) );
NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2275_), .B(_2277_), .Y(_2278_) );
NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2278_), .B(_2251_), .Y(_2279_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(entrada_hash1_contadores_15_), .C(reset_bF_buf5), .Y(_2280_) );
AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_15_), .B(_2279_), .C(_2280_), .Y(_2198__15_) );
INVX2 INVX2_61 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .Y(_2281_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_2281_), .B(_2209_), .C(_2210_), .Y(_2282_) );
NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2209_), .B(_2210_), .Y(_2283_) );
AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_2283_), .B(_2279_), .C(_2200__bF_buf3), .Y(_2284_) );
AND2X2 AND2X2_136 ( .gnd(gnd), .vdd(vdd), .A(_2282_), .B(_2284_), .Y(_2198__16_) );
AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_2283_), .B(_2279_), .C(entrada_hash1_contadores_17_), .Y(_2285_) );
NAND3X1 NAND3X1_329 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_15_), .B(entrada_hash1_contadores_16_), .C(entrada_hash1_contadores_17_), .Y(_2286_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2281_), .B(_2286_), .C(reset_bF_buf5), .Y(_2287_) );
NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_2285_), .B(_2287_), .Y(_2198__17_) );
INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(_2286_), .Y(_2288_) );
AND2X2 AND2X2_137 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(_2288_), .Y(_2289_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_2289_), .B(entrada_hash1_contadores_18_), .C(reset_bF_buf5), .Y(_2290_) );
AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_18_), .B(_2289_), .C(_2290_), .Y(_2198__18_) );
NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_18_), .B(_2289_), .Y(_2291_) );
NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_18_), .B(entrada_hash1_contadores_19_), .Y(_2292_) );
NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2292_), .B(_2286_), .Y(_2293_) );
NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2279_), .Y(_2294_) );
NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf5), .B(_2294_), .Y(_2295_) );
AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_2211_), .B(_2291_), .C(_2295_), .Y(_2198__19_) );
AND2X2 AND2X2_138 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(_2293_), .Y(_2296_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_2296_), .B(entrada_hash1_contadores_20_), .C(reset_bF_buf1), .Y(_2297_) );
AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_20_), .B(_2296_), .C(_2297_), .Y(_2198__20_) );
NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_20_), .B(_2296_), .Y(_2298_) );
NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_2212_), .B(_2213_), .Y(_2299_) );
NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .B(_2293_), .Y(_2300_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_2281_), .B(_2300_), .C(reset_bF_buf5), .Y(_2301_) );
AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_2213_), .B(_2298_), .C(_2301_), .Y(_2198__21_) );
INVX2 INVX2_62 ( .gnd(gnd), .vdd(vdd), .A(_2300_), .Y(_2302_) );
AND2X2 AND2X2_139 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(_2302_), .Y(_2303_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2303_), .B(entrada_hash1_contadores_22_), .C(reset_bF_buf1), .Y(_2304_) );
AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_22_), .B(_2303_), .C(_2304_), .Y(_2198__22_) );
NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_2302_), .B(_2279_), .Y(_2305_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_2305_), .B(_2214_), .C(entrada_hash1_contadores_23_), .Y(_2306_) );
NAND3X1 NAND3X1_330 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_22_), .B(_2215_), .C(_2303_), .Y(_2307_) );
AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_2306_), .B(_2307_), .C(_2200__bF_buf3), .Y(_2198__23_) );
NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_22_), .B(entrada_hash1_contadores_23_), .Y(_2308_) );
NOR3X1 NOR3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_2226_), .B(_101_), .C(_2308_), .Y(_2309_) );
NAND3X1 NAND3X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2248_), .B(_2250_), .C(_2309_), .Y(_2310_) );
NOR3X1 NOR3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_2300_), .B(_2278_), .C(_2310_), .Y(_2311_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_2311_), .B(entrada_hash1_contadores_24_), .C(reset_bF_buf5), .Y(_2312_) );
AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_24_), .B(_2311_), .C(_2312_), .Y(_2198__24_) );
INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(_2278_), .Y(_2313_) );
OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .B(_2247_), .Y(_2314_) );
NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_2235_), .B(_2245_), .Y(_2315_) );
AND2X2 AND2X2_140 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_22_), .B(entrada_hash1_contadores_23_), .Y(_2316_) );
NAND3X1 NAND3X1_332 ( .gnd(gnd), .vdd(vdd), .A(inicio), .B(_2223_), .C(_2316_), .Y(_2317_) );
NOR3X1 NOR3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2314_), .B(_2315_), .C(_2317_), .Y(_2318_) );
NAND3X1 NAND3X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2313_), .B(_2318_), .C(_2302_), .Y(_2319_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .B(_2216_), .C(_2217_), .Y(_2320_) );
NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2216_), .B(_2217_), .Y(_2321_) );
AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_2321_), .B(_2311_), .C(_2200__bF_buf0), .Y(_2322_) );
AND2X2 AND2X2_141 ( .gnd(gnd), .vdd(vdd), .A(_2320_), .B(_2322_), .Y(_2198__25_) );
AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_2321_), .B(_2311_), .C(entrada_hash1_contadores_26_), .Y(_2323_) );
NAND3X1 NAND3X1_334 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_24_), .B(entrada_hash1_contadores_25_), .C(entrada_hash1_contadores_26_), .Y(_2324_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_2319_), .B(_2324_), .C(reset_bF_buf3), .Y(_2325_) );
NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2323_), .B(_2325_), .Y(_2198__26_) );
NOR3X1 NOR3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_2218_), .B(_2324_), .C(_2319_), .Y(_2326_) );
INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(_2324_), .Y(_2327_) );
AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_2327_), .B(_2311_), .C(entrada_hash1_contadores_27_), .Y(_2328_) );
NOR3X1 NOR3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf0), .B(_2328_), .C(_2326_), .Y(_2198__27_) );
NAND3X1 NAND3X1_335 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_27_), .B(_2327_), .C(_2311_), .Y(_2329_) );
NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_2248_), .B(_2250_), .Y(_2330_) );
NOR3X1 NOR3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_2278_), .B(_2317_), .C(_2330_), .Y(_2331_) );
NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_27_), .B(entrada_hash1_contadores_28_), .Y(_2332_) );
NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2332_), .B(_2324_), .Y(_2333_) );
NAND3X1 NAND3X1_336 ( .gnd(gnd), .vdd(vdd), .A(_2302_), .B(_2333_), .C(_2331_), .Y(_2334_) );
NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(reset_bF_buf3), .B(_2334_), .Y(_2335_) );
AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_2219_), .B(_2329_), .C(_2335_), .Y(_2198__28_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_2334_), .B(_2220_), .C(reset_bF_buf3), .Y(_2336_) );
AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_2220_), .B(_2334_), .C(_2336_), .Y(_2198__29_) );
NAND3X1 NAND3X1_337 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_29_), .B(_2333_), .C(_2311_), .Y(_2337_) );
NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_29_), .B(entrada_hash1_contadores_30_), .Y(_2338_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_2334_), .B(_2338_), .C(reset_bF_buf3), .Y(_2339_) );
AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_2221_), .B(_2337_), .C(_2339_), .Y(_2198__30_) );
NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_contadores_29_), .B(_2333_), .Y(_2340_) );
NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2221_), .B(_2340_), .Y(_2341_) );
AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_2341_), .B(_2311_), .C(entrada_hash1_contadores_31_), .Y(_2342_) );
OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_2340_), .B(_2221_), .Y(_2343_) );
NOR3X1 NOR3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_2222_), .B(_2343_), .C(_2319_), .Y(_2344_) );
NOR3X1 NOR3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_2200__bF_buf0), .B(_2342_), .C(_2344_), .Y(_2198__31_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2199__0_), .Q(entrada_hash1_nonce_0_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2199__1_), .Q(entrada_hash1_nonce_1_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2199__2_), .Q(entrada_hash1_nonce_2_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2199__3_), .Q(entrada_hash1_nonce_3_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2199__4_), .Q(entrada_hash1_nonce_4_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2199__5_), .Q(entrada_hash1_nonce_5_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2199__6_), .Q(entrada_hash1_nonce_6_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2199__7_), .Q(entrada_hash1_nonce_7_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2199__8_), .Q(entrada_hash1_nonce_8_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2199__9_), .Q(entrada_hash1_nonce_9_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2199__10_), .Q(entrada_hash1_nonce_10_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2199__11_), .Q(entrada_hash1_nonce_11_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2199__12_), .Q(entrada_hash1_nonce_12_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2199__13_), .Q(entrada_hash1_nonce_13_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2199__14_), .Q(entrada_hash1_nonce_14_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2199__15_), .Q(entrada_hash1_nonce_15_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2199__16_), .Q(entrada_hash1_nonce_16_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2199__17_), .Q(entrada_hash1_nonce_17_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2199__18_), .Q(entrada_hash1_nonce_18_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2199__19_), .Q(entrada_hash1_nonce_19_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2199__20_), .Q(entrada_hash1_nonce_20_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_2199__21_), .Q(entrada_hash1_nonce_21_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2199__22_), .Q(entrada_hash1_nonce_22_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2199__23_), .Q(entrada_hash1_nonce_23_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2199__24_), .Q(entrada_hash1_nonce_24_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2199__25_), .Q(entrada_hash1_nonce_25_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2199__26_), .Q(entrada_hash1_nonce_26_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2199__27_), .Q(entrada_hash1_nonce_27_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2199__28_), .Q(entrada_hash1_nonce_28_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2199__29_), .Q(entrada_hash1_nonce_29_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2199__30_), .Q(entrada_hash1_nonce_30_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2199__31_), .Q(entrada_hash1_nonce_31_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2198__0_), .Q(entrada_hash1_contadores_0_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2198__1_), .Q(entrada_hash1_contadores_1_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2198__2_), .Q(entrada_hash1_contadores_2_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2198__3_), .Q(entrada_hash1_contadores_3_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2198__4_), .Q(entrada_hash1_contadores_4_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2198__5_), .Q(entrada_hash1_contadores_5_) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2198__6_), .Q(entrada_hash1_contadores_6_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_2198__7_), .Q(entrada_hash1_contadores_7_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2198__8_), .Q(entrada_hash1_contadores_8_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2198__9_), .Q(entrada_hash1_contadores_9_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2198__10_), .Q(entrada_hash1_contadores_10_) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2198__11_), .Q(entrada_hash1_contadores_11_) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2198__12_), .Q(entrada_hash1_contadores_12_) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_2198__13_), .Q(entrada_hash1_contadores_13_) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2198__14_), .Q(entrada_hash1_contadores_14_) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2198__15_), .Q(entrada_hash1_contadores_15_) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2198__16_), .Q(entrada_hash1_contadores_16_) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2198__17_), .Q(entrada_hash1_contadores_17_) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2198__18_), .Q(entrada_hash1_contadores_18_) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2198__19_), .Q(entrada_hash1_contadores_19_) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2198__20_), .Q(entrada_hash1_contadores_20_) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2198__21_), .Q(entrada_hash1_contadores_21_) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_2198__22_), .Q(entrada_hash1_contadores_22_) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2198__23_), .Q(entrada_hash1_contadores_23_) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2198__24_), .Q(entrada_hash1_contadores_24_) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2198__25_), .Q(entrada_hash1_contadores_25_) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_2198__26_), .Q(entrada_hash1_contadores_26_) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2198__27_), .Q(entrada_hash1_contadores_27_) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2198__28_), .Q(entrada_hash1_contadores_28_) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2198__29_), .Q(entrada_hash1_contadores_29_) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2198__30_), .Q(entrada_hash1_contadores_30_) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_2198__31_), .Q(entrada_hash1_contadores_31_) );
INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[24]), .Y(_2345_) );
AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[64]), .B(_2345_), .C(entrada_hash1_nonce_8_), .Y(_2346_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[64]), .B(_2345_), .C(_2346_), .Y(micro_ucr_hash1_W_17__0_) );
INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[25]), .Y(_2347_) );
AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[65]), .B(_2347_), .C(entrada_hash1_nonce_9_), .Y(_2348_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[65]), .B(_2347_), .C(_2348_), .Y(micro_ucr_hash1_W_17__1_) );
INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[26]), .Y(_2349_) );
AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[66]), .B(_2349_), .C(entrada_hash1_nonce_10_), .Y(_2350_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[66]), .B(_2349_), .C(_2350_), .Y(micro_ucr_hash1_W_17__2_) );
INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[27]), .Y(_2351_) );
AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[67]), .B(_2351_), .C(entrada_hash1_nonce_11_), .Y(_2352_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[67]), .B(_2351_), .C(_2352_), .Y(micro_ucr_hash1_W_17__3_) );
INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[28]), .Y(_2353_) );
AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[68]), .B(_2353_), .C(entrada_hash1_nonce_12_), .Y(_2354_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[68]), .B(_2353_), .C(_2354_), .Y(micro_ucr_hash1_W_17__4_) );
INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[29]), .Y(_2355_) );
AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[69]), .B(_2355_), .C(entrada_hash1_nonce_13_), .Y(_2356_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[69]), .B(_2355_), .C(_2356_), .Y(micro_ucr_hash1_W_17__5_) );
INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[30]), .Y(_2357_) );
AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[70]), .B(_2357_), .C(entrada_hash1_nonce_14_), .Y(_2358_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[70]), .B(_2357_), .C(_2358_), .Y(micro_ucr_hash1_W_17__6_) );
INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[31]), .Y(_2359_) );
AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[71]), .B(_2359_), .C(entrada_hash1_nonce_15_), .Y(_2360_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[71]), .B(_2359_), .C(_2360_), .Y(micro_ucr_hash1_W_17__7_) );
INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_16_), .Y(_2361_) );
OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[72]), .B(bloque_bytes[32]), .Y(_2362_) );
NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[72]), .B(bloque_bytes[32]), .Y(_2363_) );
NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_2363_), .B(_2362_), .Y(_2364_) );
NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_2361_), .B(_2364_), .Y(micro_ucr_hash1_W_16__0_) );
INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_17_), .Y(_2365_) );
OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[73]), .B(bloque_bytes[33]), .Y(_2366_) );
NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[73]), .B(bloque_bytes[33]), .Y(_2367_) );
NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_2367_), .B(_2366_), .Y(_2368_) );
NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(_2365_), .B(_2368_), .Y(micro_ucr_hash1_W_16__1_) );
INVX2 INVX2_63 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[34]), .Y(_2369_) );
AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[74]), .B(_2369_), .C(entrada_hash1_nonce_18_), .Y(_2370_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[74]), .B(_2369_), .C(_2370_), .Y(micro_ucr_hash1_W_16__2_) );
INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_19_), .Y(_2371_) );
OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[75]), .B(bloque_bytes[35]), .Y(_2372_) );
NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[75]), .B(bloque_bytes[35]), .Y(_2373_) );
NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2373_), .B(_2372_), .Y(_2374_) );
NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2371_), .B(_2374_), .Y(micro_ucr_hash1_W_16__3_) );
INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_20_), .Y(_2375_) );
OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[76]), .B(bloque_bytes[36]), .Y(_2376_) );
NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[76]), .B(bloque_bytes[36]), .Y(_2377_) );
NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_2377_), .B(_2376_), .Y(_2378_) );
NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2375_), .B(_2378_), .Y(micro_ucr_hash1_W_16__4_) );
INVX2 INVX2_64 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[37]), .Y(_2379_) );
AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[77]), .B(_2379_), .C(entrada_hash1_nonce_21_), .Y(_2380_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[77]), .B(_2379_), .C(_2380_), .Y(micro_ucr_hash1_W_16__5_) );
INVX2 INVX2_65 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[38]), .Y(_2381_) );
AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[78]), .B(_2381_), .C(entrada_hash1_nonce_22_), .Y(_2382_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[78]), .B(_2381_), .C(_2382_), .Y(micro_ucr_hash1_W_16__6_) );
INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[39]), .Y(_2383_) );
AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[79]), .B(_2383_), .C(entrada_hash1_nonce_23_), .Y(_2384_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[79]), .B(_2383_), .C(_2384_), .Y(micro_ucr_hash1_W_16__7_) );
INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[56]), .Y(_2385_) );
INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_0_), .Y(_2386_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_2385_), .B(bloque_bytes[16]), .C(_2386_), .Y(_2387_) );
AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_2385_), .B(bloque_bytes[16]), .C(_2387_), .Y(_2388_) );
INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(_2388_), .Y(micro_ucr_hash1_W_18__0_) );
INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[57]), .Y(_2389_) );
INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_1_), .Y(_2390_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(bloque_bytes[17]), .C(_2390_), .Y(_2391_) );
AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(bloque_bytes[17]), .C(_2391_), .Y(_2392_) );
INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(_2392_), .Y(micro_ucr_hash1_W_18__1_) );
INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[58]), .Y(_2393_) );
INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_2_), .Y(_2394_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_2393_), .B(bloque_bytes[18]), .C(_2394_), .Y(_2395_) );
AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_2393_), .B(bloque_bytes[18]), .C(_2395_), .Y(_2396_) );
INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(_2396_), .Y(micro_ucr_hash1_W_18__2_) );
INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[59]), .Y(_2397_) );
INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_3_), .Y(_2398_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_2397_), .B(bloque_bytes[19]), .C(_2398_), .Y(_2399_) );
AOI21X1 AOI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_2397_), .B(bloque_bytes[19]), .C(_2399_), .Y(_2400_) );
INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(_2400_), .Y(micro_ucr_hash1_W_18__3_) );
INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[60]), .Y(_2401_) );
INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_4_), .Y(_2402_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2401_), .B(bloque_bytes[20]), .C(_2402_), .Y(_2403_) );
AOI21X1 AOI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_2401_), .B(bloque_bytes[20]), .C(_2403_), .Y(_2404_) );
INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(_2404_), .Y(micro_ucr_hash1_W_18__4_) );
INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[61]), .Y(_2405_) );
INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_5_), .Y(_2406_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_2405_), .B(bloque_bytes[21]), .C(_2406_), .Y(_2407_) );
AOI21X1 AOI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_2405_), .B(bloque_bytes[21]), .C(_2407_), .Y(_2408_) );
INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(_2408_), .Y(micro_ucr_hash1_W_18__5_) );
INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[62]), .Y(_2409_) );
INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_6_), .Y(_2410_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_2409_), .B(bloque_bytes[22]), .C(_2410_), .Y(_2411_) );
AOI21X1 AOI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_2409_), .B(bloque_bytes[22]), .C(_2411_), .Y(_2412_) );
INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(_2412_), .Y(micro_ucr_hash1_W_18__6_) );
INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[63]), .Y(_2413_) );
INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_7_), .Y(_2414_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_2413_), .B(bloque_bytes[23]), .C(_2414_), .Y(_2415_) );
AOI21X1 AOI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_2413_), .B(bloque_bytes[23]), .C(_2415_), .Y(_2416_) );
INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(_2416_), .Y(micro_ucr_hash1_W_18__7_) );
AOI21X1 AOI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_2363_), .B(_2362_), .C(entrada_hash1_nonce_16_), .Y(_2417_) );
XNOR2X1 XNOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[48]), .B(bloque_bytes[8]), .Y(_2418_) );
NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2418_), .B(_2417_), .Y(micro_ucr_hash1_W_19__0_) );
AOI21X1 AOI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_2367_), .B(_2366_), .C(entrada_hash1_nonce_17_), .Y(_2419_) );
XNOR2X1 XNOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[49]), .B(bloque_bytes[9]), .Y(_2420_) );
NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_2420_), .B(_2419_), .Y(micro_ucr_hash1_W_19__1_) );
INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[74]), .Y(_2421_) );
INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_18_), .Y(_2422_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_2421_), .B(bloque_bytes[34]), .C(_2422_), .Y(_2423_) );
AOI21X1 AOI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_2421_), .B(bloque_bytes[34]), .C(_2423_), .Y(_2424_) );
XNOR2X1 XNOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[50]), .B(bloque_bytes[10]), .Y(_2425_) );
NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_2425_), .B(_2424_), .Y(micro_ucr_hash1_W_19__2_) );
AOI21X1 AOI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_2373_), .B(_2372_), .C(entrada_hash1_nonce_19_), .Y(_2426_) );
XNOR2X1 XNOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[51]), .B(bloque_bytes[11]), .Y(_2427_) );
NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2427_), .B(_2426_), .Y(micro_ucr_hash1_W_19__3_) );
AOI21X1 AOI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_2377_), .B(_2376_), .C(entrada_hash1_nonce_20_), .Y(_2428_) );
XNOR2X1 XNOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[52]), .B(bloque_bytes[12]), .Y(_2429_) );
NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_2429_), .B(_2428_), .Y(micro_ucr_hash1_W_19__4_) );
INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[77]), .Y(_2430_) );
INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_21_), .Y(_2431_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_2430_), .B(bloque_bytes[37]), .C(_2431_), .Y(_2432_) );
AOI21X1 AOI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_2430_), .B(bloque_bytes[37]), .C(_2432_), .Y(_2433_) );
AND2X2 AND2X2_142 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[53]), .B(bloque_bytes[13]), .Y(_2434_) );
NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[53]), .B(bloque_bytes[13]), .Y(_2435_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_2434_), .B(_2435_), .C(_2433_), .Y(micro_ucr_hash1_W_19__5_) );
XOR2X1 XOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[54]), .B(bloque_bytes[14]), .Y(_2436_) );
INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[79]), .Y(_2437_) );
NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[39]), .B(_2437_), .Y(_2438_) );
AND2X2 AND2X2_143 ( .gnd(gnd), .vdd(vdd), .A(_2384_), .B(_2438_), .Y(_2439_) );
XNOR2X1 XNOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[55]), .B(bloque_bytes[15]), .Y(_2440_) );
XOR2X1 XOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[64]), .B(bloque_bytes[24]), .Y(_2441_) );
NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_8_), .B(_2441_), .Y(_2442_) );
XNOR2X1 XNOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[40]), .B(bloque_bytes[0]), .Y(_2443_) );
NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .B(_2442_), .Y(micro_ucr_hash1_W_20__0_) );
XOR2X1 XOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[65]), .B(bloque_bytes[25]), .Y(_2444_) );
NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_9_), .B(_2444_), .Y(_2445_) );
XNOR2X1 XNOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[41]), .B(bloque_bytes[1]), .Y(_2446_) );
NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .B(_2445_), .Y(micro_ucr_hash1_W_20__1_) );
INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[66]), .Y(_2447_) );
INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_10_), .Y(_2448_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_2447_), .B(bloque_bytes[26]), .C(_2448_), .Y(_2449_) );
AOI21X1 AOI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_2447_), .B(bloque_bytes[26]), .C(_2449_), .Y(_2450_) );
XNOR2X1 XNOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[42]), .B(bloque_bytes[2]), .Y(_2451_) );
NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_2450_), .Y(micro_ucr_hash1_W_20__2_) );
XOR2X1 XOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[43]), .B(bloque_bytes[3]), .Y(_2452_) );
NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2452_), .B(micro_ucr_hash1_W_17__3_), .Y(_2453_) );
INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(_2453_), .Y(micro_ucr_hash1_W_20__3_) );
XOR2X1 XOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[44]), .B(bloque_bytes[4]), .Y(_2454_) );
NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_2454_), .B(micro_ucr_hash1_W_17__4_), .Y(_2455_) );
INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .Y(micro_ucr_hash1_W_20__4_) );
XOR2X1 XOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[45]), .B(bloque_bytes[5]), .Y(_2456_) );
NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2456_), .B(micro_ucr_hash1_W_17__5_), .Y(_2457_) );
INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(_2457_), .Y(micro_ucr_hash1_W_20__5_) );
XOR2X1 XOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[46]), .B(bloque_bytes[6]), .Y(_2458_) );
NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_2458_), .B(micro_ucr_hash1_W_17__6_), .Y(_2459_) );
INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .Y(micro_ucr_hash1_W_20__6_) );
INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[71]), .Y(_2460_) );
INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_15_), .Y(_2461_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .B(bloque_bytes[31]), .C(_2461_), .Y(_2462_) );
AOI21X1 AOI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_2460_), .B(bloque_bytes[31]), .C(_2462_), .Y(_2463_) );
XNOR2X1 XNOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[47]), .B(bloque_bytes[7]), .Y(_2464_) );
NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .B(_2463_), .Y(micro_ucr_hash1_W_20__7_) );
AND2X2 AND2X2_144 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[32]), .B(entrada_hash1_nonce_24_), .Y(_2465_) );
NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[32]), .B(entrada_hash1_nonce_24_), .Y(_2466_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_2465_), .B(_2466_), .C(_2388_), .Y(micro_ucr_hash1_W_21__0_) );
AND2X2 AND2X2_145 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[33]), .B(entrada_hash1_nonce_25_), .Y(_2467_) );
NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[33]), .B(entrada_hash1_nonce_25_), .Y(_2468_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_2467_), .B(_2468_), .C(_2392_), .Y(micro_ucr_hash1_W_21__1_) );
INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_26_), .Y(_2469_) );
NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_2369_), .B(_2469_), .Y(_2470_) );
NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[34]), .B(entrada_hash1_nonce_26_), .Y(_2471_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .B(_2471_), .C(_2396_), .Y(micro_ucr_hash1_W_21__2_) );
AND2X2 AND2X2_146 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[35]), .B(entrada_hash1_nonce_27_), .Y(_2472_) );
NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[35]), .B(entrada_hash1_nonce_27_), .Y(_2473_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_2472_), .B(_2473_), .C(_2400_), .Y(micro_ucr_hash1_W_21__3_) );
AND2X2 AND2X2_147 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[36]), .B(entrada_hash1_nonce_28_), .Y(_2474_) );
NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[36]), .B(entrada_hash1_nonce_28_), .Y(_2475_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_2474_), .B(_2475_), .C(_2404_), .Y(micro_ucr_hash1_W_21__4_) );
INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_29_), .Y(_2476_) );
NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_2379_), .B(_2476_), .Y(_2477_) );
NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[37]), .B(entrada_hash1_nonce_29_), .Y(_2478_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_2477_), .B(_2478_), .C(_2408_), .Y(micro_ucr_hash1_W_21__5_) );
INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_30_), .Y(_2479_) );
NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_2381_), .B(_2479_), .Y(_2480_) );
NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[38]), .B(entrada_hash1_nonce_30_), .Y(_2481_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_2480_), .B(_2481_), .C(_2412_), .Y(micro_ucr_hash1_W_21__6_) );
XNOR2X1 XNOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[39]), .B(entrada_hash1_nonce_31_), .Y(_2482_) );
AND2X2 AND2X2_148 ( .gnd(gnd), .vdd(vdd), .A(_2416_), .B(_2482_), .Y(_2483_) );
XNOR2X1 XNOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[24]), .B(entrada_hash1_nonce_16_), .Y(_2484_) );
NAND3X1 NAND3X1_338 ( .gnd(gnd), .vdd(vdd), .A(_2418_), .B(_2484_), .C(_2417_), .Y(micro_ucr_hash1_W_22__0_) );
XNOR2X1 XNOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[25]), .B(entrada_hash1_nonce_17_), .Y(_2485_) );
NAND3X1 NAND3X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2420_), .B(_2485_), .C(_2419_), .Y(micro_ucr_hash1_W_22__1_) );
XNOR2X1 XNOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[26]), .B(entrada_hash1_nonce_18_), .Y(_2486_) );
NAND3X1 NAND3X1_340 ( .gnd(gnd), .vdd(vdd), .A(_2425_), .B(_2486_), .C(_2424_), .Y(micro_ucr_hash1_W_22__2_) );
XNOR2X1 XNOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[27]), .B(entrada_hash1_nonce_19_), .Y(_2487_) );
NAND3X1 NAND3X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2427_), .B(_2487_), .C(_2426_), .Y(micro_ucr_hash1_W_22__3_) );
XNOR2X1 XNOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[28]), .B(entrada_hash1_nonce_20_), .Y(_2488_) );
NAND3X1 NAND3X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2429_), .B(_2488_), .C(_2428_), .Y(micro_ucr_hash1_W_22__4_) );
XOR2X1 XOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[29]), .B(entrada_hash1_nonce_21_), .Y(_2489_) );
NOR2X1 NOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_2489_), .B(micro_ucr_hash1_W_19__5_), .Y(_2490_) );
INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(_2490_), .Y(micro_ucr_hash1_W_22__5_) );
INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[78]), .Y(_2491_) );
INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_22_), .Y(_2492_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .B(bloque_bytes[38]), .C(_2492_), .Y(_2493_) );
AOI21X1 AOI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .B(bloque_bytes[38]), .C(_2493_), .Y(_2494_) );
INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(_2436_), .Y(_2495_) );
XNOR2X1 XNOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[30]), .B(entrada_hash1_nonce_22_), .Y(_2496_) );
NAND3X1 NAND3X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2495_), .B(_2496_), .C(_2494_), .Y(micro_ucr_hash1_W_22__6_) );
XNOR2X1 XNOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[31]), .B(entrada_hash1_nonce_23_), .Y(_2497_) );
NAND3X1 NAND3X1_344 ( .gnd(gnd), .vdd(vdd), .A(_2440_), .B(_2497_), .C(_2439_), .Y(micro_ucr_hash1_W_22__7_) );
XNOR2X1 XNOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_8_), .B(bloque_bytes[16]), .Y(_2498_) );
NAND3X1 NAND3X1_345 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .B(_2498_), .C(_2442_), .Y(micro_ucr_hash1_W_23__0_) );
XNOR2X1 XNOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_9_), .B(bloque_bytes[17]), .Y(_2499_) );
NAND3X1 NAND3X1_346 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .B(_2499_), .C(_2445_), .Y(micro_ucr_hash1_W_23__1_) );
XNOR2X1 XNOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_10_), .B(bloque_bytes[18]), .Y(_2500_) );
NAND3X1 NAND3X1_347 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_2500_), .C(_2450_), .Y(micro_ucr_hash1_W_23__2_) );
XNOR2X1 XNOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_11_), .B(bloque_bytes[19]), .Y(_2501_) );
AND2X2 AND2X2_149 ( .gnd(gnd), .vdd(vdd), .A(_2453_), .B(_2501_), .Y(_2502_) );
INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(_2502_), .Y(micro_ucr_hash1_W_23__3_) );
XNOR2X1 XNOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_12_), .B(bloque_bytes[20]), .Y(_2503_) );
AND2X2 AND2X2_150 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .B(_2503_), .Y(_2504_) );
XNOR2X1 XNOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_13_), .B(bloque_bytes[21]), .Y(_2505_) );
AND2X2 AND2X2_151 ( .gnd(gnd), .vdd(vdd), .A(_2457_), .B(_2505_), .Y(_2506_) );
XNOR2X1 XNOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_14_), .B(bloque_bytes[22]), .Y(_2507_) );
AND2X2 AND2X2_152 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .B(_2507_), .Y(_2508_) );
XNOR2X1 XNOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_15_), .B(bloque_bytes[23]), .Y(_2509_) );
NAND3X1 NAND3X1_348 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .B(_2509_), .C(_2463_), .Y(micro_ucr_hash1_W_23__7_) );
OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_21__0_), .B(bloque_bytes[8]), .Y(micro_ucr_hash1_W_24__0_) );
OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_21__1_), .B(bloque_bytes[9]), .Y(micro_ucr_hash1_W_24__1_) );
NOR2X1 NOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[10]), .B(micro_ucr_hash1_W_21__2_), .Y(_2510_) );
INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(_2510_), .Y(micro_ucr_hash1_W_24__2_) );
OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_21__3_), .B(bloque_bytes[11]), .Y(micro_ucr_hash1_W_24__3_) );
OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_21__4_), .B(bloque_bytes[12]), .Y(micro_ucr_hash1_W_24__4_) );
NOR2X1 NOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[13]), .B(micro_ucr_hash1_W_21__5_), .Y(_2511_) );
INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .Y(micro_ucr_hash1_W_24__5_) );
NOR2X1 NOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[14]), .B(micro_ucr_hash1_W_21__6_), .Y(_2512_) );
INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(_2512_), .Y(micro_ucr_hash1_W_24__6_) );
AND2X2 AND2X2_153 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_7_), .B(bloque_bytes[15]), .Y(_2513_) );
NOR2X1 NOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_7_), .B(bloque_bytes[15]), .Y(_2514_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .B(_2514_), .C(_2483_), .Y(micro_ucr_hash1_W_24__7_) );
NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[0]), .B(micro_ucr_hash1_W_16__0_), .Y(_2515_) );
INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[0]), .Y(_2516_) );
NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_2516_), .B(_2417_), .Y(_2517_) );
AOI21X1 AOI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .B(_2515_), .C(micro_ucr_hash1_W_22__0_), .Y(_2518_) );
INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(_2518_), .Y(micro_ucr_hash1_W_25__0_) );
NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[1]), .B(micro_ucr_hash1_W_16__1_), .Y(_2519_) );
INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[1]), .Y(_2520_) );
NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_2520_), .B(_2419_), .Y(_2521_) );
AOI21X1 AOI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .B(_2519_), .C(micro_ucr_hash1_W_22__1_), .Y(_2522_) );
INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(_2522_), .Y(micro_ucr_hash1_W_25__1_) );
NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[2]), .B(micro_ucr_hash1_W_16__2_), .Y(_2523_) );
OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__2_), .B(bloque_bytes[2]), .Y(_2524_) );
AOI21X1 AOI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_2523_), .B(_2524_), .C(micro_ucr_hash1_W_22__2_), .Y(_2525_) );
INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(_2525_), .Y(micro_ucr_hash1_W_25__2_) );
NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[3]), .B(micro_ucr_hash1_W_16__3_), .Y(_2526_) );
INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[3]), .Y(_2527_) );
NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_2527_), .B(_2426_), .Y(_2528_) );
AOI21X1 AOI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2526_), .C(micro_ucr_hash1_W_22__3_), .Y(_2529_) );
INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .Y(micro_ucr_hash1_W_25__3_) );
NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[4]), .B(micro_ucr_hash1_W_16__4_), .Y(_2530_) );
INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[4]), .Y(_2531_) );
NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .B(_2428_), .Y(_2532_) );
AOI21X1 AOI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_2532_), .B(_2530_), .C(micro_ucr_hash1_W_22__4_), .Y(_2533_) );
XNOR2X1 XNOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__5_), .B(bloque_bytes[5]), .Y(_2534_) );
NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[6]), .B(micro_ucr_hash1_W_16__6_), .Y(_2535_) );
OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__6_), .B(bloque_bytes[6]), .Y(_2536_) );
AOI21X1 AOI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .B(_2536_), .C(micro_ucr_hash1_W_22__6_), .Y(_2537_) );
NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[7]), .B(micro_ucr_hash1_W_16__7_), .Y(_2538_) );
OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__7_), .B(bloque_bytes[7]), .Y(_2539_) );
AOI21X1 AOI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_2538_), .B(_2539_), .C(micro_ucr_hash1_W_22__7_), .Y(_2540_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_2441_), .B(entrada_hash1_nonce_8_), .C(entrada_hash1_nonce_24_), .Y(_2541_) );
OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_17__0_), .B(entrada_hash1_nonce_24_), .Y(_2542_) );
AOI21X1 AOI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_2541_), .B(_2542_), .C(micro_ucr_hash1_W_23__0_), .Y(_2543_) );
INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(_2543_), .Y(micro_ucr_hash1_W_26__0_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_2444_), .B(entrada_hash1_nonce_9_), .C(entrada_hash1_nonce_25_), .Y(_2544_) );
OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_17__1_), .B(entrada_hash1_nonce_25_), .Y(_2545_) );
AOI21X1 AOI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_2544_), .B(_2545_), .C(micro_ucr_hash1_W_23__1_), .Y(_2546_) );
INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(_2546_), .Y(micro_ucr_hash1_W_26__1_) );
NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_26_), .B(micro_ucr_hash1_W_17__2_), .Y(_2547_) );
NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2469_), .B(_2450_), .Y(_2548_) );
AOI21X1 AOI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_2547_), .B(_2548_), .C(micro_ucr_hash1_W_23__2_), .Y(_2549_) );
INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(_2549_), .Y(micro_ucr_hash1_W_26__2_) );
INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_27_), .Y(_2550_) );
NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_2502_), .Y(micro_ucr_hash1_W_26__3_) );
INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_28_), .Y(_2551_) );
NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_2551_), .B(_2504_), .Y(micro_ucr_hash1_W_26__4_) );
NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_2476_), .B(_2506_), .Y(micro_ucr_hash1_W_26__5_) );
NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_2479_), .B(_2508_), .Y(micro_ucr_hash1_W_26__6_) );
NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_31_), .B(micro_ucr_hash1_W_17__7_), .Y(_2552_) );
OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_17__7_), .B(entrada_hash1_nonce_31_), .Y(_2553_) );
AOI21X1 AOI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .B(_2553_), .C(micro_ucr_hash1_W_23__7_), .Y(_2554_) );
INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(_2554_), .Y(micro_ucr_hash1_W_26__7_) );
OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__0_), .B(entrada_hash1_nonce_16_), .Y(micro_ucr_hash1_W_27__0_) );
OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__1_), .B(entrada_hash1_nonce_17_), .Y(micro_ucr_hash1_W_27__1_) );
NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_2422_), .B(_2510_), .Y(micro_ucr_hash1_W_27__2_) );
OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__3_), .B(entrada_hash1_nonce_19_), .Y(micro_ucr_hash1_W_27__3_) );
XNOR2X1 XNOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_19__0_), .B(entrada_hash1_nonce_8_), .Y(_2555_) );
NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_2518_), .B(_2555_), .Y(micro_ucr_hash1_W_28__0_) );
XNOR2X1 XNOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_19__1_), .B(entrada_hash1_nonce_9_), .Y(_2556_) );
NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_2522_), .B(_2556_), .Y(micro_ucr_hash1_W_28__1_) );
NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_2448_), .B(_2525_), .Y(micro_ucr_hash1_W_28__2_) );
XNOR2X1 XNOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_19__3_), .B(entrada_hash1_nonce_11_), .Y(_2557_) );
NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_2529_), .B(_2557_), .Y(micro_ucr_hash1_W_28__3_) );
XNOR2X1 XNOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_19__4_), .B(entrada_hash1_nonce_12_), .Y(_2558_) );
NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_2533_), .B(_2558_), .Y(micro_ucr_hash1_W_28__4_) );
INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_13_), .Y(_2559_) );
NAND3X1 NAND3X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2559_), .B(_2534_), .C(_2490_), .Y(micro_ucr_hash1_W_28__5_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_16__6_), .B(_2436_), .C(entrada_hash1_nonce_14_), .Y(_2560_) );
INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_14_), .Y(_2561_) );
NAND3X1 NAND3X1_350 ( .gnd(gnd), .vdd(vdd), .A(_2561_), .B(_2495_), .C(_2494_), .Y(_2562_) );
NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_2560_), .B(_2562_), .Y(_2563_) );
NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_2563_), .B(_2537_), .Y(micro_ucr_hash1_W_28__6_) );
NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_2461_), .B(_2540_), .Y(micro_ucr_hash1_W_28__7_) );
AOI21X1 AOI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .B(_2442_), .C(_2386_), .Y(_2564_) );
NOR2X1 NOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_0_), .B(micro_ucr_hash1_W_20__0_), .Y(_2565_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2565_), .B(_2564_), .C(_2543_), .Y(micro_ucr_hash1_W_29__0_) );
AOI21X1 AOI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_2446_), .B(_2445_), .C(_2390_), .Y(_2566_) );
NOR2X1 NOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_1_), .B(micro_ucr_hash1_W_20__1_), .Y(_2567_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_2567_), .B(_2566_), .C(_2546_), .Y(micro_ucr_hash1_W_29__1_) );
AOI21X1 AOI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_2450_), .C(_2394_), .Y(_2568_) );
NOR2X1 NOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(entrada_hash1_nonce_2_), .B(micro_ucr_hash1_W_20__2_), .Y(_2569_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_2569_), .B(_2568_), .C(_2549_), .Y(micro_ucr_hash1_W_29__2_) );
NAND3X1 NAND3X1_351 ( .gnd(gnd), .vdd(vdd), .A(_2398_), .B(_2550_), .C(_2502_), .Y(micro_ucr_hash1_W_29__3_) );
OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__0_), .B(micro_ucr_hash1_W_16__0_), .Y(micro_ucr_hash1_W_30__0_) );
OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__1_), .B(micro_ucr_hash1_W_16__1_), .Y(micro_ucr_hash1_W_30__1_) );
NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_2424_), .B(_2510_), .Y(micro_ucr_hash1_W_30__2_) );
OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__3_), .B(micro_ucr_hash1_W_16__3_), .Y(micro_ucr_hash1_W_30__3_) );
OR2X2 OR2X2_112 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__4_), .B(micro_ucr_hash1_W_16__4_), .Y(micro_ucr_hash1_W_30__4_) );
NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(_2511_), .Y(micro_ucr_hash1_W_30__5_) );
NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_2494_), .B(_2512_), .Y(micro_ucr_hash1_W_30__6_) );
OR2X2 OR2X2_113 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_W_24__7_), .B(micro_ucr_hash1_W_16__7_), .Y(micro_ucr_hash1_W_30__7_) );
AND2X2 AND2X2_154 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__0_), .B(micro_ucr_hash1_a_31__1_), .Y(_2570_) );
NOR2X1 NOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__0_), .B(micro_ucr_hash1_a_31__1_), .Y(_2571_) );
NOR2X1 NOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .B(_2570_), .Y(micro_ucr_hash1_hash_17_) );
INVX2 INVX2_66 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__2_), .Y(_2572_) );
XNOR2X1 XNOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_2570_), .B(_2572_), .Y(micro_ucr_hash1_hash_18_) );
NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__2_), .B(_2570_), .Y(_2573_) );
XNOR2X1 XNOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .B(micro_ucr_hash1_a_31__3_), .Y(micro_ucr_hash1_hash_19_) );
INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__3_), .Y(_2574_) );
NOR2X1 NOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_2572_), .B(_2574_), .Y(_2575_) );
NAND3X1 NAND3X1_352 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__4_), .B(_2570_), .C(_2575_), .Y(_2576_) );
INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__4_), .Y(_2577_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .B(_2574_), .C(_2577_), .Y(_2578_) );
AND2X2 AND2X2_155 ( .gnd(gnd), .vdd(vdd), .A(_2578_), .B(_2576_), .Y(micro_ucr_hash1_hash_20_) );
XNOR2X1 XNOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_2576_), .B(micro_ucr_hash1_a_31__5_), .Y(micro_ucr_hash1_hash_21_) );
AND2X2 AND2X2_156 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__4_), .B(micro_ucr_hash1_a_31__5_), .Y(_2579_) );
NAND3X1 NAND3X1_353 ( .gnd(gnd), .vdd(vdd), .A(_2570_), .B(_2579_), .C(_2575_), .Y(_2580_) );
XNOR2X1 XNOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_2580_), .B(micro_ucr_hash1_a_31__6_), .Y(micro_ucr_hash1_hash_22_) );
INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__6_), .Y(_2581_) );
NOR2X1 NOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2581_), .B(_2580_), .Y(_2582_) );
XOR2X1 XOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_2582_), .B(micro_ucr_hash1_a_31__7_), .Y(micro_ucr_hash1_hash_23_) );
INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_a_31__0_), .Y(micro_ucr_hash1_hash_16_) );
INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_hash_8_) );
NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2583_) );
INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(_2583_), .Y(_2584_) );
NOR2X1 NOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2585_) );
NOR2X1 NOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2585_), .B(_2584_), .Y(micro_ucr_hash1_hash_9_) );
XNOR2X1 XNOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_2583_), .B(gnd), .Y(micro_ucr_hash1_hash_10_) );
INVX2 INVX2_67 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_2586_) );
NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_2584_), .Y(_2587_) );
XNOR2X1 XNOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_2587_), .B(_2586_), .Y(micro_ucr_hash1_hash_11_) );
INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_2588_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_2583_), .B(_2588_), .C(_2586_), .Y(_2589_) );
XOR2X1 XOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .B(micro_ucr_hash1_b_31__4_), .Y(micro_ucr_hash1_hash_12_) );
AND2X2 AND2X2_157 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .B(micro_ucr_hash1_b_31__4_), .Y(_2590_) );
AND2X2 AND2X2_158 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .B(micro_ucr_hash1_b_31__5_), .Y(_2591_) );
NOR2X1 NOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__5_), .B(_2590_), .Y(_2592_) );
NOR2X1 NOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(_2592_), .B(_2591_), .Y(micro_ucr_hash1_hash_13_) );
XOR2X1 XOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_2591_), .B(micro_ucr_hash1_b_31__6_), .Y(micro_ucr_hash1_hash_14_) );
NAND3X1 NAND3X1_354 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__5_), .B(micro_ucr_hash1_b_31__6_), .C(_2590_), .Y(_2593_) );
XOR2X1 XOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_2593_), .B(micro_ucr_hash1_b_31__7_), .Y(micro_ucr_hash1_hash_15_) );
XOR2X1 XOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(vdd), .Y(micro_ucr_hash1_a_0__0_) );
XOR2X1 XOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(micro_ucr_hash1_a_0__1_) );
XOR2X1 XOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(micro_ucr_hash1_a_0__2_) );
XOR2X1 XOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(vdd), .Y(micro_ucr_hash1_a_0__3_) );
INVX2 INVX2_68 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[88]), .Y(_2663_) );
XNOR2X1 XNOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(vdd), .Y(_2664_) );
XNOR2X1 XNOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_2664_), .B(_2663_), .Y(micro_ucr_hash1_b_1__4_) );
NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_2663_), .B(_2664_), .Y(_2665_) );
OR2X2 OR2X2_114 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2666_) );
NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2667_) );
NAND3X1 NAND3X1_355 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[89]), .B(_2667_), .C(_2666_), .Y(_2668_) );
INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[89]), .Y(_2669_) );
NOR2X1 NOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2670_) );
AND2X2 AND2X2_159 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2671_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_2671_), .B(_2670_), .C(_2669_), .Y(_2672_) );
NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_2672_), .B(_2668_), .Y(_2673_) );
XNOR2X1 XNOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_2673_), .B(_2665_), .Y(micro_ucr_hash1_b_1__5_) );
NAND3X1 NAND3X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2668_), .B(_2672_), .C(_2665_), .Y(_2674_) );
NOR3X1 NOR3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_2669_), .B(_2670_), .C(_2671_), .Y(_2675_) );
INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[90]), .Y(_2676_) );
NOR2X1 NOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2677_) );
AND2X2 AND2X2_160 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2678_) );
NOR3X1 NOR3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_2676_), .B(_2677_), .C(_2678_), .Y(_2679_) );
OR2X2 OR2X2_115 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2680_) );
NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2681_) );
AOI21X1 AOI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_2681_), .B(_2680_), .C(bloque_bytes[90]), .Y(_2682_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2679_), .B(_2682_), .C(_2675_), .Y(_2683_) );
NAND3X1 NAND3X1_357 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[90]), .B(_2681_), .C(_2680_), .Y(_2684_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_2678_), .B(_2677_), .C(_2676_), .Y(_2685_) );
NAND3X1 NAND3X1_358 ( .gnd(gnd), .vdd(vdd), .A(_2685_), .B(_2668_), .C(_2684_), .Y(_2686_) );
NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_2686_), .B(_2683_), .Y(_2687_) );
XNOR2X1 XNOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_2687_), .B(_2674_), .Y(micro_ucr_hash1_b_1__6_) );
NAND3X1 NAND3X1_359 ( .gnd(gnd), .vdd(vdd), .A(_2684_), .B(_2685_), .C(_2675_), .Y(_2688_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_2679_), .B(_2682_), .C(_2668_), .Y(_2689_) );
NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_2688_), .B(_2689_), .Y(_2690_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2690_), .B(_2674_), .C(_2688_), .Y(_2691_) );
INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[91]), .Y(_2692_) );
NOR2X1 NOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(_2693_) );
AND2X2 AND2X2_161 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(_2694_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .B(_2693_), .C(_2692_), .Y(_2695_) );
OR2X2 OR2X2_116 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(_2696_) );
NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(gnd), .Y(_2697_) );
NAND3X1 NAND3X1_360 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[91]), .B(_2697_), .C(_2696_), .Y(_2698_) );
AOI21X1 AOI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .B(_2698_), .C(_2684_), .Y(_2699_) );
NAND3X1 NAND3X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2692_), .B(_2697_), .C(_2696_), .Y(_2700_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .B(_2693_), .C(bloque_bytes[91]), .Y(_2701_) );
AOI21X1 AOI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_2701_), .B(_2700_), .C(_2679_), .Y(_2702_) );
NOR2X1 NOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_2699_), .B(_2702_), .Y(_2594_) );
XOR2X1 XOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_2691_), .B(_2594_), .Y(micro_ucr_hash1_b_1__7_) );
INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[92]), .Y(_2595_) );
OR2X2 OR2X2_117 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2596_) );
NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2597_) );
NAND3X1 NAND3X1_362 ( .gnd(gnd), .vdd(vdd), .A(_2595_), .B(_2597_), .C(_2596_), .Y(_2598_) );
NOR2X1 NOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2599_) );
AND2X2 AND2X2_162 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2600_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2600_), .B(_2599_), .C(bloque_bytes[92]), .Y(_2601_) );
NAND3X1 NAND3X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .B(_2598_), .C(_2601_), .Y(_2602_) );
AOI21X1 AOI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_2697_), .B(_2696_), .C(bloque_bytes[91]), .Y(_2603_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2600_), .B(_2599_), .C(_2595_), .Y(_2604_) );
NAND3X1 NAND3X1_364 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[92]), .B(_2597_), .C(_2596_), .Y(_2605_) );
NAND3X1 NAND3X1_365 ( .gnd(gnd), .vdd(vdd), .A(_2604_), .B(_2605_), .C(_2603_), .Y(_2606_) );
AND2X2 AND2X2_163 ( .gnd(gnd), .vdd(vdd), .A(_2606_), .B(_2602_), .Y(_2607_) );
INVX2 INVX2_69 ( .gnd(gnd), .vdd(vdd), .A(_2702_), .Y(_2608_) );
NOR2X1 NOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_2682_), .B(_2679_), .Y(_2609_) );
AOI21X1 AOI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_2675_), .B(_2609_), .C(_2699_), .Y(_2610_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_2690_), .B(_2674_), .C(_2610_), .Y(_2611_) );
NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_2608_), .B(_2611_), .Y(_2612_) );
XNOR2X1 XNOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_2612_), .B(_2607_), .Y(micro_ucr_hash1_c_0__4_) );
NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_2602_), .B(_2606_), .Y(_2613_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_2612_), .B(_2613_), .C(_2602_), .Y(_2614_) );
INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[93]), .Y(_2615_) );
OR2X2 OR2X2_118 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2616_) );
NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2617_) );
NAND3X1 NAND3X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2615_), .B(_2617_), .C(_2616_), .Y(_2618_) );
NOR2X1 NOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2619_) );
AND2X2 AND2X2_164 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2620_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .B(_2619_), .C(bloque_bytes[93]), .Y(_2621_) );
NAND3X1 NAND3X1_367 ( .gnd(gnd), .vdd(vdd), .A(_2604_), .B(_2621_), .C(_2618_), .Y(_2622_) );
AOI21X1 AOI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_2597_), .B(_2596_), .C(bloque_bytes[92]), .Y(_2623_) );
NAND3X1 NAND3X1_368 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[93]), .B(_2617_), .C(_2616_), .Y(_2624_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .B(_2619_), .C(_2615_), .Y(_2625_) );
NAND3X1 NAND3X1_369 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .B(_2624_), .C(_2623_), .Y(_2626_) );
NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_2622_), .B(_2626_), .Y(_2627_) );
INVX2 INVX2_70 ( .gnd(gnd), .vdd(vdd), .A(_2627_), .Y(_2628_) );
XNOR2X1 XNOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_2614_), .B(_2628_), .Y(micro_ucr_hash1_c_0__5_) );
AOI21X1 AOI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_2622_), .B(_2626_), .C(_2613_), .Y(_2629_) );
NAND3X1 NAND3X1_370 ( .gnd(gnd), .vdd(vdd), .A(_2608_), .B(_2629_), .C(_2611_), .Y(_2630_) );
NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_2625_), .B(_2624_), .Y(_2631_) );
OR2X2 OR2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_2631_), .B(_2623_), .Y(_2632_) );
INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(_2632_), .Y(_2633_) );
AOI21X1 AOI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2623_), .B(_2631_), .C(_2602_), .Y(_2634_) );
NOR2X1 NOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2634_), .B(_2633_), .Y(_2635_) );
INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(bloque_bytes[94]), .Y(_2636_) );
XNOR2X1 XNOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(gnd), .Y(_2637_) );
OR2X2 OR2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_2637_), .B(_2636_), .Y(_2638_) );
NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_2636_), .B(_2637_), .Y(_2639_) );
NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_2639_), .B(_2638_), .Y(_2640_) );
OR2X2 OR2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_2640_), .B(_2624_), .Y(_2641_) );
NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(_2624_), .B(_2640_), .Y(_2642_) );
NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_2642_), .B(_2641_), .Y(_2643_) );
AOI21X1 AOI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_2635_), .B(_2630_), .C(_2643_), .Y(_2644_) );
NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_2627_), .B(_2607_), .Y(_2645_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_2612_), .B(_2645_), .C(_2635_), .Y(_2646_) );
INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(_2643_), .Y(_2647_) );
NOR2X1 NOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2647_), .B(_2646_), .Y(_2648_) );
NOR2X1 NOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_2644_), .B(_2648_), .Y(micro_ucr_hash1_c_0__6_) );
INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(_2688_), .Y(_2649_) );
AOI21X1 AOI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_2608_), .B(_2649_), .C(_2699_), .Y(_2650_) );
AOI21X1 AOI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_2663_), .B(_2664_), .C(_2673_), .Y(_2651_) );
NAND3X1 NAND3X1_371 ( .gnd(gnd), .vdd(vdd), .A(_2651_), .B(_2687_), .C(_2594_), .Y(_2652_) );
AOI21X1 AOI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_2650_), .B(_2652_), .C(_2645_), .Y(_2653_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_2628_), .B(_2602_), .C(_2632_), .Y(_2654_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_2653_), .B(_2654_), .C(_2647_), .Y(_2655_) );
XOR2X1 XOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(vdd), .B(bloque_bytes[95]), .Y(_2656_) );
XNOR2X1 XNOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_2656_), .B(gnd), .Y(_2657_) );
XNOR2X1 XNOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_2657_), .B(_2638_), .Y(_2658_) );
NAND3X1 NAND3X1_372 ( .gnd(gnd), .vdd(vdd), .A(_2641_), .B(_2658_), .C(_2655_), .Y(_2659_) );
INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(_2641_), .Y(_2660_) );
INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .Y(_2661_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_2644_), .B(_2660_), .C(_2661_), .Y(_2662_) );
NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_2659_), .B(_2662_), .Y(micro_ucr_hash1_c_0__7_) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_10__0_) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_10__1_) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_10__2_) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_10__3_) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_11__0_) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_11__1_) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_11__2_) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_11__3_) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_12__0_) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_12__1_) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_12__2_) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_12__3_) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_13__0_) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_13__1_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_13__2_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_13__3_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_14__0_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_14__1_) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_14__2_) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_14__3_) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_15__0_) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_15__1_) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_15__2_) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_15__3_) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_16__0_) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_16__1_) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_16__2_) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_16__3_) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_17__0_) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_17__1_) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_17__2_) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_17__3_) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_18__0_) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_18__1_) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_18__2_) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_18__3_) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_19__0_) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_19__1_) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_19__2_) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_19__3_) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_1__0_) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_1__1_) );
BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_1__2_) );
BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_1__3_) );
BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_20__0_) );
BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_20__1_) );
BUFX2 BUFX2_72 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_20__2_) );
BUFX2 BUFX2_73 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_20__3_) );
BUFX2 BUFX2_74 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_21__0_) );
BUFX2 BUFX2_75 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_21__1_) );
BUFX2 BUFX2_76 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_21__2_) );
BUFX2 BUFX2_77 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_21__3_) );
BUFX2 BUFX2_78 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_22__0_) );
BUFX2 BUFX2_79 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_22__1_) );
BUFX2 BUFX2_80 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_22__2_) );
BUFX2 BUFX2_81 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_22__3_) );
BUFX2 BUFX2_82 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_23__0_) );
BUFX2 BUFX2_83 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_23__1_) );
BUFX2 BUFX2_84 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_23__2_) );
BUFX2 BUFX2_85 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_23__3_) );
BUFX2 BUFX2_86 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_24__0_) );
BUFX2 BUFX2_87 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_24__1_) );
BUFX2 BUFX2_88 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_24__2_) );
BUFX2 BUFX2_89 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_24__3_) );
BUFX2 BUFX2_90 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_25__0_) );
BUFX2 BUFX2_91 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_25__1_) );
BUFX2 BUFX2_92 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_25__2_) );
BUFX2 BUFX2_93 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_25__3_) );
BUFX2 BUFX2_94 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_26__0_) );
BUFX2 BUFX2_95 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_26__1_) );
BUFX2 BUFX2_96 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_26__2_) );
BUFX2 BUFX2_97 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_26__3_) );
BUFX2 BUFX2_98 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_27__0_) );
BUFX2 BUFX2_99 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_27__1_) );
BUFX2 BUFX2_100 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_27__2_) );
BUFX2 BUFX2_101 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_27__3_) );
BUFX2 BUFX2_102 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_28__0_) );
BUFX2 BUFX2_103 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_28__1_) );
BUFX2 BUFX2_104 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_28__2_) );
BUFX2 BUFX2_105 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_28__3_) );
BUFX2 BUFX2_106 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_29__0_) );
BUFX2 BUFX2_107 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_29__1_) );
BUFX2 BUFX2_108 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_29__2_) );
BUFX2 BUFX2_109 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_29__3_) );
BUFX2 BUFX2_110 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_2__0_) );
BUFX2 BUFX2_111 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_2__1_) );
BUFX2 BUFX2_112 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_2__2_) );
BUFX2 BUFX2_113 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_2__3_) );
BUFX2 BUFX2_114 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_30__0_) );
BUFX2 BUFX2_115 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_30__1_) );
BUFX2 BUFX2_116 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_30__2_) );
BUFX2 BUFX2_117 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_30__3_) );
BUFX2 BUFX2_118 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_31__0_) );
BUFX2 BUFX2_119 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_31__1_) );
BUFX2 BUFX2_120 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_31__2_) );
BUFX2 BUFX2_121 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_31__3_) );
BUFX2 BUFX2_122 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_3__0_) );
BUFX2 BUFX2_123 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_3__1_) );
BUFX2 BUFX2_124 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_3__2_) );
BUFX2 BUFX2_125 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_3__3_) );
BUFX2 BUFX2_126 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_4__0_) );
BUFX2 BUFX2_127 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_4__1_) );
BUFX2 BUFX2_128 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_4__2_) );
BUFX2 BUFX2_129 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_4__3_) );
BUFX2 BUFX2_130 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_5__0_) );
BUFX2 BUFX2_131 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_5__1_) );
BUFX2 BUFX2_132 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_5__2_) );
BUFX2 BUFX2_133 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_5__3_) );
BUFX2 BUFX2_134 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_6__0_) );
BUFX2 BUFX2_135 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_6__1_) );
BUFX2 BUFX2_136 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_6__2_) );
BUFX2 BUFX2_137 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_6__3_) );
BUFX2 BUFX2_138 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_7__0_) );
BUFX2 BUFX2_139 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_7__1_) );
BUFX2 BUFX2_140 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_7__2_) );
BUFX2 BUFX2_141 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_7__3_) );
BUFX2 BUFX2_142 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_8__0_) );
BUFX2 BUFX2_143 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_8__1_) );
BUFX2 BUFX2_144 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_8__2_) );
BUFX2 BUFX2_145 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_8__3_) );
BUFX2 BUFX2_146 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_9__0_) );
BUFX2 BUFX2_147 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_9__1_) );
BUFX2 BUFX2_148 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_9__2_) );
BUFX2 BUFX2_149 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(micro_ucr_hash1_b_9__3_) );
BUFX2 BUFX2_150 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__4_), .Y(micro_ucr_hash1_c_0__0_) );
BUFX2 BUFX2_151 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__5_), .Y(micro_ucr_hash1_c_0__1_) );
BUFX2 BUFX2_152 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__6_), .Y(micro_ucr_hash1_c_0__2_) );
BUFX2 BUFX2_153 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_1__7_), .Y(micro_ucr_hash1_c_0__3_) );
BUFX2 BUFX2_154 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__4_), .Y(micro_ucr_hash1_c_10__0_) );
BUFX2 BUFX2_155 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__5_), .Y(micro_ucr_hash1_c_10__1_) );
BUFX2 BUFX2_156 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__6_), .Y(micro_ucr_hash1_c_10__2_) );
BUFX2 BUFX2_157 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_11__7_), .Y(micro_ucr_hash1_c_10__3_) );
BUFX2 BUFX2_158 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__4_), .Y(micro_ucr_hash1_c_12__0_) );
BUFX2 BUFX2_159 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__5_), .Y(micro_ucr_hash1_c_12__1_) );
BUFX2 BUFX2_160 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__6_), .Y(micro_ucr_hash1_c_12__2_) );
BUFX2 BUFX2_161 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_13__7_), .Y(micro_ucr_hash1_c_12__3_) );
BUFX2 BUFX2_162 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__4_), .Y(micro_ucr_hash1_c_14__0_) );
BUFX2 BUFX2_163 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__5_), .Y(micro_ucr_hash1_c_14__1_) );
BUFX2 BUFX2_164 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__6_), .Y(micro_ucr_hash1_c_14__2_) );
BUFX2 BUFX2_165 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_15__7_), .Y(micro_ucr_hash1_c_14__3_) );
BUFX2 BUFX2_166 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__4_), .Y(micro_ucr_hash1_c_16__0_) );
BUFX2 BUFX2_167 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__5_), .Y(micro_ucr_hash1_c_16__1_) );
BUFX2 BUFX2_168 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__6_), .Y(micro_ucr_hash1_c_16__2_) );
BUFX2 BUFX2_169 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_17__7_), .Y(micro_ucr_hash1_c_16__3_) );
BUFX2 BUFX2_170 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__4_), .Y(micro_ucr_hash1_c_18__0_) );
BUFX2 BUFX2_171 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__5_), .Y(micro_ucr_hash1_c_18__1_) );
BUFX2 BUFX2_172 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__6_), .Y(micro_ucr_hash1_c_18__2_) );
BUFX2 BUFX2_173 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_19__7_), .Y(micro_ucr_hash1_c_18__3_) );
BUFX2 BUFX2_174 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__4_), .Y(micro_ucr_hash1_c_20__0_) );
BUFX2 BUFX2_175 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__5_), .Y(micro_ucr_hash1_c_20__1_) );
BUFX2 BUFX2_176 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__6_), .Y(micro_ucr_hash1_c_20__2_) );
BUFX2 BUFX2_177 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_21__7_), .Y(micro_ucr_hash1_c_20__3_) );
BUFX2 BUFX2_178 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__4_), .Y(micro_ucr_hash1_c_22__0_) );
BUFX2 BUFX2_179 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__5_), .Y(micro_ucr_hash1_c_22__1_) );
BUFX2 BUFX2_180 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__6_), .Y(micro_ucr_hash1_c_22__2_) );
BUFX2 BUFX2_181 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_23__7_), .Y(micro_ucr_hash1_c_22__3_) );
BUFX2 BUFX2_182 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__4_), .Y(micro_ucr_hash1_c_24__0_) );
BUFX2 BUFX2_183 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__5_), .Y(micro_ucr_hash1_c_24__1_) );
BUFX2 BUFX2_184 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__6_), .Y(micro_ucr_hash1_c_24__2_) );
BUFX2 BUFX2_185 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_25__7_), .Y(micro_ucr_hash1_c_24__3_) );
BUFX2 BUFX2_186 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__4_), .Y(micro_ucr_hash1_c_26__0_) );
BUFX2 BUFX2_187 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__5_), .Y(micro_ucr_hash1_c_26__1_) );
BUFX2 BUFX2_188 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__6_), .Y(micro_ucr_hash1_c_26__2_) );
BUFX2 BUFX2_189 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_27__7_), .Y(micro_ucr_hash1_c_26__3_) );
BUFX2 BUFX2_190 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__4_), .Y(micro_ucr_hash1_c_28__0_) );
BUFX2 BUFX2_191 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__5_), .Y(micro_ucr_hash1_c_28__1_) );
BUFX2 BUFX2_192 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__6_), .Y(micro_ucr_hash1_c_28__2_) );
BUFX2 BUFX2_193 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_29__7_), .Y(micro_ucr_hash1_c_28__3_) );
BUFX2 BUFX2_194 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__4_), .Y(micro_ucr_hash1_c_2__0_) );
BUFX2 BUFX2_195 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__5_), .Y(micro_ucr_hash1_c_2__1_) );
BUFX2 BUFX2_196 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__6_), .Y(micro_ucr_hash1_c_2__2_) );
BUFX2 BUFX2_197 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_3__7_), .Y(micro_ucr_hash1_c_2__3_) );
BUFX2 BUFX2_198 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__4_), .Y(micro_ucr_hash1_c_30__0_) );
BUFX2 BUFX2_199 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__5_), .Y(micro_ucr_hash1_c_30__1_) );
BUFX2 BUFX2_200 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__6_), .Y(micro_ucr_hash1_c_30__2_) );
BUFX2 BUFX2_201 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_31__7_), .Y(micro_ucr_hash1_c_30__3_) );
BUFX2 BUFX2_202 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__4_), .Y(micro_ucr_hash1_c_4__0_) );
BUFX2 BUFX2_203 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__5_), .Y(micro_ucr_hash1_c_4__1_) );
BUFX2 BUFX2_204 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__6_), .Y(micro_ucr_hash1_c_4__2_) );
BUFX2 BUFX2_205 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_5__7_), .Y(micro_ucr_hash1_c_4__3_) );
BUFX2 BUFX2_206 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__4_), .Y(micro_ucr_hash1_c_6__0_) );
BUFX2 BUFX2_207 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__5_), .Y(micro_ucr_hash1_c_6__1_) );
BUFX2 BUFX2_208 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__6_), .Y(micro_ucr_hash1_c_6__2_) );
BUFX2 BUFX2_209 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_7__7_), .Y(micro_ucr_hash1_c_6__3_) );
BUFX2 BUFX2_210 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__4_), .Y(micro_ucr_hash1_c_8__0_) );
BUFX2 BUFX2_211 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__5_), .Y(micro_ucr_hash1_c_8__1_) );
BUFX2 BUFX2_212 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__6_), .Y(micro_ucr_hash1_c_8__2_) );
BUFX2 BUFX2_213 ( .gnd(gnd), .vdd(vdd), .A(micro_ucr_hash1_b_9__7_), .Y(micro_ucr_hash1_c_8__3_) );
endmodule
